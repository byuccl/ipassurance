module grethm
   (rst,
    clk,
    .\ahbmi[hgrant] ({ahbmi[0],ahbmi[1],ahbmi[2],ahbmi[3],ahbmi[4],ahbmi[5],ahbmi[6],ahbmi[7],ahbmi[8],ahbmi[9],ahbmi[10],ahbmi[11],ahbmi[12],ahbmi[13],ahbmi[14],ahbmi[15]}),
    \ahbmi[hready] ,
    \ahbmi[hresp] ,
    \ahbmi[hrdata] ,
    \ahbmi[hirq] ,
    \ahbmi[testen] ,
    \ahbmi[testrst] ,
    \ahbmi[scanen] ,
    \ahbmi[testoen] ,
    \ahbmi[testin] ,
    .\ahbmo[hbusreq] (ahbmo),
    \ahbmo[hlock] ,
    \ahbmo[htrans] ,
    \ahbmo[haddr] ,
    \ahbmo[hwrite] ,
    \ahbmo[hsize] ,
    \ahbmo[hburst] ,
    \ahbmo[hprot] ,
    \ahbmo[hwdata] ,
    \ahbmo[hirq] ,
    \ahbmo[hconfig][0] ,
    \ahbmo[hconfig][1] ,
    \ahbmo[hconfig][2] ,
    \ahbmo[hconfig][3] ,
    \ahbmo[hconfig][4] ,
    \ahbmo[hconfig][5] ,
    \ahbmo[hconfig][6] ,
    \ahbmo[hconfig][7] ,
    \ahbmo[hindex] ,
    .\apbi[psel] ({apbi[0],apbi[1],apbi[2],apbi[3],apbi[4],apbi[5],apbi[6],apbi[7],apbi[8],apbi[9],apbi[10],apbi[11],apbi[12],apbi[13],apbi[14],apbi[15]}),
    \apbi[penable] ,
    \apbi[paddr] ,
    \apbi[pwrite] ,
    \apbi[pwdata] ,
    \apbi[pirq] ,
    \apbi[testen] ,
    \apbi[testrst] ,
    \apbi[scanen] ,
    \apbi[testoen] ,
    \apbi[testin] ,
    \apbo[prdata] ,
    \apbo[pirq] ,
    \apbo[pconfig][0] ,
    \apbo[pconfig][1] ,
    \apbo[pindex] ,
    \ethi[gtx_clk] ,
    .\ethi[rmii_clk] (ethi),
    \ethi[tx_clk] ,
    \ethi[tx_clk_90] ,
    \ethi[tx_dv] ,
    \ethi[rx_clk] ,
    \ethi[rxd] ,
    \ethi[rx_dv] ,
    \ethi[rx_er] ,
    \ethi[rx_col] ,
    \ethi[rx_crs] ,
    \ethi[rx_en] ,
    \ethi[mdio_i] ,
    \ethi[mdint] ,
    \ethi[phyrstaddr] ,
    \ethi[edcladdr] ,
    \ethi[edclsepahb] ,
    \ethi[edcldisable] ,
    \etho[reset] ,
    \etho[txd] ,
    \etho[tx_en] ,
    \etho[tx_er] ,
    \etho[tx_clk] ,
    \etho[mdc] ,
    \etho[mdio_o] ,
    \etho[mdio_oe] ,
    \etho[gbit] ,
    \etho[speed] );
  (* sync_set_reset = "true" *) input rst;
  input clk;
  input \ahbmi[hready] ;
  input [1:0]\ahbmi[hresp] ;
  input [31:0]\ahbmi[hrdata] ;
  input [31:0]\ahbmi[hirq] ;
  input \ahbmi[testen] ;
  input \ahbmi[testrst] ;
  input \ahbmi[scanen] ;
  input \ahbmi[testoen] ;
  input [3:0]\ahbmi[testin] ;
  output \ahbmo[hlock] ;
  output [1:0]\ahbmo[htrans] ;
  output [31:0]\ahbmo[haddr] ;
  output \ahbmo[hwrite] ;
  output [2:0]\ahbmo[hsize] ;
  output [2:0]\ahbmo[hburst] ;
  output [3:0]\ahbmo[hprot] ;
  output [31:0]\ahbmo[hwdata] ;
  output [31:0]\ahbmo[hirq] ;
  output [31:0]\ahbmo[hconfig][0] ;
  output [31:0]\ahbmo[hconfig][1] ;
  output [31:0]\ahbmo[hconfig][2] ;
  output [31:0]\ahbmo[hconfig][3] ;
  output [31:0]\ahbmo[hconfig][4] ;
  output [31:0]\ahbmo[hconfig][5] ;
  output [31:0]\ahbmo[hconfig][6] ;
  output [31:0]\ahbmo[hconfig][7] ;
  output [3:0]\ahbmo[hindex] ;
  input \apbi[penable] ;
  input [31:0]\apbi[paddr] ;
  input \apbi[pwrite] ;
  input [31:0]\apbi[pwdata] ;
  input [31:0]\apbi[pirq] ;
  input \apbi[testen] ;
  input \apbi[testrst] ;
  input \apbi[scanen] ;
  input \apbi[testoen] ;
  input [3:0]\apbi[testin] ;
  output [31:0]\apbo[prdata] ;
  output [31:0]\apbo[pirq] ;
  output [31:0]\apbo[pconfig][0] ;
  output [31:0]\apbo[pconfig][1] ;
  output [3:0]\apbo[pindex] ;
  input \ethi[gtx_clk] ;
  input \ethi[tx_clk] ;
  input \ethi[tx_clk_90] ;
  input \ethi[tx_dv] ;
  input \ethi[rx_clk] ;
  input [7:0]\ethi[rxd] ;
  input \ethi[rx_dv] ;
  input \ethi[rx_er] ;
  input \ethi[rx_col] ;
  input \ethi[rx_crs] ;
  input \ethi[rx_en] ;
  input \ethi[mdio_i] ;
  input \ethi[mdint] ;
  input [4:0]\ethi[phyrstaddr] ;
  input [3:0]\ethi[edcladdr] ;
  input \ethi[edclsepahb] ;
  input \ethi[edcldisable] ;
  output \etho[reset] ;
  output [7:0]\etho[txd] ;
  output \etho[tx_en] ;
  output \etho[tx_er] ;
  output \etho[tx_clk] ;
  output \etho[mdc] ;
  output \etho[mdio_o] ;
  output \etho[mdio_oe] ;
  output \etho[gbit] ;
  output \etho[speed] ;
  input [0:15]ahbmi;
  output ahbmo;
  input [0:15]apbi;
  input ethi;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[def_state][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[def_state][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[def_state][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[def_state][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[def_state][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[main_state][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r[rx_state][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_gmiimode0.r_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire FSM_sequential_r;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[edclrstate][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[mdio_state][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[mdio_state][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[mdio_state][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[mdio_state][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[mdio_state][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[mdio_state][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[mdio_state][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[mdio_state][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[regaddr][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[regaddr][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[regaddr][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[regaddr][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[regaddr][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[regaddr][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r[rxdstate][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]FSM_sequential_r_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_16_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_16_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_22_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_22_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_30_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_30_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_31_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_31_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_31_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_38_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_38_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_38_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_43_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_43_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[edclrstate][3]_i_43_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[mdio_state][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_reg[regaddr][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire GND_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire VCC_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_101__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_101_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_103_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_104_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_105_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_107__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_107_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_108_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_110_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_111_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_111_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_111_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_111_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_111_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_111_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_111_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_111_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_114_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_19__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_20__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_21__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_23__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_24__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_25__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_26__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_27__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_28__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_29__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_30__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_31__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_32__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_33__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_34__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_34__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_35__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_36__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_37__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_38__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_39__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_40__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_41__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_42__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_43__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_44__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_45__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_46__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_47__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_48__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_49__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_50__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_51__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_52__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_53__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_54__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_55__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_56__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_57__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_58__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_60__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_61__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_62__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_63__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_64__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_65__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_66__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_67__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_68__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_69__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_70__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_71__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_72__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_73__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_73__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_73__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_73__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_73__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_73__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_73__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_73__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_74__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_75__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_76__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_77__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_78__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_79__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_80_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_81__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_82__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_83__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_84__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_85__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_86__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_86__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_86__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_86__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_86__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_86__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_86__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_86__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_87__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_87__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_87__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_87__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_87__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_87__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_87__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_87__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_88__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_89__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_90__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_91__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_92__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_93__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_93_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_94__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_94_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_95_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_96_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_97__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_97_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_98__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \a9.x[0].r0_i_99_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [0:15]ahbmi;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\ahbmi[hrdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ahbmi[hready] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\ahbmi[hresp] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ahbmo;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:1]\^ahbmo[haddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\ahbmo[htrans] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ahbmo[htrans][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\ahbmo[hwdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ahbmo[hwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [0:15]apbi;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\apbi[paddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbi[penable] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\apbi[pwdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbi[pwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire apbo;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [12:12]\^apbo[pirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[pirq][12]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[pirq][12]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\apbo[prdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][0]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][10]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][10]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][10]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][10]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][10]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][11]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][11]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][11]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][12]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][12]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][12]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][13]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][13]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][13]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][14]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][14]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][14]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][14]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][14]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][15]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][15]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][15]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][16]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][17]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][18]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][19]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][1]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][20]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][21]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][22]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][23]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][24]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][25]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][26]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][27]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][28]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][28]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][29]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][2]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][2]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][30]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][30]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][31]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][31]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][3]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][3]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][3]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][4]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][4]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][4]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][5]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][5]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][5]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][6]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][6]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][6]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][7]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][7]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][7]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][8]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][8]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][8]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][9]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][9]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][9]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][9]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ethi;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ethi[mdio_i] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ethi[rx_crs] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]\ethi[rxd] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire etho;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \etho[mdc] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \etho[mdio_o] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \etho[mdio_oe] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \etho[reset] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \etho[speed] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \etho[tx_en] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\^etho[txd] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][0]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][10]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][10]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][10]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][3]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][5]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][6]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][6]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][8]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][9]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[byte_count][9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[cnt][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[cnt][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[cnt][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[cnt][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[cnt][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[cnt][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[cnt][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[cnt][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[cnt][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[cnt][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[cnt][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][11]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][13]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][24]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][25]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][26]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][31]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crc_en]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[crs_act]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[data][27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[data][31]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[data][31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[deferring]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[delay_val][9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[done]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[done]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[done]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[dv]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[enold]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[got4b]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[gotframe]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[icnt][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[icnt][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ifg_cycls][8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[ltfound]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[odd_nibble]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[odd_nibble]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[random][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[rcnt][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[rcnt][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[rcnt][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[rcnt][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[read]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[read]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[read]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[restart]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[restart]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[retry_cnt][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[retry_cnt][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[rmii_crc_en]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[rxd2][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[rxd2][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[rxdp][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[rxdp][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[slot_count][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[slot_count][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[slot_count][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[start][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[start][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[start]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[start]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][0]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][1]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[status][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[switch]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[sync_start]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[sync_start]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[sync_start]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[transmitting]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[tx_en]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[tx_en]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[tx_en]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[tx_en]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[tx_en]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[tx_en]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[tx_en]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[tx_en]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[tx_en]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[tx_en]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[tx_en]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[tx_en]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][0]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][1]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][1]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][1]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[txd][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[write]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[zero]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r[zero]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\gmiimode0.r_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][3]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][3]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][3]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][3]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][3]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][3]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][7]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][7]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][7]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][7]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][7]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][7]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[byte_count][7]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[tx_en]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[tx_en]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[tx_en]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[tx_en]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[txd][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[txd][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \gmiimode0.r_reg[txd][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\m100.u0/datain ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_53 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_54 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_55 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_56 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_57 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_53 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_54 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_55 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_56 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_57 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [8:0]\m100.u0/eraddress ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\m100.u0/erdata ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/erenable ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\m100.u0/ethc0/a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/ahb0/nbo ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/ahb0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/ahb0/r_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/ahb0/r_reg[bb]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/ahb0/r_reg[bg]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/ahb0/r_reg[bo]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/ahb0/r_reg[error]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/ahb0/r_reg[retry]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/ahb0/v ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\m100.u0/ethc0/crcadder ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\m100.u0/ethc0/d ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/data1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/data2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\m100.u0/ethc0/p_0_in0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/p_0_in153_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/p_0_in1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/p_116_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [17:0]\m100.u0/ethc0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/p_1_in128_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/p_1_in143_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/p_1_in4_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]\m100.u0/ethc0/p_6_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[abufs_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[abufs_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[addrdone]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[addrok_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [9:0]\m100.u0/ethc0/r_reg[applength]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[bcast_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[capbil_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[capbil_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[check]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\m100.u0/ethc0/r_reg[checkdata]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[cnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[cnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[cnt_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[cnt_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[cnt_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ctrlpkt]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ecnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ecnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ecnt_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ecnt_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclactive_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclbcast]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[edclip_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/r_reg[edclrstate] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[emacaddr_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[erxidle]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[etxidle]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ewr]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[gotframe_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[init_busy_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[ipcrc_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mac_addr_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][busy]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][linkfail_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][phyadr_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][phyadr_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][phyadr_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[mdio_ctrl][write]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/r_reg[mdio_state] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[msbgood_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[nak_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[oplen_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[oplen_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[oplen_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[oplen_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[oplen_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[oplen_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[oplen_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[oplen_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[oplen_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[oplen_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[phywr]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\m100.u0/ethc0/r_reg[regaddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rfcnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rfcnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rfrpnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rfrpnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:1]\m100.u0/ethc0/r_reg[rmsto][addr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][data_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][req_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rmsto][write_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rstaneg_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rstphy]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxaddr_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxburstav]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxburstcnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxburstcnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:0]\m100.u0/ethc0/r_reg[rxbytecount]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxden]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdesc_n_0_][31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdone] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdoneack]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdoneold]__1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdsel_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdsel_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdsel_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdsel_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdsel_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdsel_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxdsel_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\m100.u0/ethc0/r_reg[rxdstate] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxirq]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxlength_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxlength_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxlength_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxlength_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxlength_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxlength_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxlength_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxlength_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxlength_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxlength_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxlength_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\m100.u0/ethc0/r_reg[rxstart]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxstatus_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxstatus_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxstatus_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxwrap_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[rxwriteack]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [13:0]\m100.u0/ethc0/r_reg[seq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[status][invaddr_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[status][rx_err_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[status][rx_int_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[status][rxahberr_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[status][toosmall_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[status][tx_err_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[status][tx_int_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[status][txahberr_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tarp]0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tarp]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tcnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tcnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tcnt_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tcnt_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tcnt_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tcnt_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tcnt_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tedcl]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tfcnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tfcnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tfcnt_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tfcnt_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tfcnt_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tfcnt_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tfcnt_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tfcnt_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:1]\m100.u0/ethc0/r_reg[tmsto][addr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][data_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][req_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tmsto][write_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[tnak]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [29:0]\m100.u0/ethc0/r_reg[txaddr]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txburstav]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txburstcnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txburstcnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txcnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txcnt_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txcnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txcnt_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txcnt_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txcnt_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txcnt_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txcnt_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txcnt_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txcnt_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txcnt_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdata_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdataav_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txden]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\m100.u0/ethc0/r_reg[txdesc]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\m100.u0/ethc0/r_reg[txdone]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdsel_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdsel_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdsel_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdsel_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdsel_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdsel_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdsel_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdstate_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdstate_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdstate_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txdstate_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txirq]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txirqgen_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txlength_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txlength_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txlength_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txlength_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txlength_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txlength_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txlength_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txlength_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txlength_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txlength_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txlength_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txread] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txreadack]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\m100.u0/ethc0/r_reg[txrestart]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txstart]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txstart_sync_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txstatus_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txstatus_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txvalid_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[txwrap_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[udpsrc_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[write_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[write_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[write_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[write_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/r_reg[writeok_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rin ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rin[status][txahberr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rin[tmsto][req] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rmsti ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rmsti[grant] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rmsti[ready] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rmsti[retry] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/crc_en ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:16]\m100.u0/ethc0/rx_rmii1.rx0/d ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/dv17_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r[lentype][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r[lentype][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[done_ack_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dv]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[en]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[enold]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][11]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][11]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][11]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[ltfound_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[odd_nibble_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[start]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[write_ack] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_0_in10_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_0_in12_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_0_in15_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_10_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_11_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_13_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_14_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_15_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_16_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_17_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_18_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_19_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_1_in6_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_20_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_22_in55_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_23_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_24_in59_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_25_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_26_in64_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_27_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_28_in69_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_29_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_30_in72_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_31_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_32_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_33_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [27:24]\m100.u0/ethc0/rx_rmii1.rx0/p_4_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/p_9_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\m100.u0/ethc0/rx_rmii1.rx0/plusOp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/rstout0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/rxrst ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/v ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:0]\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/rx_rmii1.rx0/v[cnt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:3]\m100.u0/ethc0/rx_rmii1.rx0/v[data] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/v[got4b] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/v[status] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rx_rmii1.rx0/write_req ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rxo ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:0]\m100.u0/ethc0/rxo[byte_count] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rxo[gotframe] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\m100.u0/ethc0/rxo[lentype] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rxo[start] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/rxo[status] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/rxo[write] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/setmz ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/setmz11_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/swap ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/swap12_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tmsti ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tmsti[ready] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tmsti[retry] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [9:4]\m100.u0/ethc0/tx_rmii1.tx0/conv_integer ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [8:0]\m100.u0/ethc0/tx_rmii1.tx0/d ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/frame_waiting ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_act]__1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_prev_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[deferring_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[read_ack] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[transmitting]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_0_in10_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_0_in38_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_0_in74_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_10_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_11_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_12_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_13_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_14_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/tx_rmii1.tx0/p_15_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/tx_rmii1.tx0/p_16_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_17_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/tx_rmii1.tx0/p_18_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/tx_rmii1.tx0/p_19_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_1_in75_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/tx_rmii1.tx0/p_20_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_22_in55_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_23_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_24_in59_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_25_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_26_in64_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_27_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_28_in69_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_28_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_30_in72_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_31_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_31_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_32_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_33_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_5_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_5_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_7_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_8_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/p_9_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/rin ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/rin[fullduplex] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/rin[speed] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\m100.u0/ethc0/tx_rmii1.tx0/rin[txd_msb] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/speed ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/rstout0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/txrst ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [9:0]\m100.u0/ethc0/tx_rmii1.tx0/v ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/tx_rmii1.tx0/v[cnt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\m100.u0/ethc0/tx_rmii1.tx0/v[crc] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/v[data] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [9:1]\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/v[ifg_cycls] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\m100.u0/ethc0/tx_rmii1.tx0/v[rcnt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:1]\m100.u0/ethc0/tx_rmii1.tx0/v[retry_cnt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [6:0]\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/v[switch]3_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/v[tx_en] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]14_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]9_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/tx_rmii1.tx0/v[zero]7_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/txo ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/txo[read] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/txo[restart] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\m100.u0/ethc0/txo[status] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\m100.u0/ethc0/v[abufs] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[addrok] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[addrok]62_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[check] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[cnt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[ctrl][rxen] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[ctrl][txen] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[ctrlpkt]68_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[ctrlpkt]69_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:1]\m100.u0/ethc0/v[ecnt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[edclactive]58_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[edclip] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[edclrstate] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[edclrstate]0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[edclrstate]01_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[edclrstate]1121_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[edclrstate]1124_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[edclrstate]2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[edclrstate]2126_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [47:31]\m100.u0/ethc0/v[emacaddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [17:0]\m100.u0/ethc0/v[ipcrc] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [47:31]\m100.u0/ethc0/v[mac_addr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\m100.u0/ethc0/v[mdccnt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[mdio_ctrl][busy] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[mdio_ctrl][busy]0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[mdio_ctrl][write]1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[mdio_ctrl][write]113_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[mdioen] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[mdioo] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[mdioo]5_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[nak] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[nak]1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[phywr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [6:0]\m100.u0/ethc0/v[rcntl] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [6:0]\m100.u0/ethc0/v[rcntm] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rcntm]0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[regaddr]1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\m100.u0/ethc0/v[rfcnt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\m100.u0/ethc0/v[rfcnt]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:2]\m100.u0/ethc0/v[rmsto][addr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [18:0]\m100.u0/ethc0/v[rmsto][data] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rmsto][req] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rmsto][req]2136_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rmsto][req]2137_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rmsto][req]57_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rmsto][write] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rpnt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rxaddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rxburstav] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rxbytecount] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:0]\m100.u0/ethc0/v[rxcnt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [9:3]\m100.u0/ethc0/v[rxdsel] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rxlength] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rxstatus] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rxstatus]1135_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rxstatus]2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rxstatus]2130_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[rxwrap] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[seq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[status][invaddr]45_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[status][rx_err]15_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[status][rx_err]18_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[status][rx_int]26_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[status][rxahberr]32_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[status][toosmall]2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[status][toosmall]39_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[status][toosmall]42_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[tfrpnt]1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\m100.u0/ethc0/v[tfwpnt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[tmsto][data] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[tmsto][req]0139_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[tmsto][req]1149_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[txdsel] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[txirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[udpsrc] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[writeok]1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/v[writeok]154_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ethc0/veri ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [6:0]\m100.u0/ewaddressl ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [8:0]\m100.u0/ewaddressm ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ewritel ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/ewritem ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[addrok]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[bcast]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[ctrl][edcldis]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[ctrl][full_duplex]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[ctrl][rxen]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[ctrl][speed]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[ctrl][txen]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[ctrlpkt]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[disableduplex]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[edclactive]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[edclbcast]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[erenable]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[erxidle]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[gotframe]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[init_busy]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[mdio_ctrl][busy]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[mdio_ctrl][linkfail]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[mdio_ctrl][read]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[mdio_ctrl][write]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[mdioclk]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[mdioen]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[mdioo]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[msbgood]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[phywr]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[rmsto][write]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[rstaneg]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[rstphy]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[rxden]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[rxdoneack]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[rxirq]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[rxwrap]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[status][invaddr]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[status][rx_err]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[status][rx_int]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[status][rxahberr]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[status][toosmall]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[status][tx_err]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[status][tx_int]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[status][txahberr]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[tarp]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[tedcl]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[tmsto][write]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[tnak]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[txden]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[txirq]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[txirqgen]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[txstart]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[txstart_sync]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[txwrap]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/r[writeok]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\m100.u0/rxraddress ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\m100.u0/rxrdata ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\m100.u0/rxwaddress ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\m100.u0/rxwdata ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/rxwrite ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [6:0]\m100.u0/txraddress ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\m100.u0/txrdata ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/txrenable ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [6:0]\m100.u0/txwaddress ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\m100.u0/txwdata ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m100.u0/txwrite ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]p_0_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[abufs][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[addrdone]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[addrok]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[addrok]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[addrok]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[addrok]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[addrok]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[addrok]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[addrok]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[applength][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[applength][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[applength][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[applength][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[applength][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[applength][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[applength][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[applength][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[applength][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[applength][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ba]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ba]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bb]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bb]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bb]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bb]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bcast]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bcast]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bcast]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bcast]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bcast]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bcast]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bcast]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bcast]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bcast]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bcast]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bg]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[bo]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[capbil][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[capbil][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[capbil][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[capbil][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[capbil][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cnt][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrl][full_duplex]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrl][full_duplex]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrl][rxen]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrl][rxen]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrl][rxen]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrl][speed]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrl][speed]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrl][txen]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrl][txen]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrlpkt]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrlpkt]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrlpkt]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ctrlpkt]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[duplexstate][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[duplexstate][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[duplexstate][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[duplexstate][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[duplexstate][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[duplexstate][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[duplexstate][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[duplexstate][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ecnt][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ecnt][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ecnt][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[edclactive]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[edclactive]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[edclactive]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[edclactive]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[edclactive]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[edclactive]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[edclactive]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[edclactive]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[edclactive]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[edclbcast]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[emacaddr][31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[error]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[erxidle]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[erxidle]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ewr]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[init_busy]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][11]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][11]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][11]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][11]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][11]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][11]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][11]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][15]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][15]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][15]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][7]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][7]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][7]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][7]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][7]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][7]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipcrc][7]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdccnt][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][busy]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][busy]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][busy]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][busy]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][busy]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][10]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][10]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][10]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][11]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][11]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][11]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][11]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][12]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][12]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][12]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][12]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][12]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][13]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][13]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][13]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][13]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][13]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][13]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][14]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][14]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][14]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][14]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][14]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][14]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][4]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][4]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][5]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][5]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][5]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][6]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][6]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][6]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][7]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][8]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][8]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][8]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][9]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][9]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][9]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][data][9]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][linkfail]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][linkfail]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][phyadr][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][phyadr][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][read]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][read]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][regadr][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][regadr][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][regadr][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][regadr][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][regadr][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][regadr][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][write]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][write]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][write]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][write]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][write]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdio_ctrl][write]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioclk]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioen]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[mdioo]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[msbgood]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[nak]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[nak]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[nak]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[nak]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[nak]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[nak]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[phywr]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[phywr]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][4]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][4]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][5]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntl][6]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][4]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][4]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][4]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][4]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][4]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][5]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][5]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][5]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][5]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][5]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][5]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][5]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rcntm][6]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[retry]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfcnt][2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfcnt][2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfcnt][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfcnt][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfcnt][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfcnt][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfcnt][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfrpnt][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfrpnt][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfrpnt][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfrpnt][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfrpnt][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfrpnt][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfrpnt][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfrpnt][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfwpnt][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rfwpnt][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][13]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][17]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][1]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][21]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][21]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][25]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][25]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][addr][9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][data][18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][data][31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rmsto][req]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rpnt][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rpnt][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rpnt][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rstaneg]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxburstcnt][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxburstcnt][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxburstcnt][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxbytecount][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxbytecount][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxbytecount][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxbytecount][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxbytecount][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxbytecount][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxbytecount][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxbytecount][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxbytecount][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxbytecount][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxbytecount][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][10]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxcnt][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxdesc][31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxdoneold]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxdsel][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxdsel][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxdsel][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxdsel][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxdsel][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxdsel][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxdsel][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxdsel][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxdsel][9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][10]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][10]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][10]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][10]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxlength][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstart][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstart][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[rxstatus][4]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[seq][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][invaddr]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][rx_int]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][toosmall]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][tx_int]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[status][txahberr]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tarp]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tarp]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tarp]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tarp]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][4]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][4]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tcnt][6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tedcl]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfcnt][7]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfrpnt][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfrpnt][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfrpnt][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfrpnt][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfrpnt][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfrpnt][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfrpnt][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfrpnt][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfrpnt][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfrpnt][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfrpnt][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfrpnt][6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfwpnt][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfwpnt][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfwpnt][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfwpnt][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfwpnt][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfwpnt][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfwpnt][6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfwpnt][6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfwpnt][6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tfwpnt][6]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][13]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][17]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][21]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][25]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][29]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][29]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][29]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][29]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][29]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][29]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][29]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][29]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][29]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][5]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][addr][9]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][data][14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][data][14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][data][15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][data][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][data][31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][data][31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][data][31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][data][31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][data][31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][req]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][write]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][write]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][write]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][write]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][write]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][write]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][write]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tmsto][write]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tpnt][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[tpnt][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txaddr][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txburstav]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txburstav]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txburstav]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txburstav]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txburstcnt][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txburstcnt][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txburstcnt][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txburstcnt][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txburstcnt][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][10]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][10]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][10]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][6]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][6]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][6]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][9]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txcnt][9]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdataav]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdone][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdone][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdsel][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdsel][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdsel][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdsel][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdsel][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdsel][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdsel][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdsel][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdsel][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdsel][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdsel][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdsel][9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txdstate][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][10]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txlength][9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txrestart][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txstart]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txstart]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txstart_sync]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txstart_sync]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txstart_sync]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txstart_sync]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txstatus][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txstatus][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[txstatus][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[udpsrc][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[write][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[write][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[write][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[write][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[write][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[writeok]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]r_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[addrok]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[addrok]_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[addrok]_i_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[addrok]_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[edclactive]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[edclactive]_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[edclactive]_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[edclactive]_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[edclactive]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[edclactive]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[edclactive]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[edclactive]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][11]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][11]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][11]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][11]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][11]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][11]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][15]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][15]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][15]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][15]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][15]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][15]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][16]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][16]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][17]_i_4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][17]_i_4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][3]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][3]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][3]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][3]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][3]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][3]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][7]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][7]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][7]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][7]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][7]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ipcrc][7]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[mdio_ctrl][write]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[mdioo]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[msbgood]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[msbgood]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[msbgood]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[msbgood]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[msbgood]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[msbgood]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[msbgood]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[msbgood]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[msbgood]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[msbgood]_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[msbgood]_i_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[msbgood]_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[nak]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[nak]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[nak]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[nak]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[nak]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[nak]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[nak]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_10_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_10_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_10_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_10_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][13]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_10_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_10_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_10_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_10_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][17]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_10_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_10_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_10_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_10_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][1]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_10_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_10_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_10_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_10_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][21]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_10_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_10_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_10_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_10_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][25]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][29]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][29]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][29]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][29]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][29]_i_8_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][29]_i_8_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][29]_i_8_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][29]_i_8_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_10_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_10_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_10_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_10_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][5]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_10_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_10_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_10_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_10_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][addr][9]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_15_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_15_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_15_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rmsto][req]_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rxcnt][10]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rxcnt][10]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rxcnt][10]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rxcnt][10]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rxcnt][10]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rxcnt][10]_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rxcnt][10]_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rxcnt][10]_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rxstatus][4]_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rxstatus][4]_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[rxstatus][4]_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[seq][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[status][toosmall]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[status][toosmall]_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[status][toosmall]_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[status][toosmall]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[status][toosmall]_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[status][toosmall]_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[status][toosmall]_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][3]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][7]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][7]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][7]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][7]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][7]_i_4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][7]_i_4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][7]_i_4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tfcnt][7]_i_4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_14_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_14_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_14_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_14_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][13]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_14_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_14_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_14_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_14_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][17]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_17_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_17_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_17_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_17_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][1]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_14_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_14_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_14_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_14_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][21]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_14_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_14_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_14_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_14_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][25]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][29]_i_11_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][29]_i_11_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][29]_i_11_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][29]_i_11_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][29]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][29]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][29]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][29]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_14_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_14_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_14_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_14_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][5]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_14_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_14_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_14_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_14_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][addr][9]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[tmsto][write]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[txlength][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[txlength][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rst;

  assign \ahbmo[haddr] [31:1] = \^ahbmo[haddr] [31:1];
  assign \ahbmo[haddr] [0] = etho;
  assign \ahbmo[hburst] [2] = etho;
  assign \ahbmo[hburst] [1] = etho;
  assign \ahbmo[hburst] [0] = apbo;
  assign \ahbmo[hconfig][0] [31] = etho;
  assign \ahbmo[hconfig][0] [30] = etho;
  assign \ahbmo[hconfig][0] [29] = etho;
  assign \ahbmo[hconfig][0] [28] = etho;
  assign \ahbmo[hconfig][0] [27] = etho;
  assign \ahbmo[hconfig][0] [26] = etho;
  assign \ahbmo[hconfig][0] [25] = etho;
  assign \ahbmo[hconfig][0] [24] = apbo;
  assign \ahbmo[hconfig][0] [23] = etho;
  assign \ahbmo[hconfig][0] [22] = etho;
  assign \ahbmo[hconfig][0] [21] = etho;
  assign \ahbmo[hconfig][0] [20] = etho;
  assign \ahbmo[hconfig][0] [19] = etho;
  assign \ahbmo[hconfig][0] [18] = etho;
  assign \ahbmo[hconfig][0] [17] = etho;
  assign \ahbmo[hconfig][0] [16] = apbo;
  assign \ahbmo[hconfig][0] [15] = apbo;
  assign \ahbmo[hconfig][0] [14] = apbo;
  assign \ahbmo[hconfig][0] [13] = etho;
  assign \ahbmo[hconfig][0] [12] = apbo;
  assign \ahbmo[hconfig][0] [11] = etho;
  assign \ahbmo[hconfig][0] [10] = etho;
  assign \ahbmo[hconfig][0] [9] = etho;
  assign \ahbmo[hconfig][0] [8] = etho;
  assign \ahbmo[hconfig][0] [7] = etho;
  assign \ahbmo[hconfig][0] [6] = etho;
  assign \ahbmo[hconfig][0] [5] = etho;
  assign \ahbmo[hconfig][0] [4] = etho;
  assign \ahbmo[hconfig][0] [3] = etho;
  assign \ahbmo[hconfig][0] [2] = etho;
  assign \ahbmo[hconfig][0] [1] = etho;
  assign \ahbmo[hconfig][0] [0] = etho;
  assign \ahbmo[hconfig][1] [31] = etho;
  assign \ahbmo[hconfig][1] [30] = etho;
  assign \ahbmo[hconfig][1] [29] = etho;
  assign \ahbmo[hconfig][1] [28] = etho;
  assign \ahbmo[hconfig][1] [27] = etho;
  assign \ahbmo[hconfig][1] [26] = etho;
  assign \ahbmo[hconfig][1] [25] = etho;
  assign \ahbmo[hconfig][1] [24] = etho;
  assign \ahbmo[hconfig][1] [23] = etho;
  assign \ahbmo[hconfig][1] [22] = etho;
  assign \ahbmo[hconfig][1] [21] = etho;
  assign \ahbmo[hconfig][1] [20] = etho;
  assign \ahbmo[hconfig][1] [19] = etho;
  assign \ahbmo[hconfig][1] [18] = etho;
  assign \ahbmo[hconfig][1] [17] = etho;
  assign \ahbmo[hconfig][1] [16] = etho;
  assign \ahbmo[hconfig][1] [15] = etho;
  assign \ahbmo[hconfig][1] [14] = etho;
  assign \ahbmo[hconfig][1] [13] = etho;
  assign \ahbmo[hconfig][1] [12] = etho;
  assign \ahbmo[hconfig][1] [11] = etho;
  assign \ahbmo[hconfig][1] [10] = etho;
  assign \ahbmo[hconfig][1] [9] = etho;
  assign \ahbmo[hconfig][1] [8] = etho;
  assign \ahbmo[hconfig][1] [7] = etho;
  assign \ahbmo[hconfig][1] [6] = etho;
  assign \ahbmo[hconfig][1] [5] = etho;
  assign \ahbmo[hconfig][1] [4] = etho;
  assign \ahbmo[hconfig][1] [3] = etho;
  assign \ahbmo[hconfig][1] [2] = etho;
  assign \ahbmo[hconfig][1] [1] = etho;
  assign \ahbmo[hconfig][1] [0] = etho;
  assign \ahbmo[hconfig][2] [31] = etho;
  assign \ahbmo[hconfig][2] [30] = etho;
  assign \ahbmo[hconfig][2] [29] = etho;
  assign \ahbmo[hconfig][2] [28] = etho;
  assign \ahbmo[hconfig][2] [27] = etho;
  assign \ahbmo[hconfig][2] [26] = etho;
  assign \ahbmo[hconfig][2] [25] = etho;
  assign \ahbmo[hconfig][2] [24] = etho;
  assign \ahbmo[hconfig][2] [23] = etho;
  assign \ahbmo[hconfig][2] [22] = etho;
  assign \ahbmo[hconfig][2] [21] = etho;
  assign \ahbmo[hconfig][2] [20] = etho;
  assign \ahbmo[hconfig][2] [19] = etho;
  assign \ahbmo[hconfig][2] [18] = etho;
  assign \ahbmo[hconfig][2] [17] = etho;
  assign \ahbmo[hconfig][2] [16] = etho;
  assign \ahbmo[hconfig][2] [15] = etho;
  assign \ahbmo[hconfig][2] [14] = etho;
  assign \ahbmo[hconfig][2] [13] = etho;
  assign \ahbmo[hconfig][2] [12] = etho;
  assign \ahbmo[hconfig][2] [11] = etho;
  assign \ahbmo[hconfig][2] [10] = etho;
  assign \ahbmo[hconfig][2] [9] = etho;
  assign \ahbmo[hconfig][2] [8] = etho;
  assign \ahbmo[hconfig][2] [7] = etho;
  assign \ahbmo[hconfig][2] [6] = etho;
  assign \ahbmo[hconfig][2] [5] = etho;
  assign \ahbmo[hconfig][2] [4] = etho;
  assign \ahbmo[hconfig][2] [3] = etho;
  assign \ahbmo[hconfig][2] [2] = etho;
  assign \ahbmo[hconfig][2] [1] = etho;
  assign \ahbmo[hconfig][2] [0] = etho;
  assign \ahbmo[hconfig][3] [31] = etho;
  assign \ahbmo[hconfig][3] [30] = etho;
  assign \ahbmo[hconfig][3] [29] = etho;
  assign \ahbmo[hconfig][3] [28] = etho;
  assign \ahbmo[hconfig][3] [27] = etho;
  assign \ahbmo[hconfig][3] [26] = etho;
  assign \ahbmo[hconfig][3] [25] = etho;
  assign \ahbmo[hconfig][3] [24] = etho;
  assign \ahbmo[hconfig][3] [23] = etho;
  assign \ahbmo[hconfig][3] [22] = etho;
  assign \ahbmo[hconfig][3] [21] = etho;
  assign \ahbmo[hconfig][3] [20] = etho;
  assign \ahbmo[hconfig][3] [19] = etho;
  assign \ahbmo[hconfig][3] [18] = etho;
  assign \ahbmo[hconfig][3] [17] = etho;
  assign \ahbmo[hconfig][3] [16] = etho;
  assign \ahbmo[hconfig][3] [15] = etho;
  assign \ahbmo[hconfig][3] [14] = etho;
  assign \ahbmo[hconfig][3] [13] = etho;
  assign \ahbmo[hconfig][3] [12] = etho;
  assign \ahbmo[hconfig][3] [11] = etho;
  assign \ahbmo[hconfig][3] [10] = etho;
  assign \ahbmo[hconfig][3] [9] = etho;
  assign \ahbmo[hconfig][3] [8] = etho;
  assign \ahbmo[hconfig][3] [7] = etho;
  assign \ahbmo[hconfig][3] [6] = etho;
  assign \ahbmo[hconfig][3] [5] = etho;
  assign \ahbmo[hconfig][3] [4] = etho;
  assign \ahbmo[hconfig][3] [3] = etho;
  assign \ahbmo[hconfig][3] [2] = etho;
  assign \ahbmo[hconfig][3] [1] = etho;
  assign \ahbmo[hconfig][3] [0] = etho;
  assign \ahbmo[hconfig][4] [31] = etho;
  assign \ahbmo[hconfig][4] [30] = etho;
  assign \ahbmo[hconfig][4] [29] = etho;
  assign \ahbmo[hconfig][4] [28] = etho;
  assign \ahbmo[hconfig][4] [27] = etho;
  assign \ahbmo[hconfig][4] [26] = etho;
  assign \ahbmo[hconfig][4] [25] = etho;
  assign \ahbmo[hconfig][4] [24] = etho;
  assign \ahbmo[hconfig][4] [23] = etho;
  assign \ahbmo[hconfig][4] [22] = etho;
  assign \ahbmo[hconfig][4] [21] = etho;
  assign \ahbmo[hconfig][4] [20] = etho;
  assign \ahbmo[hconfig][4] [19] = etho;
  assign \ahbmo[hconfig][4] [18] = etho;
  assign \ahbmo[hconfig][4] [17] = etho;
  assign \ahbmo[hconfig][4] [16] = etho;
  assign \ahbmo[hconfig][4] [15] = etho;
  assign \ahbmo[hconfig][4] [14] = etho;
  assign \ahbmo[hconfig][4] [13] = etho;
  assign \ahbmo[hconfig][4] [12] = etho;
  assign \ahbmo[hconfig][4] [11] = etho;
  assign \ahbmo[hconfig][4] [10] = etho;
  assign \ahbmo[hconfig][4] [9] = etho;
  assign \ahbmo[hconfig][4] [8] = etho;
  assign \ahbmo[hconfig][4] [7] = etho;
  assign \ahbmo[hconfig][4] [6] = etho;
  assign \ahbmo[hconfig][4] [5] = etho;
  assign \ahbmo[hconfig][4] [4] = etho;
  assign \ahbmo[hconfig][4] [3] = etho;
  assign \ahbmo[hconfig][4] [2] = etho;
  assign \ahbmo[hconfig][4] [1] = etho;
  assign \ahbmo[hconfig][4] [0] = etho;
  assign \ahbmo[hconfig][5] [31] = etho;
  assign \ahbmo[hconfig][5] [30] = etho;
  assign \ahbmo[hconfig][5] [29] = etho;
  assign \ahbmo[hconfig][5] [28] = etho;
  assign \ahbmo[hconfig][5] [27] = etho;
  assign \ahbmo[hconfig][5] [26] = etho;
  assign \ahbmo[hconfig][5] [25] = etho;
  assign \ahbmo[hconfig][5] [24] = etho;
  assign \ahbmo[hconfig][5] [23] = etho;
  assign \ahbmo[hconfig][5] [22] = etho;
  assign \ahbmo[hconfig][5] [21] = etho;
  assign \ahbmo[hconfig][5] [20] = etho;
  assign \ahbmo[hconfig][5] [19] = etho;
  assign \ahbmo[hconfig][5] [18] = etho;
  assign \ahbmo[hconfig][5] [17] = etho;
  assign \ahbmo[hconfig][5] [16] = etho;
  assign \ahbmo[hconfig][5] [15] = etho;
  assign \ahbmo[hconfig][5] [14] = etho;
  assign \ahbmo[hconfig][5] [13] = etho;
  assign \ahbmo[hconfig][5] [12] = etho;
  assign \ahbmo[hconfig][5] [11] = etho;
  assign \ahbmo[hconfig][5] [10] = etho;
  assign \ahbmo[hconfig][5] [9] = etho;
  assign \ahbmo[hconfig][5] [8] = etho;
  assign \ahbmo[hconfig][5] [7] = etho;
  assign \ahbmo[hconfig][5] [6] = etho;
  assign \ahbmo[hconfig][5] [5] = etho;
  assign \ahbmo[hconfig][5] [4] = etho;
  assign \ahbmo[hconfig][5] [3] = etho;
  assign \ahbmo[hconfig][5] [2] = etho;
  assign \ahbmo[hconfig][5] [1] = etho;
  assign \ahbmo[hconfig][5] [0] = etho;
  assign \ahbmo[hconfig][6] [31] = etho;
  assign \ahbmo[hconfig][6] [30] = etho;
  assign \ahbmo[hconfig][6] [29] = etho;
  assign \ahbmo[hconfig][6] [28] = etho;
  assign \ahbmo[hconfig][6] [27] = etho;
  assign \ahbmo[hconfig][6] [26] = etho;
  assign \ahbmo[hconfig][6] [25] = etho;
  assign \ahbmo[hconfig][6] [24] = etho;
  assign \ahbmo[hconfig][6] [23] = etho;
  assign \ahbmo[hconfig][6] [22] = etho;
  assign \ahbmo[hconfig][6] [21] = etho;
  assign \ahbmo[hconfig][6] [20] = etho;
  assign \ahbmo[hconfig][6] [19] = etho;
  assign \ahbmo[hconfig][6] [18] = etho;
  assign \ahbmo[hconfig][6] [17] = etho;
  assign \ahbmo[hconfig][6] [16] = etho;
  assign \ahbmo[hconfig][6] [15] = etho;
  assign \ahbmo[hconfig][6] [14] = etho;
  assign \ahbmo[hconfig][6] [13] = etho;
  assign \ahbmo[hconfig][6] [12] = etho;
  assign \ahbmo[hconfig][6] [11] = etho;
  assign \ahbmo[hconfig][6] [10] = etho;
  assign \ahbmo[hconfig][6] [9] = etho;
  assign \ahbmo[hconfig][6] [8] = etho;
  assign \ahbmo[hconfig][6] [7] = etho;
  assign \ahbmo[hconfig][6] [6] = etho;
  assign \ahbmo[hconfig][6] [5] = etho;
  assign \ahbmo[hconfig][6] [4] = etho;
  assign \ahbmo[hconfig][6] [3] = etho;
  assign \ahbmo[hconfig][6] [2] = etho;
  assign \ahbmo[hconfig][6] [1] = etho;
  assign \ahbmo[hconfig][6] [0] = etho;
  assign \ahbmo[hconfig][7] [31] = etho;
  assign \ahbmo[hconfig][7] [30] = etho;
  assign \ahbmo[hconfig][7] [29] = etho;
  assign \ahbmo[hconfig][7] [28] = etho;
  assign \ahbmo[hconfig][7] [27] = etho;
  assign \ahbmo[hconfig][7] [26] = etho;
  assign \ahbmo[hconfig][7] [25] = etho;
  assign \ahbmo[hconfig][7] [24] = etho;
  assign \ahbmo[hconfig][7] [23] = etho;
  assign \ahbmo[hconfig][7] [22] = etho;
  assign \ahbmo[hconfig][7] [21] = etho;
  assign \ahbmo[hconfig][7] [20] = etho;
  assign \ahbmo[hconfig][7] [19] = etho;
  assign \ahbmo[hconfig][7] [18] = etho;
  assign \ahbmo[hconfig][7] [17] = etho;
  assign \ahbmo[hconfig][7] [16] = etho;
  assign \ahbmo[hconfig][7] [15] = etho;
  assign \ahbmo[hconfig][7] [14] = etho;
  assign \ahbmo[hconfig][7] [13] = etho;
  assign \ahbmo[hconfig][7] [12] = etho;
  assign \ahbmo[hconfig][7] [11] = etho;
  assign \ahbmo[hconfig][7] [10] = etho;
  assign \ahbmo[hconfig][7] [9] = etho;
  assign \ahbmo[hconfig][7] [8] = etho;
  assign \ahbmo[hconfig][7] [7] = etho;
  assign \ahbmo[hconfig][7] [6] = etho;
  assign \ahbmo[hconfig][7] [5] = etho;
  assign \ahbmo[hconfig][7] [4] = etho;
  assign \ahbmo[hconfig][7] [3] = etho;
  assign \ahbmo[hconfig][7] [2] = etho;
  assign \ahbmo[hconfig][7] [1] = etho;
  assign \ahbmo[hconfig][7] [0] = etho;
  assign \ahbmo[hindex] [3] = etho;
  assign \ahbmo[hindex] [2] = apbo;
  assign \ahbmo[hindex] [1] = apbo;
  assign \ahbmo[hindex] [0] = etho;
  assign \ahbmo[hirq] [31] = etho;
  assign \ahbmo[hirq] [30] = etho;
  assign \ahbmo[hirq] [29] = etho;
  assign \ahbmo[hirq] [28] = etho;
  assign \ahbmo[hirq] [27] = etho;
  assign \ahbmo[hirq] [26] = etho;
  assign \ahbmo[hirq] [25] = etho;
  assign \ahbmo[hirq] [24] = etho;
  assign \ahbmo[hirq] [23] = etho;
  assign \ahbmo[hirq] [22] = etho;
  assign \ahbmo[hirq] [21] = etho;
  assign \ahbmo[hirq] [20] = etho;
  assign \ahbmo[hirq] [19] = etho;
  assign \ahbmo[hirq] [18] = etho;
  assign \ahbmo[hirq] [17] = etho;
  assign \ahbmo[hirq] [16] = etho;
  assign \ahbmo[hirq] [15] = etho;
  assign \ahbmo[hirq] [14] = etho;
  assign \ahbmo[hirq] [13] = etho;
  assign \ahbmo[hirq] [12] = etho;
  assign \ahbmo[hirq] [11] = etho;
  assign \ahbmo[hirq] [10] = etho;
  assign \ahbmo[hirq] [9] = etho;
  assign \ahbmo[hirq] [8] = etho;
  assign \ahbmo[hirq] [7] = etho;
  assign \ahbmo[hirq] [6] = etho;
  assign \ahbmo[hirq] [5] = etho;
  assign \ahbmo[hirq] [4] = etho;
  assign \ahbmo[hirq] [3] = etho;
  assign \ahbmo[hirq] [2] = etho;
  assign \ahbmo[hirq] [1] = etho;
  assign \ahbmo[hirq] [0] = etho;
  assign \ahbmo[hlock]  = etho;
  assign \ahbmo[hprot] [3] = etho;
  assign \ahbmo[hprot] [2] = etho;
  assign \ahbmo[hprot] [1] = apbo;
  assign \ahbmo[hprot] [0] = apbo;
  assign \ahbmo[hsize] [2] = etho;
  assign \ahbmo[hsize] [1] = apbo;
  assign \ahbmo[hsize] [0] = etho;
  assign \apbo[pconfig][0] [31] = etho;
  assign \apbo[pconfig][0] [30] = etho;
  assign \apbo[pconfig][0] [29] = etho;
  assign \apbo[pconfig][0] [28] = etho;
  assign \apbo[pconfig][0] [27] = etho;
  assign \apbo[pconfig][0] [26] = etho;
  assign \apbo[pconfig][0] [25] = etho;
  assign \apbo[pconfig][0] [24] = apbo;
  assign \apbo[pconfig][0] [23] = etho;
  assign \apbo[pconfig][0] [22] = etho;
  assign \apbo[pconfig][0] [21] = etho;
  assign \apbo[pconfig][0] [20] = etho;
  assign \apbo[pconfig][0] [19] = etho;
  assign \apbo[pconfig][0] [18] = etho;
  assign \apbo[pconfig][0] [17] = etho;
  assign \apbo[pconfig][0] [16] = apbo;
  assign \apbo[pconfig][0] [15] = apbo;
  assign \apbo[pconfig][0] [14] = apbo;
  assign \apbo[pconfig][0] [13] = etho;
  assign \apbo[pconfig][0] [12] = apbo;
  assign \apbo[pconfig][0] [11] = etho;
  assign \apbo[pconfig][0] [10] = etho;
  assign \apbo[pconfig][0] [9] = etho;
  assign \apbo[pconfig][0] [8] = etho;
  assign \apbo[pconfig][0] [7] = etho;
  assign \apbo[pconfig][0] [6] = etho;
  assign \apbo[pconfig][0] [5] = etho;
  assign \apbo[pconfig][0] [4] = etho;
  assign \apbo[pconfig][0] [3] = apbo;
  assign \apbo[pconfig][0] [2] = apbo;
  assign \apbo[pconfig][0] [1] = etho;
  assign \apbo[pconfig][0] [0] = etho;
  assign \apbo[pconfig][1] [31] = etho;
  assign \apbo[pconfig][1] [30] = etho;
  assign \apbo[pconfig][1] [29] = etho;
  assign \apbo[pconfig][1] [28] = etho;
  assign \apbo[pconfig][1] [27] = etho;
  assign \apbo[pconfig][1] [26] = etho;
  assign \apbo[pconfig][1] [25] = etho;
  assign \apbo[pconfig][1] [24] = etho;
  assign \apbo[pconfig][1] [23] = apbo;
  assign \apbo[pconfig][1] [22] = apbo;
  assign \apbo[pconfig][1] [21] = apbo;
  assign \apbo[pconfig][1] [20] = apbo;
  assign \apbo[pconfig][1] [19] = etho;
  assign \apbo[pconfig][1] [18] = etho;
  assign \apbo[pconfig][1] [17] = etho;
  assign \apbo[pconfig][1] [16] = etho;
  assign \apbo[pconfig][1] [15] = apbo;
  assign \apbo[pconfig][1] [14] = apbo;
  assign \apbo[pconfig][1] [13] = apbo;
  assign \apbo[pconfig][1] [12] = apbo;
  assign \apbo[pconfig][1] [11] = apbo;
  assign \apbo[pconfig][1] [10] = apbo;
  assign \apbo[pconfig][1] [9] = apbo;
  assign \apbo[pconfig][1] [8] = apbo;
  assign \apbo[pconfig][1] [7] = apbo;
  assign \apbo[pconfig][1] [6] = apbo;
  assign \apbo[pconfig][1] [5] = apbo;
  assign \apbo[pconfig][1] [4] = apbo;
  assign \apbo[pconfig][1] [3] = etho;
  assign \apbo[pconfig][1] [2] = etho;
  assign \apbo[pconfig][1] [1] = etho;
  assign \apbo[pconfig][1] [0] = apbo;
  assign \apbo[pindex] [3] = apbo;
  assign \apbo[pindex] [2] = apbo;
  assign \apbo[pindex] [1] = apbo;
  assign \apbo[pindex] [0] = apbo;
  assign \apbo[pirq] [31] = etho;
  assign \apbo[pirq] [30] = etho;
  assign \apbo[pirq] [29] = etho;
  assign \apbo[pirq] [28] = etho;
  assign \apbo[pirq] [27] = etho;
  assign \apbo[pirq] [26] = etho;
  assign \apbo[pirq] [25] = etho;
  assign \apbo[pirq] [24] = etho;
  assign \apbo[pirq] [23] = etho;
  assign \apbo[pirq] [22] = etho;
  assign \apbo[pirq] [21] = etho;
  assign \apbo[pirq] [20] = etho;
  assign \apbo[pirq] [19] = etho;
  assign \apbo[pirq] [18] = etho;
  assign \apbo[pirq] [17] = etho;
  assign \apbo[pirq] [16] = etho;
  assign \apbo[pirq] [15] = etho;
  assign \apbo[pirq] [14] = etho;
  assign \apbo[pirq] [13] = etho;
  assign \apbo[pirq] [12] = \^apbo[pirq] [12];
  assign \apbo[pirq] [11] = etho;
  assign \apbo[pirq] [10] = etho;
  assign \apbo[pirq] [9] = etho;
  assign \apbo[pirq] [8] = etho;
  assign \apbo[pirq] [7] = etho;
  assign \apbo[pirq] [6] = etho;
  assign \apbo[pirq] [5] = etho;
  assign \apbo[pirq] [4] = etho;
  assign \apbo[pirq] [3] = etho;
  assign \apbo[pirq] [2] = etho;
  assign \apbo[pirq] [1] = etho;
  assign \apbo[pirq] [0] = etho;
  assign \etho[gbit]  = etho;
  assign \etho[tx_clk]  = etho;
  assign \etho[tx_er]  = etho;
  assign \etho[txd] [7] = etho;
  assign \etho[txd] [6] = etho;
  assign \etho[txd] [5] = etho;
  assign \etho[txd] [4] = etho;
  assign \etho[txd] [3:0] = \^etho[txd] [3:0];
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0455AAAA)) 
    \FSM_sequential_gmiimode0.r[def_state][0]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/frame_waiting ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [2]),
        .I4(\FSM_sequential_gmiimode0.r[def_state][2]_i_3_n_0 ),
        .O(\FSM_sequential_gmiimode0.r ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000060)) 
    \FSM_sequential_gmiimode0.r[def_state][0]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[deferring_n_0_] ),
        .I3(\gmiimode0.r[start][1]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/frame_waiting ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h06AA)) 
    \FSM_sequential_gmiimode0.r[def_state][1]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [2]),
        .I3(\FSM_sequential_gmiimode0.r[def_state][2]_i_3_n_0 ),
        .O(\FSM_sequential_gmiimode0.r[def_state][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \FSM_sequential_gmiimode0.r[def_state][2]_i_1 
       (.I0(\FSM_sequential_gmiimode0.r[def_state][2]_i_2_n_0 ),
        .I1(\FSM_sequential_gmiimode0.r[def_state][2]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [2]),
        .O(\FSM_sequential_gmiimode0.r[def_state][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00204020)) 
    \FSM_sequential_gmiimode0.r[def_state][2]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/frame_waiting ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in38_in ),
        .O(\FSM_sequential_gmiimode0.r[def_state][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBFBFBFB0F00FFF0)) 
    \FSM_sequential_gmiimode0.r[def_state][2]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/frame_waiting ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .I3(\FSM_sequential_gmiimode0.r[def_state][2]_i_4_n_0 ),
        .I4(\gmiimode0.r[ifg_cycls][7]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [2]),
        .O(\FSM_sequential_gmiimode0.r[def_state][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6562626265626562)) 
    \FSM_sequential_gmiimode0.r[def_state][2]_i_4 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[transmitting]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in38_in ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/rin ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_prev_n_0_] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_act]__1 ),
        .O(\FSM_sequential_gmiimode0.r[def_state][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1777155517771455)) 
    \FSM_sequential_gmiimode0.r[main_state][0]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_31_out ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_28_out ),
        .O(\FSM_sequential_gmiimode0.r[main_state][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h82)) 
    \FSM_sequential_gmiimode0.r[main_state][0]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txvalid_n_0_] ),
        .I1(\m100.u0/ethc0/txo[read] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[read_ack] ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/p_28_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF62426260)) 
    \FSM_sequential_gmiimode0.r[main_state][1]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\FSM_sequential_gmiimode0.r[main_state][1]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\FSM_sequential_gmiimode0.r[main_state][1]_i_3_n_0 ),
        .O(\FSM_sequential_gmiimode0.r[main_state][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \FSM_sequential_gmiimode0.r[main_state][1]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .O(\FSM_sequential_gmiimode0.r[main_state][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111101011111000)) 
    \FSM_sequential_gmiimode0.r[main_state][1]_i_3 
       (.I0(\FSM_sequential_gmiimode0.r[main_state][1]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_31_out ),
        .I2(\gmiimode0.r[byte_count][6]_i_2_n_0 ),
        .I3(\FSM_sequential_gmiimode0.r[main_state][1]_i_5_n_0 ),
        .I4(\FSM_sequential_gmiimode0.r[main_state][1]_i_6_n_0 ),
        .I5(\FSM_sequential_gmiimode0.r[main_state][1]_i_7_n_0 ),
        .O(\FSM_sequential_gmiimode0.r[main_state][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4004000000000000)) 
    \FSM_sequential_gmiimode0.r[main_state][1]_i_4 
       (.I0(\gmiimode0.r_reg[tx_en]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txvalid_n_0_] ),
        .I2(\m100.u0/ethc0/txo[read] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[read_ack] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\FSM_sequential_gmiimode0.r[main_state][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000008000000)) 
    \FSM_sequential_gmiimode0.r[main_state][1]_i_5 
       (.I0(\FSM_sequential_gmiimode0.r[main_state][1]_i_8_n_0 ),
        .I1(\FSM_sequential_gmiimode0.r[main_state][1]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .O(\FSM_sequential_gmiimode0.r[main_state][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0332)) 
    \FSM_sequential_gmiimode0.r[main_state][1]_i_6 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .O(\FSM_sequential_gmiimode0.r[main_state][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA00C000)) 
    \FSM_sequential_gmiimode0.r[main_state][1]_i_7 
       (.I0(\gmiimode0.r[cnt][3]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\gmiimode0.r_reg[tx_en]_i_7_n_0 ),
        .O(\FSM_sequential_gmiimode0.r[main_state][1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h04400000)) 
    \FSM_sequential_gmiimode0.r[main_state][1]_i_8 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][6] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][5] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .I3(\gmiimode0.r[byte_count][6]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ),
        .O(\FSM_sequential_gmiimode0.r[main_state][1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000010101)) 
    \FSM_sequential_gmiimode0.r[main_state][1]_i_9 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][9] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][10] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][8] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][6] ),
        .I4(\gmiimode0.r[byte_count][10]_i_6_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][7] ),
        .O(\FSM_sequential_gmiimode0.r[main_state][1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0CAA30AA)) 
    \FSM_sequential_gmiimode0.r[main_state][2]_i_1 
       (.I0(\FSM_sequential_gmiimode0.r[main_state][2]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\FSM_sequential_gmiimode0.r[main_state][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAEAFAAAAAAABA)) 
    \FSM_sequential_gmiimode0.r[main_state][2]_i_2 
       (.I0(\FSM_sequential_gmiimode0.r[main_state][2]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_28_out ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_31_out ),
        .I5(\gmiimode0.r_reg[tx_en]_i_7_n_0 ),
        .O(\FSM_sequential_gmiimode0.r[main_state][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAB22AA22AA22AA22)) 
    \FSM_sequential_gmiimode0.r[main_state][2]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_31_out ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_28_out ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .O(\FSM_sequential_gmiimode0.r[main_state][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAEAEAEAEFFAEAEAE)) 
    \FSM_sequential_gmiimode0.r[main_state][3]_i_1 
       (.I0(\FSM_sequential_gmiimode0.r[main_state][3]_i_3_n_0 ),
        .I1(\FSM_sequential_gmiimode0.r[main_state][3]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\FSM_sequential_gmiimode0.r[main_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5342FFFF53420000)) 
    \FSM_sequential_gmiimode0.r[main_state][3]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_31_out ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I5(\FSM_sequential_gmiimode0.r[main_state][3]_i_6_n_0 ),
        .O(\FSM_sequential_gmiimode0.r[main_state][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000DFFFDFFFDFFF))
    \FSM_sequential_gmiimode0.r[main_state][3]_i_3 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I5(\FSM_sequential_gmiimode0.r[main_state][3]_i_7_n_0 ),
        .O(\FSM_sequential_gmiimode0.r[main_state][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF1FF01000)) 
    \FSM_sequential_gmiimode0.r[main_state][3]_i_4 
       (.I0(\gmiimode0.r[delay_val][9]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/v [9]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I4(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I5(\FSM_sequential_gmiimode0.r[main_state][3]_i_8_n_0 ),
        .O(\FSM_sequential_gmiimode0.r[main_state][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h20002020)) 
    \FSM_sequential_gmiimode0.r[main_state][3]_i_5 
       (.I0(\etho[tx_en] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in38_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/rin ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_prev_n_0_] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_act]__1 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/p_31_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFAAFFAA0A22)) 
    \FSM_sequential_gmiimode0.r[main_state][3]_i_6 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_28_out ),
        .I2(\gmiimode0.r_reg[tx_en]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_31_out ),
        .O(\FSM_sequential_gmiimode0.r[main_state][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F0C0F0CAA0CEACC)) 
    \FSM_sequential_gmiimode0.r[main_state][3]_i_7 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]14_out ),
        .I1(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I4(\FSM_sequential_gmiimode0.r[main_state][3]_i_9_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\FSM_sequential_gmiimode0.r[main_state][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00F800F800FF0000)) 
    \FSM_sequential_gmiimode0.r[main_state][3]_i_8 
       (.I0(\gmiimode0.r[ifg_cycls][8]_i_5_n_0 ),
        .I1(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]14_out ),
        .I3(\gmiimode0.r[tx_en]_i_5_n_0 ),
        .I4(\gmiimode0.r[byte_count][10]_i_4__0_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\FSM_sequential_gmiimode0.r[main_state][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \FSM_sequential_gmiimode0.r[main_state][3]_i_9 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .O(\FSM_sequential_gmiimode0.r[main_state][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB88888BBB8BB88BB)) 
    \FSM_sequential_gmiimode0.r[rx_state][0]_i_1 
       (.I0(\FSM_sequential_gmiimode0.r[rx_state][0]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I5(\FSM_sequential_gmiimode0.r[rx_state][0]_i_3_n_0 ),
        .O(\FSM_sequential_gmiimode0.r[rx_state][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h20003000)) 
    \FSM_sequential_gmiimode0.r[rx_state][0]_i_2 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .O(\FSM_sequential_gmiimode0.r[rx_state][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \FSM_sequential_gmiimode0.r[rx_state][0]_i_3 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [10]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [8]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [7]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [6]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [9]),
        .O(\FSM_sequential_gmiimode0.r[rx_state][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8CCFF)) 
    \FSM_sequential_gmiimode0.r[rx_state][1]_i_2 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\FSM_sequential_gmiimode0.r[rx_state][0]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .O(\FSM_sequential_gmiimode0.r[rx_state][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FFEA)) 
    \FSM_sequential_gmiimode0.r[rx_state][1]_i_3 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .O(\FSM_sequential_gmiimode0.r[rx_state][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30FF3F0430FFFF77)) 
    \FSM_sequential_gmiimode0.r[rx_state][2]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\FSM_sequential_gmiimode0.r[rx_state][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8A88)) 
    \FSM_sequential_gmiimode0.r[rx_state][2]_i_2 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [10]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [9]),
        .I2(\FSM_sequential_gmiimode0.r[rx_state][2]_i_4_n_0 ),
        .I3(\FSM_sequential_gmiimode0.r[rx_state][2]_i_5_n_0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8880)) 
    \FSM_sequential_gmiimode0.r[rx_state][2]_i_3 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dv]__0 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[en]__0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \FSM_sequential_gmiimode0.r[rx_state][2]_i_4 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [5]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [8]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [7]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [6]),
        .O(\FSM_sequential_gmiimode0.r[rx_state][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEAAAAAAA)) 
    \FSM_sequential_gmiimode0.r[rx_state][2]_i_5 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [4]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [3]),
        .O(\FSM_sequential_gmiimode0.r[rx_state][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \FSM_sequential_gmiimode0.r[rx_state][3]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/rxrst ),
        .O(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \FSM_sequential_gmiimode0.r[rx_state][3]_i_2 
       (.I0(\FSM_sequential_gmiimode0.r[rx_state][3]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I2(\FSM_sequential_gmiimode0.r[rx_state][3]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\FSM_sequential_gmiimode0.r[rx_state][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \FSM_sequential_gmiimode0.r[rx_state][3]_i_3 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .O(\FSM_sequential_gmiimode0.r[rx_state][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB888B888B8BBB8)) 
    \FSM_sequential_gmiimode0.r[rx_state][3]_i_4 
       (.I0(\FSM_sequential_gmiimode0.r[rx_state][3]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\gmiimode0.r[sync_start]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I4(\m100.u0/ethc0/rxo[write] ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[write_ack] ),
        .O(\FSM_sequential_gmiimode0.r[rx_state][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3F32FFFF)) 
    \FSM_sequential_gmiimode0.r[rx_state][3]_i_5 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .O(\FSM_sequential_gmiimode0.r[rx_state][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h909F)) 
    \FSM_sequential_gmiimode0.r[rx_state][3]_i_6 
       (.I0(\m100.u0/ethc0/rxo ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[done_ack_n_0_][0] ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .O(\FSM_sequential_gmiimode0.r[rx_state][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \FSM_sequential_gmiimode0.r_reg[rx_state][1]_i_1 
       (.I0(\FSM_sequential_gmiimode0.r[rx_state][1]_i_2_n_0 ),
        .I1(\FSM_sequential_gmiimode0.r[rx_state][1]_i_3_n_0 ),
        .O(\FSM_sequential_gmiimode0.r_reg ),
        .S(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B888B8B8B8B8)) 
    \FSM_sequential_r[edclrstate][0]_i_1 
       (.I0(\FSM_sequential_r[edclrstate][0]_i_2_n_0 ),
        .I1(\FSM_sequential_r[edclrstate][0]_i_3_n_0 ),
        .I2(\FSM_sequential_r[edclrstate][0]_i_4_n_0 ),
        .I3(\FSM_sequential_r[edclrstate][2]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(FSM_sequential_r));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4703440000000000)) 
    \FSM_sequential_r[edclrstate][0]_i_2 
       (.I0(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\FSM_sequential_r[edclrstate][2]_i_11_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\FSM_sequential_r[edclrstate][0]_i_5_n_0 ),
        .O(\FSM_sequential_r[edclrstate][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8A8A8)) 
    \FSM_sequential_r[edclrstate][0]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I4(\FSM_sequential_r[edclrstate][2]_i_11_n_0 ),
        .I5(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\FSM_sequential_r[edclrstate][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h011F)) 
    \FSM_sequential_r[edclrstate][0]_i_4 
       (.I0(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\FSM_sequential_r[edclrstate][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFBEAAAABE)) 
    \FSM_sequential_r[edclrstate][0]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rxdone] ),
        .I3(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I4(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\FSM_sequential_r[edclrstate][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAEEAE)) 
    \FSM_sequential_r[edclrstate][1]_i_1 
       (.I0(\FSM_sequential_r[edclrstate][1]_i_2_n_0 ),
        .I1(\FSM_sequential_r[edclrstate][1]_i_3_n_0 ),
        .I2(\FSM_sequential_r[edclrstate][2]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I4(\FSM_sequential_r[edclrstate][1]_i_4_n_0 ),
        .I5(\FSM_sequential_r[edclrstate][1]_i_5_n_0 ),
        .O(\FSM_sequential_r[edclrstate][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000044440000000C)) 
    \FSM_sequential_r[edclrstate][1]_i_2 
       (.I0(\FSM_sequential_r[edclrstate][2]_i_11_n_0 ),
        .I1(\FSM_sequential_r[edclrstate][1]_i_6_n_0 ),
        .I2(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I3(\m100.u0/ethc0/v[edclrstate]1124_out ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\FSM_sequential_r[edclrstate][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_r[edclrstate][1]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\FSM_sequential_r[edclrstate][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF00FFDFFFFF)) 
    \FSM_sequential_r[edclrstate][1]_i_4 
       (.I0(\FSM_sequential_r[edclrstate][2]_i_8_n_0 ),
        .I1(\FSM_sequential_r[edclrstate][2]_i_9_n_0 ),
        .I2(\FSM_sequential_r[edclrstate][2]_i_10_n_0 ),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\FSM_sequential_r[edclrstate][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0400)) 
    \FSM_sequential_r[edclrstate][1]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\FSM_sequential_r[edclrstate][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_r[edclrstate][1]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\FSM_sequential_r[edclrstate][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAA8AAA8AAA80000)) 
    \FSM_sequential_r[edclrstate][2]_i_1 
       (.I0(\FSM_sequential_r[edclrstate][2]_i_2_n_0 ),
        .I1(\FSM_sequential_r[edclrstate][2]_i_3_n_0 ),
        .I2(\FSM_sequential_r[edclrstate][2]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I4(\FSM_sequential_r[edclrstate][2]_i_6_n_0 ),
        .I5(\FSM_sequential_r[edclrstate][2]_i_7_n_0 ),
        .O(\FSM_sequential_r[edclrstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \FSM_sequential_r[edclrstate][2]_i_10 
       (.I0(\m100.u0/rxwdata [23]),
        .I1(\m100.u0/rxwdata [30]),
        .I2(\m100.u0/rxwdata [26]),
        .I3(\FSM_sequential_r[edclrstate][2]_i_12_n_0 ),
        .I4(\FSM_sequential_r[edclrstate][2]_i_13_n_0 ),
        .O(\FSM_sequential_r[edclrstate][2]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEFEAEAEA)) 
    \FSM_sequential_r[edclrstate][2]_i_11 
       (.I0(\FSM_sequential_r[edclrstate][2]_i_14_n_0 ),
        .I1(\m100.u0/ethc0/rxo[status] [0]),
        .I2(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I3(\FSM_sequential_r[edclrstate][2]_i_15_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[rxstatus_n_0_][0] ),
        .I5(\r[rxstatus][1]_i_1_n_0 ),
        .O(\FSM_sequential_r[edclrstate][2]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \FSM_sequential_r[edclrstate][2]_i_12 
       (.I0(\m100.u0/rxwdata [28]),
        .I1(\m100.u0/rxwdata [21]),
        .I2(\m100.u0/rxwdata [16]),
        .I3(\m100.u0/rxwdata [25]),
        .O(\FSM_sequential_r[edclrstate][2]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \FSM_sequential_r[edclrstate][2]_i_13 
       (.I0(\m100.u0/rxwdata [31]),
        .I1(\m100.u0/rxwdata [24]),
        .I2(\m100.u0/rxwdata [29]),
        .I3(\m100.u0/rxwdata [22]),
        .O(\FSM_sequential_r[edclrstate][2]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFAEEEAAAAAEEE)) 
    \FSM_sequential_r[edclrstate][2]_i_14 
       (.I0(\r[rxstatus][3]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxstatus_n_0_][2] ),
        .I2(\FSM_sequential_r[edclrstate][2]_i_16_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I5(\m100.u0/ethc0/rxo[status] [2]),
        .O(\FSM_sequential_r[edclrstate][2]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \FSM_sequential_r[edclrstate][2]_i_15 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .O(\FSM_sequential_r[edclrstate][2]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_r[edclrstate][2]_i_16 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .O(\FSM_sequential_r[edclrstate][2]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFDF)) 
    \FSM_sequential_r[edclrstate][2]_i_2 
       (.I0(\FSM_sequential_r[edclrstate][2]_i_8_n_0 ),
        .I1(\FSM_sequential_r[edclrstate][2]_i_9_n_0 ),
        .I2(\FSM_sequential_r[edclrstate][2]_i_10_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\FSM_sequential_r[edclrstate][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \FSM_sequential_r[edclrstate][2]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\FSM_sequential_r[edclrstate][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h04FF0404)) 
    \FSM_sequential_r[edclrstate][2]_i_4 
       (.I0(\m100.u0/ethc0/r_reg ),
        .I1(\m100.u0/ethc0/r_reg[abufs_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .I3(\FSM_sequential_r[edclrstate][3]_i_15_n_0 ),
        .I4(\m100.u0/ethc0/v[edclrstate]2126_in ),
        .O(\FSM_sequential_r[edclrstate][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6006)) 
    \FSM_sequential_r[edclrstate][2]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdone] ),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .O(\m100.u0/ethc0/v[rxstatus]1135_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0500000005550450)) 
    \FSM_sequential_r[edclrstate][2]_i_6 
       (.I0(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I1(\m100.u0/ethc0/v[edclrstate]1124_out ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\FSM_sequential_r[edclrstate][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0400)) 
    \FSM_sequential_r[edclrstate][2]_i_7 
       (.I0(\FSM_sequential_r[edclrstate][2]_i_11_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\FSM_sequential_r[edclrstate][2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \FSM_sequential_r[edclrstate][2]_i_8 
       (.I0(\m100.u0/rxwdata [19]),
        .I1(\m100.u0/rxwdata [18]),
        .I2(\m100.u0/rxwdata [17]),
        .I3(\m100.u0/ethc0/r_reg[edclbcast]__0 ),
        .I4(\m100.u0/rxwdata [20]),
        .I5(\m100.u0/rxwdata [27]),
        .O(\FSM_sequential_r[edclrstate][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF7FFF)) 
    \FSM_sequential_r[edclrstate][2]_i_9 
       (.I0(\m100.u0/rxwdata [17]),
        .I1(\m100.u0/rxwdata [18]),
        .I2(\m100.u0/rxwdata [27]),
        .I3(\m100.u0/ethc0/r_reg[edclbcast]__0 ),
        .I4(\m100.u0/rxwdata [19]),
        .I5(\m100.u0/rxwdata [20]),
        .O(\FSM_sequential_r[edclrstate][2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAEFEAEAE)) 
    \FSM_sequential_r[edclrstate][3]_i_1 
       (.I0(\FSM_sequential_r[edclrstate][3]_i_3_n_0 ),
        .I1(\FSM_sequential_r[edclrstate][3]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\FSM_sequential_r[edclrstate][3]_i_5_n_0 ),
        .O(\FSM_sequential_r[edclrstate][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4000)) 
    \FSM_sequential_r[edclrstate][3]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\FSM_sequential_r[edclrstate][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2AAA2AAA00002AAA)) 
    \FSM_sequential_r[edclrstate][3]_i_11 
       (.I0(\FSM_sequential_r[edclrstate][3]_i_14_n_0 ),
        .I1(\FSM_sequential_r[edclrstate][3]_i_20_n_0 ),
        .I2(\FSM_sequential_r[edclrstate][3]_i_21_n_0 ),
        .I3(\r_reg[edclactive]_i_6_n_2 ),
        .I4(\m100.u0/ethc0/v[edclrstate]01_out ),
        .I5(\FSM_sequential_r[edclrstate][3]_i_23_n_0 ),
        .O(\FSM_sequential_r[edclrstate][3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \FSM_sequential_r[edclrstate][3]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/p_6_in [14]),
        .O(\m100.u0/ethc0/v[edclrstate]0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6666F66FF66F6666)) 
    \FSM_sequential_r[edclrstate][3]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I1(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I3(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I4(\m100.u0/ethc0/r_reg[rxdone] ),
        .I5(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\m100.u0/ethc0/v[edclrstate] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55545555)) 
    \FSM_sequential_r[edclrstate][3]_i_14 
       (.I0(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_r[edclrstate][3]_i_15 
       (.I0(\FSM_sequential_r[edclrstate][3]_i_24_n_0 ),
        .I1(\FSM_sequential_r[edclrstate][3]_i_25_n_0 ),
        .O(\FSM_sequential_r[edclrstate][3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \FSM_sequential_r[edclrstate][3]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[abufs_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg ),
        .O(\FSM_sequential_r[edclrstate][3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_r[edclrstate][3]_i_18 
       (.I0(\m100.u0/ethc0/v[edclrstate]2 ),
        .I1(\FSM_sequential_r[edclrstate][3]_i_24_n_0 ),
        .O(\m100.u0/ethc0/v[edclrstate]1124_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_r[edclrstate][3]_i_19 
       (.I0(\FSM_sequential_r[edclrstate][2]_i_10_n_0 ),
        .I1(\FSM_sequential_r[edclrstate][2]_i_8_n_0 ),
        .O(\m100.u0/ethc0/v[edclrstate]1121_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF00EA)) 
    \FSM_sequential_r[edclrstate][3]_i_2 
       (.I0(\FSM_sequential_r[edclrstate][3]_i_6_n_0 ),
        .I1(\FSM_sequential_r[edclrstate][3]_i_7_n_0 ),
        .I2(\FSM_sequential_r[edclrstate][3]_i_8_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I4(\FSM_sequential_r[edclrstate][3]_i_9_n_0 ),
        .I5(\FSM_sequential_r[edclrstate][3]_i_10_n_0 ),
        .O(\FSM_sequential_r[edclrstate][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_r[edclrstate][3]_i_20 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_r[edclrstate][3]_i_21 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFDF)) 
    \FSM_sequential_r[edclrstate][3]_i_23 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \FSM_sequential_r[edclrstate][3]_i_24 
       (.I0(\FSM_sequential_r[edclrstate][3]_i_34_n_0 ),
        .I1(\m100.u0/rxwdata [20]),
        .I2(\m100.u0/rxwdata [19]),
        .I3(\m100.u0/rxwdata [27]),
        .I4(\m100.u0/rxwdata [25]),
        .I5(\FSM_sequential_r[edclrstate][3]_i_35_n_0 ),
        .O(\FSM_sequential_r[edclrstate][3]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    \FSM_sequential_r[edclrstate][3]_i_25 
       (.I0(\FSM_sequential_r[edclrstate][3]_i_36_n_0 ),
        .I1(\m100.u0/rxwdata [13]),
        .I2(\m100.u0/rxwdata [12]),
        .I3(\m100.u0/rxwdata [9]),
        .I4(\m100.u0/rxwdata [7]),
        .I5(\FSM_sequential_r[edclrstate][3]_i_37_n_0 ),
        .O(\FSM_sequential_r[edclrstate][3]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \FSM_sequential_r[edclrstate][3]_i_27 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][47] ),
        .I1(\m100.u0/rxwdata [31]),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][46] ),
        .I3(\m100.u0/rxwdata [30]),
        .O(\FSM_sequential_r[edclrstate][3]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_28 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][45] ),
        .I1(\m100.u0/rxwdata [29]),
        .I2(\m100.u0/rxwdata [27]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][43] ),
        .I4(\m100.u0/rxwdata [28]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][44] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_29 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][42] ),
        .I1(\m100.u0/rxwdata [26]),
        .I2(\m100.u0/rxwdata [24]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][40] ),
        .I4(\m100.u0/rxwdata [25]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][41] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h20202C202C202020)) 
    \FSM_sequential_r[edclrstate][3]_i_3 
       (.I0(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .I5(\m100.u0/ethc0/r_reg[rxdone] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \FSM_sequential_r[edclrstate][3]_i_32 
       (.I0(\m100.u0/ethc0/p_0_in0_in [15]),
        .I1(\m100.u0/rxwdata [15]),
        .O(\FSM_sequential_r[edclrstate][3]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_33 
       (.I0(\m100.u0/ethc0/p_0_in0_in [14]),
        .I1(\m100.u0/rxwdata [14]),
        .I2(\m100.u0/rxwdata [12]),
        .I3(\m100.u0/ethc0/p_0_in0_in [12]),
        .I4(\m100.u0/rxwdata [13]),
        .I5(\m100.u0/ethc0/p_0_in0_in [13]),
        .O(\FSM_sequential_r[edclrstate][3]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \FSM_sequential_r[edclrstate][3]_i_34 
       (.I0(\m100.u0/rxwdata [17]),
        .I1(\m100.u0/rxwdata [18]),
        .I2(\m100.u0/rxwdata [28]),
        .I3(\m100.u0/rxwdata [22]),
        .O(\FSM_sequential_r[edclrstate][3]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    \FSM_sequential_r[edclrstate][3]_i_35 
       (.I0(\m100.u0/rxwdata [24]),
        .I1(\m100.u0/rxwdata [30]),
        .I2(\m100.u0/rxwdata [26]),
        .I3(\m100.u0/rxwdata [29]),
        .I4(\FSM_sequential_r[edclrstate][3]_i_50_n_0 ),
        .O(\FSM_sequential_r[edclrstate][3]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \FSM_sequential_r[edclrstate][3]_i_36 
       (.I0(\m100.u0/rxwdata [15]),
        .I1(\m100.u0/rxwdata [14]),
        .I2(\m100.u0/rxwdata [11]),
        .I3(\m100.u0/rxwdata [0]),
        .O(\FSM_sequential_r[edclrstate][3]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    \FSM_sequential_r[edclrstate][3]_i_37 
       (.I0(\m100.u0/rxwdata [2]),
        .I1(\m100.u0/rxwdata [6]),
        .I2(\m100.u0/rxwdata [5]),
        .I3(\m100.u0/rxwdata [8]),
        .I4(\FSM_sequential_r[edclrstate][3]_i_51_n_0 ),
        .O(\FSM_sequential_r[edclrstate][3]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_39 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][39] ),
        .I1(\m100.u0/rxwdata [23]),
        .I2(\m100.u0/rxwdata [21]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][37] ),
        .I4(\m100.u0/rxwdata [22]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][38] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5FFF0FFFFFFC000C)) 
    \FSM_sequential_r[edclrstate][3]_i_4 
       (.I0(\FSM_sequential_r[edclrstate][3]_i_11_n_0 ),
        .I1(\m100.u0/ethc0/v[edclrstate]0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/v[edclrstate] ),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\FSM_sequential_r[edclrstate][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_40 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][36] ),
        .I1(\m100.u0/rxwdata [20]),
        .I2(\m100.u0/rxwdata [19]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][35] ),
        .I4(\m100.u0/rxwdata [18]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][34] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_41 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][32] ),
        .I1(\m100.u0/rxwdata [16]),
        .I2(\m100.u0/rxwdata [17]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][33] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][31] ),
        .I5(\m100.u0/rxwdata [15]),
        .O(\FSM_sequential_r[edclrstate][3]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_42 
       (.I0(\m100.u0/rxwdata [14]),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][30] ),
        .I2(\m100.u0/rxwdata [12]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][28] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][29] ),
        .I5(\m100.u0/rxwdata [13]),
        .O(\FSM_sequential_r[edclrstate][3]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \FSM_sequential_r[edclrstate][3]_i_44 
       (.I0(\m100.u0/rxwdata [31]),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][15] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_45 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][14] ),
        .I1(\m100.u0/rxwdata [30]),
        .I2(\m100.u0/rxwdata [28]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][12] ),
        .I4(\m100.u0/rxwdata [29]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][13] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_46 
       (.I0(\m100.u0/ethc0/p_0_in0_in [11]),
        .I1(\m100.u0/rxwdata [11]),
        .I2(\m100.u0/rxwdata [9]),
        .I3(\m100.u0/ethc0/p_0_in0_in [9]),
        .I4(\m100.u0/rxwdata [10]),
        .I5(\m100.u0/ethc0/p_0_in0_in [10]),
        .O(\FSM_sequential_r[edclrstate][3]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_47 
       (.I0(\m100.u0/rxwdata [6]),
        .I1(\m100.u0/ethc0/p_0_in0_in [6]),
        .I2(\m100.u0/rxwdata [7]),
        .I3(\m100.u0/ethc0/p_0_in0_in [7]),
        .I4(\m100.u0/ethc0/p_0_in0_in [8]),
        .I5(\m100.u0/rxwdata [8]),
        .O(\FSM_sequential_r[edclrstate][3]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_48 
       (.I0(\m100.u0/ethc0/p_0_in0_in [5]),
        .I1(\m100.u0/rxwdata [5]),
        .I2(\m100.u0/rxwdata [3]),
        .I3(\m100.u0/ethc0/p_0_in0_in [3]),
        .I4(\m100.u0/rxwdata [4]),
        .I5(\m100.u0/ethc0/p_0_in0_in [4]),
        .O(\FSM_sequential_r[edclrstate][3]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_49 
       (.I0(\m100.u0/rxwdata [2]),
        .I1(\m100.u0/ethc0/p_0_in0_in [2]),
        .I2(\m100.u0/rxwdata [0]),
        .I3(\m100.u0/ethc0/p_0_in0_in [0]),
        .I4(\m100.u0/ethc0/p_0_in0_in [1]),
        .I5(\m100.u0/rxwdata [1]),
        .O(\FSM_sequential_r[edclrstate][3]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD3D3D3D3C0D3D3C0)) 
    \FSM_sequential_r[edclrstate][3]_i_5 
       (.I0(\FSM_sequential_r[edclrstate][3]_i_14_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I5(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\FSM_sequential_r[edclrstate][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \FSM_sequential_r[edclrstate][3]_i_50 
       (.I0(\m100.u0/rxwdata [16]),
        .I1(\m100.u0/rxwdata [21]),
        .I2(\m100.u0/rxwdata [31]),
        .I3(\m100.u0/rxwdata [23]),
        .O(\FSM_sequential_r[edclrstate][3]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \FSM_sequential_r[edclrstate][3]_i_51 
       (.I0(\m100.u0/rxwdata [4]),
        .I1(\m100.u0/rxwdata [3]),
        .I2(\m100.u0/rxwdata [10]),
        .I3(\m100.u0/rxwdata [1]),
        .O(\FSM_sequential_r[edclrstate][3]_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_52 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][26] ),
        .I1(\m100.u0/rxwdata [10]),
        .I2(\m100.u0/rxwdata [11]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][27] ),
        .I4(\m100.u0/rxwdata [9]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][25] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_53 
       (.I0(\m100.u0/rxwdata [8]),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][24] ),
        .I2(\m100.u0/rxwdata [6]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][22] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][23] ),
        .I5(\m100.u0/rxwdata [7]),
        .O(\FSM_sequential_r[edclrstate][3]_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_54 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][21] ),
        .I1(\m100.u0/rxwdata [5]),
        .I2(\m100.u0/rxwdata [3]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][19] ),
        .I4(\m100.u0/rxwdata [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][20] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_55 
       (.I0(\m100.u0/rxwdata [0]),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][16] ),
        .I2(\m100.u0/rxwdata [1]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][17] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][18] ),
        .I5(\m100.u0/rxwdata [2]),
        .O(\FSM_sequential_r[edclrstate][3]_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_56 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][11] ),
        .I1(\m100.u0/rxwdata [27]),
        .I2(\m100.u0/rxwdata [25]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][9] ),
        .I4(\m100.u0/rxwdata [26]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][10] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_57 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][8] ),
        .I1(\m100.u0/rxwdata [24]),
        .I2(\m100.u0/rxwdata [23]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][7] ),
        .I4(\m100.u0/rxwdata [22]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][6] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_58 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][4] ),
        .I1(\m100.u0/rxwdata [20]),
        .I2(\m100.u0/rxwdata [21]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][5] ),
        .I4(\m100.u0/rxwdata [19]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][3] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_sequential_r[edclrstate][3]_i_59 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][2] ),
        .I1(\m100.u0/rxwdata [18]),
        .I2(\m100.u0/rxwdata [16]),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][0] ),
        .I4(\m100.u0/rxwdata [17]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][1] ),
        .O(\FSM_sequential_r[edclrstate][3]_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_r[edclrstate][3]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\FSM_sequential_r[edclrstate][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FFF4)) 
    \FSM_sequential_r[edclrstate][3]_i_7 
       (.I0(\FSM_sequential_r[edclrstate][3]_i_15_n_0 ),
        .I1(\m100.u0/ethc0/v[edclrstate]2126_in ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\FSM_sequential_r[edclrstate][3]_i_17_n_0 ),
        .I4(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\FSM_sequential_r[edclrstate][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hDD20)) 
    \FSM_sequential_r[edclrstate][3]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ethc0/v[edclrstate]1124_out ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\FSM_sequential_r[edclrstate][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \FSM_sequential_r[edclrstate][3]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/v[edclrstate]1121_out ),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\FSM_sequential_r[edclrstate][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000DFF)) 
    \FSM_sequential_r[mdio_state][0]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][write]__0 ),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .O(\FSM_sequential_r[mdio_state][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h003F3F20)) 
    \FSM_sequential_r[mdio_state][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][write]__0 ),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .O(\FSM_sequential_r[mdio_state][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0078)) 
    \FSM_sequential_r[mdio_state][2]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .O(\FSM_sequential_r[mdio_state][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h402A)) 
    \FSM_sequential_r[mdio_state][3]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .O(\FSM_sequential_r[mdio_state][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hED00FFFFED000000)) 
    \FSM_sequential_r[mdio_state][3]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I1(\r[cnt][0]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I3(\m100.u0/ethc0/v[mdio_ctrl][write]1 ),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I5(\r[mdioo]_i_9_n_0 ),
        .O(\FSM_sequential_r[mdio_state][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000AAAA2A22)) 
    \FSM_sequential_r[mdio_state][3]_i_4 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][write]1 ),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I2(\FSM_sequential_r[mdio_state][3]_i_5_n_0 ),
        .I3(\FSM_sequential_r[mdio_state][3]_i_6_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I5(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .O(\FSM_sequential_r[mdio_state][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_r[mdio_state][3]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .O(\FSM_sequential_r[mdio_state][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \FSM_sequential_r[mdio_state][3]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .O(\FSM_sequential_r[mdio_state][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h1505F0F0)) 
    \FSM_sequential_r[regaddr][0]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I1(\m100.u0/ethc0/v[regaddr]1 ),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I4(\FSM_sequential_r[regaddr][2]_i_2_n_0 ),
        .O(\FSM_sequential_r[regaddr][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_r[regaddr][0]_i_2 
       (.I0(\m100.u0/ethc0/p_1_in128_in ),
        .I1(\m100.u0/ethc0/r_reg[rstaneg_n_0_] ),
        .O(\m100.u0/ethc0/v[regaddr]1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h40AA)) 
    \FSM_sequential_r[regaddr][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I1(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I3(\FSM_sequential_r[regaddr][2]_i_2_n_0 ),
        .O(\FSM_sequential_r[regaddr][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \FSM_sequential_r[regaddr][2]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\FSM_sequential_r[regaddr][2]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .O(\FSM_sequential_r[regaddr][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000F800000000)) 
    \FSM_sequential_r[regaddr][2]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I1(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I2(\FSM_sequential_r_reg[regaddr][2]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .O(\FSM_sequential_r[regaddr][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00004500)) 
    \FSM_sequential_r[regaddr][2]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][15] ),
        .I1(\m100.u0/ethc0/r_reg[rstaneg_n_0_] ),
        .I2(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][12] ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .O(\FSM_sequential_r[regaddr][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFEFFFEF)) 
    \FSM_sequential_r[regaddr][2]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I1(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/p_1_in128_in ),
        .I4(\m100.u0/ethc0/r_reg[rstaneg_n_0_] ),
        .O(\FSM_sequential_r[regaddr][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \FSM_sequential_r[rxdstate][0]_i_1 
       (.I0(\FSM_sequential_r[rxdstate][0]_i_2_n_0 ),
        .I1(\FSM_sequential_r[rxdstate][2]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .O(\FSM_sequential_r[rxdstate][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0FAF0FA0CFCFCFCF)) 
    \FSM_sequential_r[rxdstate][0]_i_2 
       (.I0(\FSM_sequential_r[rxdstate][0]_i_3_n_0 ),
        .I1(\FSM_sequential_r[rxdstate][2]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[rxden]__0 ),
        .I5(\m100.u0/ethc0/v[rmsto][write] ),
        .O(\FSM_sequential_r[rxdstate][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF0200FFFF7777)) 
    \FSM_sequential_r[rxdstate][0]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I1(\m100.u0/ethc0/p_0_in153_in ),
        .I2(\m100.u0/ethc0/r_reg[gotframe_n_0_] ),
        .I3(\m100.u0/ethc0/v[status][toosmall]2 ),
        .I4(\m100.u0/ethc0/r_reg[edclactive_n_0_] ),
        .I5(\r[status][toosmall]_i_4_n_0 ),
        .O(\FSM_sequential_r[rxdstate][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \FSM_sequential_r[rxdstate][1]_i_1 
       (.I0(\FSM_sequential_r[rxdstate][1]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I2(\FSM_sequential_r[rxdstate][1]_i_3_n_0 ),
        .I3(\FSM_sequential_r[rxdstate][2]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .O(\FSM_sequential_r[rxdstate][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000088883303BBBB)) 
    \FSM_sequential_r[rxdstate][1]_i_2 
       (.I0(\FSM_sequential_r[rxdstate][1]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/p_0_in153_in ),
        .I3(\m100.u0/ethc0/p_1_in4_in ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I5(\m100.u0/ethc0/rmsti ),
        .O(\FSM_sequential_r[rxdstate][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hC8CB)) 
    \FSM_sequential_r[rxdstate][1]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxden]__0 ),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/p_6_in [1]),
        .O(\FSM_sequential_r[rxdstate][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF5F7F7F7F7F7F7F7)) 
    \FSM_sequential_r[rxdstate][1]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I1(\m100.u0/ethc0/p_0_in153_in ),
        .I2(\m100.u0/ethc0/r_reg[edclactive_n_0_] ),
        .I3(\m100.u0/ethc0/r_reg[gotframe_n_0_] ),
        .I4(\r[status][toosmall]_i_4_n_0 ),
        .I5(\m100.u0/ethc0/v[status][toosmall]2 ),
        .O(\FSM_sequential_r[rxdstate][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \FSM_sequential_r[rxdstate][2]_i_1 
       (.I0(\FSM_sequential_r[rxdstate][2]_i_2_n_0 ),
        .I1(\FSM_sequential_r[rxdstate][2]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .O(\FSM_sequential_r[rxdstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30BBCC8830BBCCBB)) 
    \FSM_sequential_r[rxdstate][2]_i_2 
       (.I0(\FSM_sequential_r[rxdstate][2]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I2(\m100.u0/ethc0/rmsti ),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I5(\m100.u0/ethc0/p_6_in [1]),
        .O(\FSM_sequential_r[rxdstate][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \FSM_sequential_r[rxdstate][2]_i_3 
       (.I0(\FSM_sequential_r[rxdstate][2]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\FSM_sequential_r[rxdstate][2]_i_6_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\FSM_sequential_r[rxdstate][2]_i_7_n_0 ),
        .O(\FSM_sequential_r[rxdstate][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4500)) 
    \FSM_sequential_r[rxdstate][2]_i_4 
       (.I0(\m100.u0/ethc0/rmsti ),
        .I1(\m100.u0/ethc0/p_1_in4_in ),
        .I2(\m100.u0/ethc0/p_0_in153_in ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .O(\FSM_sequential_r[rxdstate][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFBF0F0FBFBF0F00)) 
    \FSM_sequential_r[rxdstate][2]_i_5 
       (.I0(\m100.u0/ethc0/p_0_in153_in ),
        .I1(\r_reg[rxcnt][10]_i_8_n_2 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\FSM_sequential_r[rxdstate][2]_i_8_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I5(\m100.u0/ethc0/r_reg[rxburstav]__0 ),
        .O(\FSM_sequential_r[rxdstate][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFCCEECC)) 
    \FSM_sequential_r[rxdstate][2]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/rmsti ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/rmsti[ready] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .O(\FSM_sequential_r[rxdstate][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFAFAFAFFF3FFF30)) 
    \FSM_sequential_r[rxdstate][2]_i_7 
       (.I0(\FSM_sequential_r[rxdstate][2]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxden]__0 ),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\r[erxidle]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/p_6_in [1]),
        .I5(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .O(\FSM_sequential_r[rxdstate][2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFAE)) 
    \FSM_sequential_r[rxdstate][2]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[edclactive_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[addrdone]__0 ),
        .I2(\m100.u0/ethc0/r_reg[addrok_n_0_] ),
        .I3(\m100.u0/ethc0/r_reg[ctrlpkt]__0 ),
        .O(\FSM_sequential_r[rxdstate][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000D000000000000)) 
    \FSM_sequential_r[rxdstate][2]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I1(\ahbmi[hresp] [0]),
        .I2(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I3(\ahbmi[hresp] [1]),
        .I4(\ahbmi[hready] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg ),
        .O(\FSM_sequential_r[rxdstate][2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \FSM_sequential_r_reg[edclrstate][3]_i_16 
       (.CI(FSM_sequential_r_reg[3]),
        .CO({\FSM_sequential_r_reg[edclrstate][3]_i_16_n_0 ,\m100.u0/ethc0/v[edclrstate]2126_in ,\FSM_sequential_r_reg[edclrstate][3]_i_16_n_2 ,\FSM_sequential_r_reg[edclrstate][3]_i_16_n_3 }),
        .CYINIT(etho),
        .DI({etho,apbo,apbo,apbo}),
        .S({etho,\FSM_sequential_r[edclrstate][3]_i_27_n_0 ,\FSM_sequential_r[edclrstate][3]_i_28_n_0 ,\FSM_sequential_r[edclrstate][3]_i_29_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_r_reg[edclrstate][3]_i_22 
       (.CI(\FSM_sequential_r_reg[edclrstate][3]_i_31_n_0 ),
        .CO({\FSM_sequential_r_reg[edclrstate][3]_i_22_n_0 ,\FSM_sequential_r_reg[edclrstate][3]_i_22_n_1 ,\m100.u0/ethc0/v[edclrstate]01_out ,\FSM_sequential_r_reg[edclrstate][3]_i_22_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,apbo,apbo}),
        .S({etho,etho,\FSM_sequential_r[edclrstate][3]_i_32_n_0 ,\FSM_sequential_r[edclrstate][3]_i_33_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \FSM_sequential_r_reg[edclrstate][3]_i_26 
       (.CI(\FSM_sequential_r_reg[edclrstate][3]_i_38_n_0 ),
        .CO(FSM_sequential_r_reg),
        .CYINIT(etho),
        .DI({apbo,apbo,apbo,apbo}),
        .S({\FSM_sequential_r[edclrstate][3]_i_39_n_0 ,\FSM_sequential_r[edclrstate][3]_i_40_n_0 ,\FSM_sequential_r[edclrstate][3]_i_41_n_0 ,\FSM_sequential_r[edclrstate][3]_i_42_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \FSM_sequential_r_reg[edclrstate][3]_i_30 
       (.CI(\FSM_sequential_r_reg[edclrstate][3]_i_43_n_0 ),
        .CO({\FSM_sequential_r_reg[edclrstate][3]_i_30_n_0 ,\FSM_sequential_r_reg[edclrstate][3]_i_30_n_1 ,\m100.u0/ethc0/v[edclrstate]2 ,\FSM_sequential_r_reg[edclrstate][3]_i_30_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,apbo,apbo}),
        .S({etho,etho,\FSM_sequential_r[edclrstate][3]_i_44_n_0 ,\FSM_sequential_r[edclrstate][3]_i_45_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_r_reg[edclrstate][3]_i_31 
       (.CI(etho),
        .CO({\FSM_sequential_r_reg[edclrstate][3]_i_31_n_0 ,\FSM_sequential_r_reg[edclrstate][3]_i_31_n_1 ,\FSM_sequential_r_reg[edclrstate][3]_i_31_n_2 ,\FSM_sequential_r_reg[edclrstate][3]_i_31_n_3 }),
        .CYINIT(etho),
        .DI({apbo,apbo,apbo,apbo}),
        .S({\FSM_sequential_r[edclrstate][3]_i_46_n_0 ,\FSM_sequential_r[edclrstate][3]_i_47_n_0 ,\FSM_sequential_r[edclrstate][3]_i_48_n_0 ,\FSM_sequential_r[edclrstate][3]_i_49_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \FSM_sequential_r_reg[edclrstate][3]_i_38 
       (.CI(etho),
        .CO({\FSM_sequential_r_reg[edclrstate][3]_i_38_n_0 ,\FSM_sequential_r_reg[edclrstate][3]_i_38_n_1 ,\FSM_sequential_r_reg[edclrstate][3]_i_38_n_2 ,\FSM_sequential_r_reg[edclrstate][3]_i_38_n_3 }),
        .CYINIT(etho),
        .DI({apbo,apbo,apbo,apbo}),
        .S({\FSM_sequential_r[edclrstate][3]_i_52_n_0 ,\FSM_sequential_r[edclrstate][3]_i_53_n_0 ,\FSM_sequential_r[edclrstate][3]_i_54_n_0 ,\FSM_sequential_r[edclrstate][3]_i_55_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \FSM_sequential_r_reg[edclrstate][3]_i_43 
       (.CI(etho),
        .CO({\FSM_sequential_r_reg[edclrstate][3]_i_43_n_0 ,\FSM_sequential_r_reg[edclrstate][3]_i_43_n_1 ,\FSM_sequential_r_reg[edclrstate][3]_i_43_n_2 ,\FSM_sequential_r_reg[edclrstate][3]_i_43_n_3 }),
        .CYINIT(etho),
        .DI({apbo,apbo,apbo,apbo}),
        .S({\FSM_sequential_r[edclrstate][3]_i_56_n_0 ,\FSM_sequential_r[edclrstate][3]_i_57_n_0 ,\FSM_sequential_r[edclrstate][3]_i_58_n_0 ,\FSM_sequential_r[edclrstate][3]_i_59_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \FSM_sequential_r_reg[mdio_state][3]_i_1 
       (.I0(\FSM_sequential_r[mdio_state][3]_i_3_n_0 ),
        .I1(\FSM_sequential_r[mdio_state][3]_i_4_n_0 ),
        .O(\FSM_sequential_r_reg[mdio_state][3]_i_1_n_0 ),
        .S(\m100.u0/ethc0/r_reg[mdio_state] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \FSM_sequential_r_reg[regaddr][2]_i_3 
       (.I0(\FSM_sequential_r[regaddr][2]_i_4_n_0 ),
        .I1(\FSM_sequential_r[regaddr][2]_i_5_n_0 ),
        .O(\FSM_sequential_r_reg[regaddr][2]_i_3_n_0 ),
        .S(\m100.u0/ethc0/r_reg[regaddr] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_1
       (.G(GND_2));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(apbo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_1
       (.P(VCC_2));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBAAAFAFABAAABAAA)) 
    \a9.x[0].r0_i_1 
       (.I0(\a9.x[0].r0_i_18_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ethc0/v[writeok]1 ),
        .I3(\a9.x[0].r0_i_19_n_0 ),
        .I4(\r[erxidle]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\m100.u0/ewritem ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \a9.x[0].r0_i_10 
       (.I0(\a9.x[0].r0_i_38_n_0 ),
        .I1(\r[rcntl][6]_i_5_n_0 ),
        .I2(\a9.x[0].r0_i_39__0_n_0 ),
        .I3(\m100.u0/ethc0/swap ),
        .I4(\m100.u0/rxwdata [7]),
        .I5(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_100 
       (.I0(\m100.u0/rxwdata [0]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][32] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][0] ),
        .O(\a9.x ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_101 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][32] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [0]),
        .O(\a9.x[0].r0_i_101_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \a9.x[0].r0_i_101__0 
       (.I0(\m100.u0/ethc0/r_reg[applength]__0 [5]),
        .O(\a9.x[0].r0_i_101__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \a9.x[0].r0_i_103 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/rxwdata [6]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I4(\m100.u0/rxwdata [22]),
        .O(\a9.x[0].r0_i_103_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \a9.x[0].r0_i_104 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/rxwdata [5]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I4(\m100.u0/rxwdata [21]),
        .O(\a9.x[0].r0_i_104_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \a9.x[0].r0_i_105 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/rxwdata [4]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I4(\m100.u0/rxwdata [20]),
        .O(\a9.x[0].r0_i_105_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \a9.x[0].r0_i_107 
       (.I0(\m100.u0/ethc0/r_reg[applength]__0 [4]),
        .O(\a9.x[0].r0_i_107_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \a9.x[0].r0_i_107__0 
       (.I0(\m100.u0/ethc0/r_reg[applength]__0 [2]),
        .O(\a9.x[0].r0_i_107__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \a9.x[0].r0_i_108 
       (.I0(\m100.u0/ethc0/r_reg[applength]__0 [1]),
        .O(\a9.x[0].r0_i_108_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB8BB8888B888)) 
    \a9.x[0].r0_i_10__0 
       (.I0(\m100.u0/rxwdata [23]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_37_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\a9.x[0].r0_i_38__0_n_0 ),
        .O(\m100.u0/datain [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_10__1 
       (.I0(\m100.u0/erdata [23]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [23]),
        .O(\m100.u0/txwdata [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \a9.x[0].r0_i_11 
       (.I0(\a9.x[0].r0_i_40__0_n_0 ),
        .I1(\r[rcntl][6]_i_5_n_0 ),
        .I2(\a9.x[0].r0_i_41__0_n_0 ),
        .I3(\m100.u0/ethc0/swap ),
        .I4(\m100.u0/rxwdata [6]),
        .I5(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \a9.x[0].r0_i_110 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/rxwdata [2]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I4(\m100.u0/rxwdata [18]),
        .O(\a9.x[0].r0_i_110_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \a9.x[0].r0_i_111 
       (.CI(etho),
        .CO({\a9.x[0].r0_i_111_n_0 ,\a9.x[0].r0_i_111_n_1 ,\a9.x[0].r0_i_111_n_2 ,\a9.x[0].r0_i_111_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,\m100.u0/ethc0/r_reg[applength]__0 [1],etho}),
        .O({\a9.x[0].r0_i_111_n_4 ,\a9.x[0].r0_i_111_n_5 ,\a9.x[0].r0_i_111_n_6 ,\a9.x[0].r0_i_111_n_7 }),
        .S({\m100.u0/ethc0/r_reg[applength]__0 [3:2],\a9.x[0].r0_i_114_n_0 ,\m100.u0/ethc0/r_reg[applength]__0 [0]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \a9.x[0].r0_i_114 
       (.I0(\m100.u0/ethc0/r_reg[applength]__0 [1]),
        .O(\a9.x[0].r0_i_114_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB8BB8888B888)) 
    \a9.x[0].r0_i_11__0 
       (.I0(\m100.u0/rxwdata [22]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_39_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\m100.u0/rxwdata [6]),
        .O(\m100.u0/datain [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_11__1 
       (.I0(\m100.u0/erdata [22]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [22]),
        .O(\m100.u0/txwdata [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \a9.x[0].r0_i_12 
       (.I0(\a9.x[0].r0_i_42__0_n_0 ),
        .I1(\r[rcntl][6]_i_5_n_0 ),
        .I2(\a9.x[0].r0_i_43__0_n_0 ),
        .I3(\m100.u0/ethc0/swap ),
        .I4(\m100.u0/rxwdata [5]),
        .I5(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB8BB8888B888)) 
    \a9.x[0].r0_i_12__0 
       (.I0(\m100.u0/rxwdata [21]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_40_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\m100.u0/rxwdata [5]),
        .O(\m100.u0/datain [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_12__1 
       (.I0(\m100.u0/erdata [21]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [21]),
        .O(\m100.u0/txwdata [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \a9.x[0].r0_i_13 
       (.I0(\a9.x[0].r0_i_44__0_n_0 ),
        .I1(\r[rcntl][6]_i_5_n_0 ),
        .I2(\a9.x[0].r0_i_45__0_n_0 ),
        .I3(\m100.u0/ethc0/swap ),
        .I4(\m100.u0/rxwdata [4]),
        .I5(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB8BB8888B888)) 
    \a9.x[0].r0_i_13__0 
       (.I0(\m100.u0/rxwdata [20]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_41_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\m100.u0/rxwdata [4]),
        .O(\m100.u0/datain [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_13__1 
       (.I0(\m100.u0/erdata [20]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [20]),
        .O(\m100.u0/txwdata [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \a9.x[0].r0_i_14 
       (.I0(\a9.x[0].r0_i_46_n_0 ),
        .I1(\r[rcntl][6]_i_5_n_0 ),
        .I2(\a9.x[0].r0_i_47_n_0 ),
        .I3(\m100.u0/ethc0/swap ),
        .I4(\m100.u0/rxwdata [3]),
        .I5(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB8BB8888B888)) 
    \a9.x[0].r0_i_14__0 
       (.I0(\m100.u0/rxwdata [19]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_42_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\m100.u0/rxwdata [3]),
        .O(\m100.u0/datain [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_14__1 
       (.I0(\m100.u0/erdata [19]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [19]),
        .O(\m100.u0/txwdata [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \a9.x[0].r0_i_15 
       (.I0(\a9.x[0].r0_i_48_n_0 ),
        .I1(\r[rcntl][6]_i_5_n_0 ),
        .I2(\a9.x[0].r0_i_49_n_0 ),
        .I3(\m100.u0/ethc0/swap ),
        .I4(\m100.u0/rxwdata [2]),
        .I5(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB8BB8888B888)) 
    \a9.x[0].r0_i_15__0 
       (.I0(\m100.u0/rxwdata [18]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_43_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\m100.u0/rxwdata [2]),
        .O(\m100.u0/datain [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_15__1 
       (.I0(\m100.u0/erdata [18]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [18]),
        .O(\m100.u0/txwdata [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \a9.x[0].r0_i_16 
       (.I0(\a9.x[0].r0_i_50_n_0 ),
        .I1(\r[rcntl][6]_i_5_n_0 ),
        .I2(\a9.x[0].r0_i_51_n_0 ),
        .I3(\m100.u0/ethc0/swap ),
        .I4(\m100.u0/rxwdata [1]),
        .I5(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB8BB8888B888)) 
    \a9.x[0].r0_i_16__0 
       (.I0(\m100.u0/rxwdata [17]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_44_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\m100.u0/rxwdata [1]),
        .O(\m100.u0/datain [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_16__1 
       (.I0(\m100.u0/erdata [17]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [17]),
        .O(\m100.u0/txwdata [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \a9.x[0].r0_i_17 
       (.I0(\a9.x[0].r0_i_52_n_0 ),
        .I1(\r[rcntl][6]_i_5_n_0 ),
        .I2(\a9.x[0].r0_i_53_n_0 ),
        .I3(\m100.u0/ethc0/swap ),
        .I4(\m100.u0/rxwdata [0]),
        .I5(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB8BB8888B888)) 
    \a9.x[0].r0_i_17__0 
       (.I0(\m100.u0/rxwdata [16]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_45_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\m100.u0/rxwdata [0]),
        .O(\m100.u0/datain [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_17__1 
       (.I0(\m100.u0/erdata [16]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [16]),
        .O(\m100.u0/txwdata [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAABFAABFF000C000)) 
    \a9.x[0].r0_i_18 
       (.I0(\a9.x[0].r0_i_54_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/ethc0/v[rcntm]0 ),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\a9.x[0].r0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6666666066666666)) 
    \a9.x[0].r0_i_18__0 
       (.I0(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I1(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\m100.u0/ethc0/veri ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_18__1 
       (.I0(\m100.u0/erdata [15]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [15]),
        .O(\m100.u0/txwdata [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFABA)) 
    \a9.x[0].r0_i_19 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/v[rcntm]0 ),
        .O(\a9.x[0].r0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000005DFA0800)) 
    \a9.x[0].r0_i_19__0 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\m100.u0/ethc0/v[rcntm]0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/ethc0/v[writeok]1 ),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\a9.x[0].r0_i_19__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_19__1 
       (.I0(\m100.u0/erdata [14]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [14]),
        .O(\m100.u0/txwdata [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFA03F0000)) 
    \a9.x[0].r0_i_1__0 
       (.I0(\m100.u0/ethc0/veri ),
        .I1(\r[erxidle]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\r[rcntl][6]_i_5_n_0 ),
        .I5(\a9.x[0].r0_i_19__0_n_0 ),
        .O(\m100.u0/ewritel ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000C004)) 
    \a9.x[0].r0_i_1__1 
       (.I0(\a9.x[0].r0_i_34__1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\m100.u0/txwrite ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FE0E)) 
    \a9.x[0].r0_i_2 
       (.I0(\a9.x[0].r0_i_20__0_n_0 ),
        .I1(\a9.x[0].r0_i_21_n_0 ),
        .I2(\m100.u0/ethc0/swap ),
        .I3(\m100.u0/rxwdata [15]),
        .I4(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDBD0000DDFD0000)) 
    \a9.x[0].r0_i_20 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/rxwdata [15]),
        .I5(\a9.x[0].r0_i_90_n_0 ),
        .O(\a9.x[0].r0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0080008088880080)) 
    \a9.x[0].r0_i_20__0 
       (.I0(\r[rcntl][6]_i_5_n_0 ),
        .I1(\a9.x[0].r0_i_22_n_0 ),
        .I2(\m100.u0/rxwdata [31]),
        .I3(\a9.x[0].r0_i_55_n_0 ),
        .I4(\m100.u0/ethc0/v[writeok]1 ),
        .I5(\a9.x[0].r0_i_56__0_n_0 ),
        .O(\a9.x[0].r0_i_20__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_20__1 
       (.I0(\m100.u0/erdata [13]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [13]),
        .O(\m100.u0/txwdata [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F808F8F8F808F80)) 
    \a9.x[0].r0_i_21 
       (.I0(\m100.u0/ethc0/r_reg[udpsrc_n_0_][15] ),
        .I1(\a9.x[0].r0_i_57__0_n_0 ),
        .I2(\r[rcntl][6]_i_5_n_0 ),
        .I3(\a9.x[0].r0_i_58_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ipcrc_n_0_][15] ),
        .I5(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB8B8FF00B8B800)) 
    \a9.x[0].r0_i_21__0 
       (.I0(\a9.x[0].r0_i_46__0_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\a9.x[0].r0_i_47__0_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I4(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I5(\m100.u0/rxwdata [15]),
        .O(\a9.x[0].r0_i_21__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_21__1 
       (.I0(\m100.u0/erdata [12]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [12]),
        .O(\m100.u0/txwdata [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4080)) 
    \a9.x[0].r0_i_22 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000008080FC00)) 
    \a9.x[0].r0_i_22__0 
       (.I0(\m100.u0/ethc0/swap12_out ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\m100.u0/ethc0/swap ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_22__1 
       (.I0(\m100.u0/erdata [11]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [11]),
        .O(\m100.u0/txwdata [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00080000)) 
    \a9.x[0].r0_i_23 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/ethc0/setmz11_out ),
        .O(\m100.u0/ethc0/setmz ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDBD0000DDFD0000)) 
    \a9.x[0].r0_i_23__0 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/rxwdata [14]),
        .I5(\a9.x[0].r0_i_90_n_0 ),
        .O(\a9.x[0].r0_i_23__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_23__1 
       (.I0(\m100.u0/erdata [10]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [10]),
        .O(\m100.u0/txwdata [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0020002000200000)) 
    \a9.x[0].r0_i_24 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\a9.x[0].r0_i_61__0_n_0 ),
        .I4(\m100.u0/rxwdata [30]),
        .I5(\a9.x[0].r0_i_55_n_0 ),
        .O(\a9.x[0].r0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB8B8FF00B8B800)) 
    \a9.x[0].r0_i_24__0 
       (.I0(\a9.x[0].r0_i_48__0_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\a9.x[0].r0_i_49__0_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I4(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I5(\m100.u0/rxwdata [14]),
        .O(\a9.x[0].r0_i_24__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_24__1 
       (.I0(\m100.u0/erdata [9]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [9]),
        .O(\m100.u0/txwdata [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F808F8F8F808F80)) 
    \a9.x[0].r0_i_25 
       (.I0(\m100.u0/ethc0/r_reg[udpsrc_n_0_][14] ),
        .I1(\a9.x[0].r0_i_57__0_n_0 ),
        .I2(\r[rcntl][6]_i_5_n_0 ),
        .I3(\a9.x[0].r0_i_62_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ipcrc_n_0_][14] ),
        .I5(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDBD0000DDFD0000)) 
    \a9.x[0].r0_i_25__0 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/rxwdata [13]),
        .I5(\a9.x[0].r0_i_90_n_0 ),
        .O(\a9.x[0].r0_i_25__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_25__1 
       (.I0(\m100.u0/erdata [8]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [8]),
        .O(\m100.u0/txwdata [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0020002000200000)) 
    \a9.x[0].r0_i_26 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\a9.x[0].r0_i_63__0_n_0 ),
        .I4(\m100.u0/rxwdata [29]),
        .I5(\a9.x[0].r0_i_55_n_0 ),
        .O(\a9.x[0].r0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB8B8FF00B8B800)) 
    \a9.x[0].r0_i_26__0 
       (.I0(\a9.x[0].r0_i_50__0_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\a9.x[0].r0_i_51__0_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I4(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I5(\m100.u0/rxwdata [13]),
        .O(\a9.x[0].r0_i_26__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_26__1 
       (.I0(\m100.u0/erdata [7]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [7]),
        .O(\m100.u0/txwdata [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F808F8F8F808F80)) 
    \a9.x[0].r0_i_27 
       (.I0(\m100.u0/ethc0/r_reg[udpsrc_n_0_][13] ),
        .I1(\a9.x[0].r0_i_57__0_n_0 ),
        .I2(\r[rcntl][6]_i_5_n_0 ),
        .I3(\a9.x[0].r0_i_64_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ipcrc_n_0_][13] ),
        .I5(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDBD0000DDFD0000)) 
    \a9.x[0].r0_i_27__0 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/rxwdata [12]),
        .I5(\a9.x[0].r0_i_90_n_0 ),
        .O(\a9.x[0].r0_i_27__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_27__1 
       (.I0(\m100.u0/erdata [6]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [6]),
        .O(\m100.u0/txwdata [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0020002000200000)) 
    \a9.x[0].r0_i_28 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\a9.x[0].r0_i_65__0_n_0 ),
        .I4(\m100.u0/rxwdata [28]),
        .I5(\a9.x[0].r0_i_55_n_0 ),
        .O(\a9.x[0].r0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB8B8FF00B8B800)) 
    \a9.x[0].r0_i_28__0 
       (.I0(\a9.x[0].r0_i_52__0_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\a9.x[0].r0_i_53__0_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I4(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I5(\m100.u0/rxwdata [12]),
        .O(\a9.x[0].r0_i_28__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_28__1 
       (.I0(\m100.u0/erdata [5]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [5]),
        .O(\m100.u0/txwdata [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F808F8F8F808F80)) 
    \a9.x[0].r0_i_29 
       (.I0(\m100.u0/ethc0/r_reg[udpsrc_n_0_][12] ),
        .I1(\a9.x[0].r0_i_57__0_n_0 ),
        .I2(\r[rcntl][6]_i_5_n_0 ),
        .I3(\a9.x[0].r0_i_66_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ipcrc_n_0_][12] ),
        .I5(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDBD0000DDFD0000)) 
    \a9.x[0].r0_i_29__0 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/rxwdata [11]),
        .I5(\a9.x[0].r0_i_90_n_0 ),
        .O(\a9.x[0].r0_i_29__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_29__1 
       (.I0(\m100.u0/erdata [4]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [4]),
        .O(\m100.u0/txwdata [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B8B8B8B8B8)) 
    \a9.x[0].r0_i_2__0 
       (.I0(\m100.u0/rxwdata [31]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_20_n_0 ),
        .I3(\a9.x[0].r0_i_21__0_n_0 ),
        .I4(\a9.x[0].r0_i_22_n_0 ),
        .I5(\r[rcntl][6]_i_5_n_0 ),
        .O(\m100.u0/datain [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_2__1 
       (.I0(\m100.u0/erdata [31]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [31]),
        .O(\m100.u0/txwdata [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FE0E)) 
    \a9.x[0].r0_i_3 
       (.I0(\a9.x[0].r0_i_24_n_0 ),
        .I1(\a9.x[0].r0_i_25_n_0 ),
        .I2(\m100.u0/ethc0/swap ),
        .I3(\m100.u0/rxwdata [14]),
        .I4(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0020002000200000)) 
    \a9.x[0].r0_i_30 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\a9.x[0].r0_i_67__0_n_0 ),
        .I4(\m100.u0/rxwdata [27]),
        .I5(\a9.x[0].r0_i_55_n_0 ),
        .O(\a9.x[0].r0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB8B8FF00B8B800)) 
    \a9.x[0].r0_i_30__0 
       (.I0(\a9.x[0].r0_i_54__0_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\a9.x[0].r0_i_55__0_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I4(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I5(\m100.u0/rxwdata [11]),
        .O(\a9.x[0].r0_i_30__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_30__1 
       (.I0(\m100.u0/erdata [3]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [3]),
        .O(\m100.u0/txwdata [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF8C888C8)) 
    \a9.x[0].r0_i_31 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\m100.u0/rxwdata [10]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\a9.x[0].r0_i_56_n_0 ),
        .I5(\a9.x[0].r0_i_57_n_0 ),
        .O(\a9.x[0].r0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F808F8F8F808F80)) 
    \a9.x[0].r0_i_31__0 
       (.I0(\m100.u0/ethc0/r_reg[udpsrc_n_0_][11] ),
        .I1(\a9.x[0].r0_i_57__0_n_0 ),
        .I2(\r[rcntl][6]_i_5_n_0 ),
        .I3(\a9.x[0].r0_i_68_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ipcrc_n_0_][11] ),
        .I5(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_31__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_31__1 
       (.I0(\m100.u0/erdata [2]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [2]),
        .O(\m100.u0/txwdata [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFF0F0E2E20000)) 
    \a9.x[0].r0_i_32 
       (.I0(\m100.u0/ethc0/r_reg[seq] [8]),
        .I1(\a9.x[0].r0_i_69__0_n_0 ),
        .I2(\m100.u0/rxwdata [26]),
        .I3(\m100.u0/ethc0/r_reg[ipcrc_n_0_][10] ),
        .I4(\a9.x[0].r0_i_70_n_0 ),
        .I5(\a9.x[0].r0_i_71__0_n_0 ),
        .O(\a9.x[0].r0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFDBF0000FFFF0000)) 
    \a9.x[0].r0_i_32__0 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/rxwdata [10]),
        .I5(\a9.x[0].r0_i_90_n_0 ),
        .O(\a9.x[0].r0_i_32__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_32__1 
       (.I0(\m100.u0/erdata [1]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [1]),
        .O(\m100.u0/txwdata [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF8C888C8)) 
    \a9.x[0].r0_i_33 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\m100.u0/rxwdata [9]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\a9.x[0].r0_i_58__0_n_0 ),
        .I5(\a9.x[0].r0_i_59_n_0 ),
        .O(\a9.x[0].r0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \a9.x[0].r0_i_33__0 
       (.I0(\a9.x[0].r0_i_57__0_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[udpsrc_n_0_][10] ),
        .I2(\a9.x[0].r0_i_72_n_0 ),
        .I3(\a9.x[0].r0_i_73__0_n_1 ),
        .I4(\a9.x[0].r0_i_74_n_0 ),
        .I5(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_33__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_33__1 
       (.I0(\m100.u0/erdata [0]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [0]),
        .O(\m100.u0/txwdata [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFF0F0E2E20000)) 
    \a9.x[0].r0_i_34 
       (.I0(\m100.u0/ethc0/r_reg[seq] [7]),
        .I1(\a9.x[0].r0_i_69__0_n_0 ),
        .I2(\m100.u0/rxwdata [25]),
        .I3(\m100.u0/ethc0/r_reg[ipcrc_n_0_][9] ),
        .I4(\a9.x[0].r0_i_70_n_0 ),
        .I5(\a9.x[0].r0_i_71__0_n_0 ),
        .O(\a9.x[0].r0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFDBF0000FFFF0000)) 
    \a9.x[0].r0_i_34__0 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/rxwdata [9]),
        .I5(\a9.x[0].r0_i_90_n_0 ),
        .O(\a9.x[0].r0_i_34__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF4FFFFFFFFFFFFF)) 
    \a9.x[0].r0_i_34__1 
       (.I0(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I1(\ahbmi[hresp] [0]),
        .I2(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I3(\ahbmi[hresp] [1]),
        .I4(\ahbmi[hready] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg ),
        .O(\a9.x[0].r0_i_34__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF8C888C8)) 
    \a9.x[0].r0_i_35 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\m100.u0/rxwdata [8]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\a9.x[0].r0_i_60__0_n_0 ),
        .I5(\a9.x[0].r0_i_61_n_0 ),
        .O(\a9.x[0].r0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAFEAAAA)) 
    \a9.x[0].r0_i_35__0 
       (.I0(\a9.x[0].r0_i_75__0_n_0 ),
        .I1(\a9.x[0].r0_i_55_n_0 ),
        .I2(\m100.u0/rxwdata [25]),
        .I3(\a9.x[0].r0_i_76_n_0 ),
        .I4(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_35__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFF0F0E2E20000)) 
    \a9.x[0].r0_i_36 
       (.I0(\m100.u0/ethc0/r_reg[seq] [6]),
        .I1(\a9.x[0].r0_i_69__0_n_0 ),
        .I2(\m100.u0/rxwdata [24]),
        .I3(\m100.u0/ethc0/r_reg[ipcrc_n_0_][8] ),
        .I4(\a9.x[0].r0_i_70_n_0 ),
        .I5(\a9.x[0].r0_i_71__0_n_0 ),
        .O(\a9.x[0].r0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFDBF0000FFFF0000)) 
    \a9.x[0].r0_i_36__0 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/rxwdata [8]),
        .I5(\a9.x[0].r0_i_90_n_0 ),
        .O(\a9.x[0].r0_i_36__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF8C888C8)) 
    \a9.x[0].r0_i_37 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\m100.u0/rxwdata [7]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\a9.x[0].r0_i_62__0_n_0 ),
        .I5(\a9.x[0].r0_i_63_n_0 ),
        .O(\a9.x[0].r0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \a9.x[0].r0_i_37__0 
       (.I0(\a9.x[0].r0_i_57__0_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[udpsrc_n_0_][8] ),
        .I2(\a9.x[0].r0_i_72_n_0 ),
        .I3(\a9.x[0].r0_i_73__0_n_7 ),
        .I4(\a9.x[0].r0_i_77__0_n_0 ),
        .I5(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_37__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFF0F0E2E20000)) 
    \a9.x[0].r0_i_38 
       (.I0(\m100.u0/ethc0/r_reg[seq] [5]),
        .I1(\a9.x[0].r0_i_69__0_n_0 ),
        .I2(\m100.u0/rxwdata [23]),
        .I3(\m100.u0/ethc0/r_reg[ipcrc_n_0_][7] ),
        .I4(\a9.x[0].r0_i_70_n_0 ),
        .I5(\a9.x[0].r0_i_71__0_n_0 ),
        .O(\a9.x[0].r0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFDBF0000FFFF0000)) 
    \a9.x[0].r0_i_38__0 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/rxwdata [7]),
        .I5(\a9.x[0].r0_i_90_n_0 ),
        .O(\a9.x[0].r0_i_38__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF8C888C8)) 
    \a9.x[0].r0_i_39 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\m100.u0/rxwdata [6]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\a9.x[0].r0_i_64__0_n_0 ),
        .I5(\a9.x[0].r0_i_65_n_0 ),
        .O(\a9.x[0].r0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAFEAAAA)) 
    \a9.x[0].r0_i_39__0 
       (.I0(\a9.x[0].r0_i_78_n_0 ),
        .I1(\a9.x[0].r0_i_55_n_0 ),
        .I2(\m100.u0/rxwdata [23]),
        .I3(\a9.x[0].r0_i_79_n_0 ),
        .I4(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_39__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B8B8B8B8B8)) 
    \a9.x[0].r0_i_3__0 
       (.I0(\m100.u0/rxwdata [30]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_23__0_n_0 ),
        .I3(\a9.x[0].r0_i_24__0_n_0 ),
        .I4(\a9.x[0].r0_i_22_n_0 ),
        .I5(\r[rcntl][6]_i_5_n_0 ),
        .O(\m100.u0/datain [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_3__1 
       (.I0(\m100.u0/erdata [30]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [30]),
        .O(\m100.u0/txwdata [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FE0E)) 
    \a9.x[0].r0_i_4 
       (.I0(\a9.x[0].r0_i_26_n_0 ),
        .I1(\a9.x[0].r0_i_27_n_0 ),
        .I2(\m100.u0/ethc0/swap ),
        .I3(\m100.u0/rxwdata [13]),
        .I4(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF8C888C8)) 
    \a9.x[0].r0_i_40 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\m100.u0/rxwdata [5]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\a9.x[0].r0_i_66__0_n_0 ),
        .I5(\a9.x[0].r0_i_67_n_0 ),
        .O(\a9.x[0].r0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFF0F0E2E20000)) 
    \a9.x[0].r0_i_40__0 
       (.I0(\m100.u0/ethc0/r_reg[seq] [4]),
        .I1(\a9.x[0].r0_i_69__0_n_0 ),
        .I2(\m100.u0/rxwdata [22]),
        .I3(\m100.u0/ethc0/r_reg[ipcrc_n_0_][6] ),
        .I4(\a9.x[0].r0_i_70_n_0 ),
        .I5(\a9.x[0].r0_i_71__0_n_0 ),
        .O(\a9.x[0].r0_i_40__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF8C888C8)) 
    \a9.x[0].r0_i_41 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\m100.u0/rxwdata [4]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\a9.x[0].r0_i_68__0_n_0 ),
        .I5(\a9.x[0].r0_i_69_n_0 ),
        .O(\a9.x[0].r0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \a9.x[0].r0_i_41__0 
       (.I0(\a9.x[0].r0_i_57__0_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[udpsrc_n_0_][6] ),
        .I2(\a9.x[0].r0_i_72_n_0 ),
        .I3(\a9.x[0].r0_i_80__0_n_5 ),
        .I4(\a9.x[0].r0_i_81_n_0 ),
        .I5(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_41__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF8C888C8)) 
    \a9.x[0].r0_i_42 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\m100.u0/rxwdata [3]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\a9.x[0].r0_i_70__0_n_0 ),
        .I5(\a9.x[0].r0_i_71_n_0 ),
        .O(\a9.x[0].r0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFF0F0E2E20000)) 
    \a9.x[0].r0_i_42__0 
       (.I0(\m100.u0/ethc0/r_reg[seq] [3]),
        .I1(\a9.x[0].r0_i_69__0_n_0 ),
        .I2(\m100.u0/rxwdata [21]),
        .I3(\m100.u0/ethc0/r_reg[ipcrc_n_0_][5] ),
        .I4(\a9.x[0].r0_i_70_n_0 ),
        .I5(\a9.x[0].r0_i_71__0_n_0 ),
        .O(\a9.x[0].r0_i_42__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF8C888C8)) 
    \a9.x[0].r0_i_43 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\m100.u0/rxwdata [2]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\a9.x[0].r0_i_72__0_n_0 ),
        .I5(\a9.x[0].r0_i_73_n_0 ),
        .O(\a9.x[0].r0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \a9.x[0].r0_i_43__0 
       (.I0(\a9.x[0].r0_i_57__0_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[udpsrc_n_0_][5] ),
        .I2(\a9.x[0].r0_i_72_n_0 ),
        .I3(\a9.x[0].r0_i_80__0_n_6 ),
        .I4(\a9.x[0].r0_i_82_n_0 ),
        .I5(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_43__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF8C888C8)) 
    \a9.x[0].r0_i_44 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\m100.u0/rxwdata [1]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\a9.x[0].r0_i_74__0_n_0 ),
        .I5(\a9.x[0].r0_i_75_n_0 ),
        .O(\a9.x[0].r0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFF0F0E2E20000)) 
    \a9.x[0].r0_i_44__0 
       (.I0(\m100.u0/ethc0/r_reg[seq] [2]),
        .I1(\a9.x[0].r0_i_69__0_n_0 ),
        .I2(\m100.u0/rxwdata [20]),
        .I3(\m100.u0/ethc0/r_reg[ipcrc_n_0_][4] ),
        .I4(\a9.x[0].r0_i_70_n_0 ),
        .I5(\a9.x[0].r0_i_71__0_n_0 ),
        .O(\a9.x[0].r0_i_44__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF8C888C8)) 
    \a9.x[0].r0_i_45 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\m100.u0/rxwdata [0]),
        .I2(\a9.x[0].r0_i_22_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\a9.x[0].r0_i_76__0_n_0 ),
        .I5(\a9.x[0].r0_i_77_n_0 ),
        .O(\a9.x[0].r0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \a9.x[0].r0_i_45__0 
       (.I0(\a9.x[0].r0_i_57__0_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[udpsrc_n_0_][4] ),
        .I2(\a9.x[0].r0_i_72_n_0 ),
        .I3(\a9.x[0].r0_i_80__0_n_7 ),
        .I4(\a9.x[0].r0_i_83_n_0 ),
        .I5(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_45__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFF0F0E2E20000)) 
    \a9.x[0].r0_i_46 
       (.I0(\m100.u0/ethc0/r_reg[seq] [1]),
        .I1(\a9.x[0].r0_i_69__0_n_0 ),
        .I2(\m100.u0/rxwdata [19]),
        .I3(\m100.u0/ethc0/r_reg[ipcrc_n_0_][3] ),
        .I4(\a9.x[0].r0_i_70_n_0 ),
        .I5(\a9.x[0].r0_i_71__0_n_0 ),
        .O(\a9.x[0].r0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_46__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][47] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][15] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [15]),
        .O(\a9.x[0].r0_i_46__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAFEAAAA)) 
    \a9.x[0].r0_i_47 
       (.I0(\a9.x[0].r0_i_84_n_0 ),
        .I1(\a9.x[0].r0_i_55_n_0 ),
        .I2(\m100.u0/rxwdata [19]),
        .I3(\a9.x[0].r0_i_85_n_0 ),
        .I4(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_47__0 
       (.I0(\m100.u0/rxwdata [15]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][47] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][15] ),
        .O(\a9.x[0].r0_i_47__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFF0F0E2E20000)) 
    \a9.x[0].r0_i_48 
       (.I0(\m100.u0/ethc0/r_reg[seq] [0]),
        .I1(\a9.x[0].r0_i_69__0_n_0 ),
        .I2(\m100.u0/rxwdata [18]),
        .I3(\m100.u0/ethc0/r_reg[ipcrc_n_0_][2] ),
        .I4(\a9.x[0].r0_i_70_n_0 ),
        .I5(\a9.x[0].r0_i_71__0_n_0 ),
        .O(\a9.x[0].r0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_48__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][46] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][14] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [14]),
        .O(\a9.x[0].r0_i_48__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \a9.x[0].r0_i_49 
       (.I0(\a9.x[0].r0_i_57__0_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[udpsrc_n_0_][2] ),
        .I2(\a9.x[0].r0_i_72_n_0 ),
        .I3(\a9.x[0].r0_i_86__0_n_5 ),
        .I4(\a9.x[0].r0_i_87_n_0 ),
        .I5(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_49__0 
       (.I0(\m100.u0/rxwdata [14]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][46] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][14] ),
        .O(\a9.x[0].r0_i_49__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B8B8B8B8B8)) 
    \a9.x[0].r0_i_4__0 
       (.I0(\m100.u0/rxwdata [29]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_25__0_n_0 ),
        .I3(\a9.x[0].r0_i_26__0_n_0 ),
        .I4(\a9.x[0].r0_i_22_n_0 ),
        .I5(\r[rcntl][6]_i_5_n_0 ),
        .O(\m100.u0/datain [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_4__1 
       (.I0(\m100.u0/erdata [29]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [29]),
        .O(\m100.u0/txwdata [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FE0E)) 
    \a9.x[0].r0_i_5 
       (.I0(\a9.x[0].r0_i_28_n_0 ),
        .I1(\a9.x[0].r0_i_29_n_0 ),
        .I2(\m100.u0/ethc0/swap ),
        .I3(\m100.u0/rxwdata [12]),
        .I4(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0FFF77FF0F0022FF)) 
    \a9.x[0].r0_i_50 
       (.I0(\r[ewr]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/v[nak]1 ),
        .I2(\m100.u0/ethc0/r_reg[ipcrc_n_0_][1] ),
        .I3(\a9.x[0].r0_i_70_n_0 ),
        .I4(\a9.x[0].r0_i_71__0_n_0 ),
        .I5(\m100.u0/rxwdata [17]),
        .O(\a9.x[0].r0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_50__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][45] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][13] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [13]),
        .O(\a9.x[0].r0_i_50__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAFEAAAA)) 
    \a9.x[0].r0_i_51 
       (.I0(\a9.x[0].r0_i_88_n_0 ),
        .I1(\a9.x[0].r0_i_55_n_0 ),
        .I2(\m100.u0/rxwdata [17]),
        .I3(\a9.x[0].r0_i_89_n_0 ),
        .I4(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_51__0 
       (.I0(\m100.u0/rxwdata [13]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][45] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][13] ),
        .O(\a9.x[0].r0_i_51__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCC04FFFFCC04CC04)) 
    \a9.x[0].r0_i_52 
       (.I0(\a9.x[0].r0_i_90_n_0 ),
        .I1(\m100.u0/rxwdata [16]),
        .I2(\a9.x[0].r0_i_91_n_0 ),
        .I3(\a9.x[0].r0_i_72_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ipcrc_n_0_][0] ),
        .I5(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_52__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][44] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][12] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [12]),
        .O(\a9.x[0].r0_i_52__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAFEAAAA)) 
    \a9.x[0].r0_i_53 
       (.I0(\a9.x[0].r0_i_92_n_0 ),
        .I1(\a9.x[0].r0_i_55_n_0 ),
        .I2(\m100.u0/rxwdata [16]),
        .I3(\a9.x[0].r0_i_93_n_0 ),
        .I4(\a9.x[0].r0_i_22_n_0 ),
        .O(\a9.x[0].r0_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_53__0 
       (.I0(\m100.u0/rxwdata [12]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][44] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][12] ),
        .O(\a9.x[0].r0_i_53__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00007070000000FF)) 
    \a9.x[0].r0_i_54 
       (.I0(\FSM_sequential_r[edclrstate][3]_i_21_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/v[writeok]1 ),
        .I3(\r[erxidle]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\a9.x[0].r0_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_54__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][43] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][11] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [11]),
        .O(\a9.x[0].r0_i_54__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000001400003C00)) 
    \a9.x[0].r0_i_55 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I2(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\a9.x[0].r0_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_55__0 
       (.I0(\m100.u0/rxwdata [11]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][43] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][11] ),
        .O(\a9.x[0].r0_i_55__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \a9.x[0].r0_i_56 
       (.I0(\a9.x[0].r0_i_78__0_n_0 ),
        .I1(\a9.x[0].r0_i_79__0_n_0 ),
        .O(\a9.x[0].r0_i_56_n_0 ),
        .S(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFDFFFDFFFCF3FFFF)) 
    \a9.x[0].r0_i_56__0 
       (.I0(\m100.u0/rxwdata [15]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][31] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\a9.x[0].r0_i_56__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0C00AC000A000C0)) 
    \a9.x[0].r0_i_57 
       (.I0(\m100.u0/ethc0/r_reg[nak_n_0_] ),
        .I1(\a9.x[0].r0_i_80_n_1 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA202)) 
    \a9.x[0].r0_i_57__0 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_57__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0B3B0A0)) 
    \a9.x[0].r0_i_58 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\a9.x[0].r0_i_91_n_0 ),
        .I2(\m100.u0/rxwdata [31]),
        .I3(\a9.x[0].r0_i_69__0_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[seq] [13]),
        .O(\a9.x[0].r0_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \a9.x[0].r0_i_58__0 
       (.I0(\a9.x[0].r0_i_81__0_n_0 ),
        .I1(\a9.x[0].r0_i_82__0_n_0 ),
        .O(\a9.x[0].r0_i_58__0_n_0 ),
        .S(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0C00AC000A000C0)) 
    \a9.x[0].r0_i_59 
       (.I0(\m100.u0/ethc0/r_reg[oplen_n_0_][9] ),
        .I1(\a9.x[0].r0_i_80_n_6 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000140014141400)) 
    \a9.x[0].r0_i_59__0 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I2(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .O(\m100.u0/ethc0/swap12_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B8B8B8B8B8)) 
    \a9.x[0].r0_i_5__0 
       (.I0(\m100.u0/rxwdata [28]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_27__0_n_0 ),
        .I3(\a9.x[0].r0_i_28__0_n_0 ),
        .I4(\a9.x[0].r0_i_22_n_0 ),
        .I5(\r[rcntl][6]_i_5_n_0 ),
        .O(\m100.u0/datain [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_5__1 
       (.I0(\m100.u0/erdata [28]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [28]),
        .O(\m100.u0/txwdata [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FE0E)) 
    \a9.x[0].r0_i_6 
       (.I0(\a9.x[0].r0_i_30_n_0 ),
        .I1(\a9.x[0].r0_i_31__0_n_0 ),
        .I2(\m100.u0/ethc0/swap ),
        .I3(\m100.u0/rxwdata [11]),
        .I4(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000060000000000)) 
    \a9.x[0].r0_i_60 
       (.I0(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I1(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\m100.u0/ethc0/setmz11_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \a9.x[0].r0_i_60__0 
       (.I0(\a9.x[0].r0_i_83__0_n_0 ),
        .I1(\a9.x[0].r0_i_84__0_n_0 ),
        .O(\a9.x[0].r0_i_60__0_n_0 ),
        .S(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0C00AC000A000C0)) 
    \a9.x[0].r0_i_61 
       (.I0(\m100.u0/ethc0/r_reg[oplen_n_0_][8] ),
        .I1(\a9.x[0].r0_i_80_n_7 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \a9.x[0].r0_i_61__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][30] ),
        .I1(\m100.u0/ethc0/v[writeok]1 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\a9.x[0].r0_i_94__0_n_0 ),
        .I4(\m100.u0/rxwdata [14]),
        .I5(\m100.u0/ethc0/setmz11_out ),
        .O(\a9.x[0].r0_i_61__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0B3B0A0)) 
    \a9.x[0].r0_i_62 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\a9.x[0].r0_i_91_n_0 ),
        .I2(\m100.u0/rxwdata [30]),
        .I3(\a9.x[0].r0_i_69__0_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[seq] [12]),
        .O(\a9.x[0].r0_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \a9.x[0].r0_i_62__0 
       (.I0(\a9.x[0].r0_i_85__0_n_0 ),
        .I1(\a9.x[0].r0_i_86_n_0 ),
        .O(\a9.x[0].r0_i_62__0_n_0 ),
        .S(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0C00AC000A000C0)) 
    \a9.x[0].r0_i_63 
       (.I0(\m100.u0/ethc0/r_reg[oplen_n_0_][7] ),
        .I1(\a9.x[0].r0_i_87__0_n_4 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \a9.x[0].r0_i_63__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][29] ),
        .I1(\m100.u0/ethc0/v[writeok]1 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\a9.x[0].r0_i_94__0_n_0 ),
        .I4(\m100.u0/rxwdata [13]),
        .I5(\m100.u0/ethc0/setmz11_out ),
        .O(\a9.x[0].r0_i_63__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0B3B0A0)) 
    \a9.x[0].r0_i_64 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\a9.x[0].r0_i_91_n_0 ),
        .I2(\m100.u0/rxwdata [29]),
        .I3(\a9.x[0].r0_i_69__0_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[seq] [11]),
        .O(\a9.x[0].r0_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \a9.x[0].r0_i_64__0 
       (.I0(\a9.x[0].r0_i_88__0_n_0 ),
        .I1(\a9.x[0].r0_i_89__0_n_0 ),
        .O(\a9.x[0].r0_i_64__0_n_0 ),
        .S(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0C00AC000A000C0)) 
    \a9.x[0].r0_i_65 
       (.I0(\m100.u0/ethc0/r_reg[oplen_n_0_][6] ),
        .I1(\a9.x[0].r0_i_87__0_n_5 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \a9.x[0].r0_i_65__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][28] ),
        .I1(\m100.u0/ethc0/v[writeok]1 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\a9.x[0].r0_i_94__0_n_0 ),
        .I4(\m100.u0/rxwdata [12]),
        .I5(\m100.u0/ethc0/setmz11_out ),
        .O(\a9.x[0].r0_i_65__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0B3B0A0)) 
    \a9.x[0].r0_i_66 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\a9.x[0].r0_i_91_n_0 ),
        .I2(\m100.u0/rxwdata [28]),
        .I3(\a9.x[0].r0_i_69__0_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[seq] [10]),
        .O(\a9.x[0].r0_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \a9.x[0].r0_i_66__0 
       (.I0(\a9.x[0].r0_i_90__0_n_0 ),
        .I1(\a9.x[0].r0_i_91__0_n_0 ),
        .O(\a9.x[0].r0_i_66__0_n_0 ),
        .S(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0C00AC000A000C0)) 
    \a9.x[0].r0_i_67 
       (.I0(\m100.u0/ethc0/r_reg[oplen_n_0_][5] ),
        .I1(\a9.x[0].r0_i_87__0_n_6 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \a9.x[0].r0_i_67__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][27] ),
        .I1(\m100.u0/ethc0/v[writeok]1 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\a9.x[0].r0_i_94__0_n_0 ),
        .I4(\m100.u0/rxwdata [11]),
        .I5(\m100.u0/ethc0/setmz11_out ),
        .O(\a9.x[0].r0_i_67__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0B3B0A0)) 
    \a9.x[0].r0_i_68 
       (.I0(\a9.x[0].r0_i_72_n_0 ),
        .I1(\a9.x[0].r0_i_91_n_0 ),
        .I2(\m100.u0/rxwdata [27]),
        .I3(\a9.x[0].r0_i_69__0_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[seq] [9]),
        .O(\a9.x[0].r0_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \a9.x[0].r0_i_68__0 
       (.I0(\a9.x[0].r0_i_92__0_n_0 ),
        .I1(\a9.x[0].r0_i_93__0_n_0 ),
        .O(\a9.x[0].r0_i_68__0_n_0 ),
        .S(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0C00AC000A000C0)) 
    \a9.x[0].r0_i_69 
       (.I0(\m100.u0/ethc0/r_reg[oplen_n_0_][4] ),
        .I1(\a9.x[0].r0_i_87__0_n_7 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    \a9.x[0].r0_i_69__0 
       (.I0(\m100.u0/ethc0/v[nak]1 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/v[writeok]1 ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\a9.x[0].r0_i_69__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B8B8B8B8B8)) 
    \a9.x[0].r0_i_6__0 
       (.I0(\m100.u0/rxwdata [27]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_29__0_n_0 ),
        .I3(\a9.x[0].r0_i_30__0_n_0 ),
        .I4(\a9.x[0].r0_i_22_n_0 ),
        .I5(\r[rcntl][6]_i_5_n_0 ),
        .O(\m100.u0/datain [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_6__1 
       (.I0(\m100.u0/erdata [27]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [27]),
        .O(\m100.u0/txwdata [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \a9.x[0].r0_i_7 
       (.I0(\a9.x[0].r0_i_32_n_0 ),
        .I1(\r[rcntl][6]_i_5_n_0 ),
        .I2(\a9.x[0].r0_i_33__0_n_0 ),
        .I3(\m100.u0/ethc0/swap ),
        .I4(\m100.u0/rxwdata [10]),
        .I5(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22C0)) 
    \a9.x[0].r0_i_70 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\a9.x[0].r0_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \a9.x[0].r0_i_70__0 
       (.I0(\a9.x[0].r0_i_94_n_0 ),
        .I1(\a9.x[0].r0_i_95_n_0 ),
        .O(\a9.x[0].r0_i_70__0_n_0 ),
        .S(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0C00AC000A000C0)) 
    \a9.x[0].r0_i_71 
       (.I0(\m100.u0/ethc0/r_reg[oplen_n_0_][3] ),
        .I1(\a9.x[0].r0_i_111_n_4 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h70DF)) 
    \a9.x[0].r0_i_71__0 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\a9.x[0].r0_i_71__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h159D)) 
    \a9.x[0].r0_i_72 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\a9.x[0].r0_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \a9.x[0].r0_i_72__0 
       (.I0(\a9.x[0].r0_i_96_n_0 ),
        .I1(\a9.x[0].r0_i_97_n_0 ),
        .O(\a9.x[0].r0_i_72__0_n_0 ),
        .S(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0C00AC000A000C0)) 
    \a9.x[0].r0_i_73 
       (.I0(\m100.u0/ethc0/r_reg[oplen_n_0_][2] ),
        .I1(\a9.x[0].r0_i_111_n_5 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \a9.x[0].r0_i_73__0 
       (.CI(\a9.x[0].r0_i_80__0_n_0 ),
        .CO({\a9.x[0].r0_i_73__0_n_0 ,\a9.x[0].r0_i_73__0_n_1 ,\a9.x[0].r0_i_73__0_n_2 ,\a9.x[0].r0_i_73__0_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\a9.x[0].r0_i_73__0_n_4 ,\a9.x[0].r0_i_73__0_n_5 ,\a9.x[0].r0_i_73__0_n_6 ,\a9.x[0].r0_i_73__0_n_7 }),
        .S({etho,apbo,\m100.u0/ethc0/r_reg[applength]__0 [9:8]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8FFFF8B880000)) 
    \a9.x[0].r0_i_74 
       (.I0(\a9.x[0].r0_i_97__0_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\a9.x[0].r0_i_94__0_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][26] ),
        .I4(\m100.u0/ethc0/v[writeok]1 ),
        .I5(\m100.u0/rxwdata [26]),
        .O(\a9.x[0].r0_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \a9.x[0].r0_i_74__0 
       (.I0(\a9.x[0].r0_i_98__0_n_0 ),
        .I1(\a9.x[0].r0_i_99_n_0 ),
        .O(\a9.x[0].r0_i_74__0_n_0 ),
        .S(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0C00AC000A000C0)) 
    \a9.x[0].r0_i_75 
       (.I0(\m100.u0/ethc0/r_reg[oplen_n_0_][1] ),
        .I1(\a9.x[0].r0_i_111_n_6 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0CAA0CA0A0AAACA)) 
    \a9.x[0].r0_i_75__0 
       (.I0(\a9.x[0].r0_i_73__0_n_6 ),
        .I1(\m100.u0/ethc0/r_reg[udpsrc_n_0_][9] ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_75__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \a9.x[0].r0_i_76 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][25] ),
        .I1(\m100.u0/ethc0/v[writeok]1 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\a9.x[0].r0_i_94__0_n_0 ),
        .I4(\m100.u0/rxwdata [9]),
        .I5(\m100.u0/ethc0/setmz11_out ),
        .O(\a9.x[0].r0_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \a9.x[0].r0_i_76__0 
       (.I0(\a9.x ),
        .I1(\a9.x[0].r0_i_101_n_0 ),
        .O(\a9.x[0].r0_i_76__0_n_0 ),
        .S(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0C00AC000A000C0)) 
    \a9.x[0].r0_i_77 
       (.I0(\m100.u0/ethc0/r_reg[oplen_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[applength]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8FFFF8B880000)) 
    \a9.x[0].r0_i_77__0 
       (.I0(\a9.x[0].r0_i_98_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\a9.x[0].r0_i_94__0_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][24] ),
        .I4(\m100.u0/ethc0/v[writeok]1 ),
        .I5(\m100.u0/rxwdata [24]),
        .O(\a9.x[0].r0_i_77__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0CAA0CA0A0AAACA)) 
    \a9.x[0].r0_i_78 
       (.I0(\a9.x[0].r0_i_80__0_n_4 ),
        .I1(\m100.u0/ethc0/r_reg[udpsrc_n_0_][7] ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_78__0 
       (.I0(\m100.u0/rxwdata [10]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][42] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][10] ),
        .O(\a9.x[0].r0_i_78__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \a9.x[0].r0_i_79 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][23] ),
        .I1(\m100.u0/ethc0/v[writeok]1 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\a9.x[0].r0_i_94__0_n_0 ),
        .I4(\m100.u0/rxwdata [7]),
        .I5(\m100.u0/ethc0/setmz11_out ),
        .O(\a9.x[0].r0_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_79__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][42] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][10] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [10]),
        .O(\a9.x[0].r0_i_79__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB8BB8888B888)) 
    \a9.x[0].r0_i_7__0 
       (.I0(\m100.u0/rxwdata [26]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_31_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\a9.x[0].r0_i_32__0_n_0 ),
        .O(\m100.u0/datain [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_7__1 
       (.I0(\m100.u0/erdata [26]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [26]),
        .O(\m100.u0/txwdata [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \a9.x[0].r0_i_8 
       (.I0(\a9.x[0].r0_i_34_n_0 ),
        .I1(\r[rcntl][6]_i_5_n_0 ),
        .I2(\a9.x[0].r0_i_35__0_n_0 ),
        .I3(\m100.u0/ethc0/swap ),
        .I4(\m100.u0/rxwdata [9]),
        .I5(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \a9.x[0].r0_i_80 
       (.CI(\a9.x[0].r0_i_87__0_n_0 ),
        .CO({\a9.x[0].r0_i_80_n_0 ,\a9.x[0].r0_i_80_n_1 ,\a9.x[0].r0_i_80_n_2 ,\a9.x[0].r0_i_80_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\a9.x[0].r0_i_80_n_4 ,\a9.x[0].r0_i_80_n_5 ,\a9.x[0].r0_i_80_n_6 ,\a9.x[0].r0_i_80_n_7 }),
        .S({etho,apbo,\m100.u0/ethc0/r_reg[applength]__0 [9:8]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \a9.x[0].r0_i_80__0 
       (.CI(\a9.x[0].r0_i_86__0_n_0 ),
        .CO({\a9.x[0].r0_i_80__0_n_0 ,\a9.x[0].r0_i_80__0_n_1 ,\a9.x[0].r0_i_80__0_n_2 ,\a9.x[0].r0_i_80__0_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,\m100.u0/ethc0/r_reg[applength]__0 [5],etho}),
        .O({\a9.x[0].r0_i_80__0_n_4 ,\a9.x[0].r0_i_80__0_n_5 ,\a9.x[0].r0_i_80__0_n_6 ,\a9.x[0].r0_i_80__0_n_7 }),
        .S({\m100.u0/ethc0/r_reg[applength]__0 [7:6],\a9.x[0].r0_i_101__0_n_0 ,\m100.u0/ethc0/r_reg[applength]__0 [4]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8FFFF8B880000)) 
    \a9.x[0].r0_i_81 
       (.I0(\a9.x[0].r0_i_103_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\a9.x[0].r0_i_94__0_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][22] ),
        .I4(\m100.u0/ethc0/v[writeok]1 ),
        .I5(\m100.u0/rxwdata [22]),
        .O(\a9.x[0].r0_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_81__0 
       (.I0(\m100.u0/rxwdata [9]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][41] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][9] ),
        .O(\a9.x[0].r0_i_81__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8FFFF8B880000)) 
    \a9.x[0].r0_i_82 
       (.I0(\a9.x[0].r0_i_104_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\a9.x[0].r0_i_94__0_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][21] ),
        .I4(\m100.u0/ethc0/v[writeok]1 ),
        .I5(\m100.u0/rxwdata [21]),
        .O(\a9.x[0].r0_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_82__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][41] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][9] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [9]),
        .O(\a9.x[0].r0_i_82__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8FFFF8B880000)) 
    \a9.x[0].r0_i_83 
       (.I0(\a9.x[0].r0_i_105_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\a9.x[0].r0_i_94__0_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][20] ),
        .I4(\m100.u0/ethc0/v[writeok]1 ),
        .I5(\m100.u0/rxwdata [20]),
        .O(\a9.x[0].r0_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_83__0 
       (.I0(\m100.u0/rxwdata [8]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][40] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][8] ),
        .O(\a9.x[0].r0_i_83__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0CAA0CA0A0AAACA)) 
    \a9.x[0].r0_i_84 
       (.I0(\a9.x[0].r0_i_86__0_n_4 ),
        .I1(\m100.u0/ethc0/r_reg[udpsrc_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_84__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][40] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][8] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [8]),
        .O(\a9.x[0].r0_i_84__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \a9.x[0].r0_i_85 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][19] ),
        .I1(\m100.u0/ethc0/v[writeok]1 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\a9.x[0].r0_i_94__0_n_0 ),
        .I4(\m100.u0/rxwdata [3]),
        .I5(\m100.u0/ethc0/setmz11_out ),
        .O(\a9.x[0].r0_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_85__0 
       (.I0(\m100.u0/rxwdata [7]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][39] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][7] ),
        .O(\a9.x[0].r0_i_85__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_86 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][39] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][7] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [7]),
        .O(\a9.x[0].r0_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \a9.x[0].r0_i_86__0 
       (.CI(etho),
        .CO({\a9.x[0].r0_i_86__0_n_0 ,\a9.x[0].r0_i_86__0_n_1 ,\a9.x[0].r0_i_86__0_n_2 ,\a9.x[0].r0_i_86__0_n_3 }),
        .CYINIT(etho),
        .DI({etho,\m100.u0/ethc0/r_reg[applength]__0 [2:1],etho}),
        .O({\a9.x[0].r0_i_86__0_n_4 ,\a9.x[0].r0_i_86__0_n_5 ,\a9.x[0].r0_i_86__0_n_6 ,\a9.x[0].r0_i_86__0_n_7 }),
        .S({\m100.u0/ethc0/r_reg[applength]__0 [3],\a9.x[0].r0_i_107__0_n_0 ,\a9.x[0].r0_i_108_n_0 ,\m100.u0/ethc0/r_reg[applength]__0 [0]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8FFFF8B880000)) 
    \a9.x[0].r0_i_87 
       (.I0(\a9.x[0].r0_i_110_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\a9.x[0].r0_i_94__0_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][18] ),
        .I4(\m100.u0/ethc0/v[writeok]1 ),
        .I5(\m100.u0/rxwdata [18]),
        .O(\a9.x[0].r0_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \a9.x[0].r0_i_87__0 
       (.CI(\a9.x[0].r0_i_111_n_0 ),
        .CO({\a9.x[0].r0_i_87__0_n_0 ,\a9.x[0].r0_i_87__0_n_1 ,\a9.x[0].r0_i_87__0_n_2 ,\a9.x[0].r0_i_87__0_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,\m100.u0/ethc0/r_reg[applength]__0 [4]}),
        .O({\a9.x[0].r0_i_87__0_n_4 ,\a9.x[0].r0_i_87__0_n_5 ,\a9.x[0].r0_i_87__0_n_6 ,\a9.x[0].r0_i_87__0_n_7 }),
        .S({\m100.u0/ethc0/r_reg[applength]__0 [7:5],\a9.x[0].r0_i_107_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0CAA0CA0A0AAACA)) 
    \a9.x[0].r0_i_88 
       (.I0(\a9.x[0].r0_i_86__0_n_6 ),
        .I1(\m100.u0/ethc0/r_reg[udpsrc_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_88__0 
       (.I0(\m100.u0/rxwdata [6]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][38] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][6] ),
        .O(\a9.x[0].r0_i_88__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \a9.x[0].r0_i_89 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][17] ),
        .I1(\m100.u0/ethc0/v[writeok]1 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\a9.x[0].r0_i_94__0_n_0 ),
        .I4(\m100.u0/rxwdata [1]),
        .I5(\m100.u0/ethc0/setmz11_out ),
        .O(\a9.x[0].r0_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_89__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][38] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][6] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [6]),
        .O(\a9.x[0].r0_i_89__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB8BB8888B888)) 
    \a9.x[0].r0_i_8__0 
       (.I0(\m100.u0/rxwdata [25]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_33_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\a9.x[0].r0_i_34__0_n_0 ),
        .O(\m100.u0/datain [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_8__1 
       (.I0(\m100.u0/erdata [25]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [25]),
        .O(\m100.u0/txwdata [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \a9.x[0].r0_i_9 
       (.I0(\a9.x[0].r0_i_36_n_0 ),
        .I1(\r[rcntl][6]_i_5_n_0 ),
        .I2(\a9.x[0].r0_i_37__0_n_0 ),
        .I3(\m100.u0/ethc0/swap ),
        .I4(\m100.u0/rxwdata [8]),
        .I5(\m100.u0/ethc0/setmz ),
        .O(\m100.u0/datain [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \a9.x[0].r0_i_90 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/v[writeok]1 ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\r[ipcrc][11]_i_13_n_0 ),
        .O(\a9.x[0].r0_i_90_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_90__0 
       (.I0(\m100.u0/rxwdata [5]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][37] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][5] ),
        .O(\a9.x[0].r0_i_90__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFDBF)) 
    \a9.x[0].r0_i_91 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\a9.x[0].r0_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_91__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][37] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][5] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [5]),
        .O(\a9.x[0].r0_i_91__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0CAA0CA0A0AAACA)) 
    \a9.x[0].r0_i_92 
       (.I0(\a9.x[0].r0_i_111_n_7 ),
        .I1(\m100.u0/ethc0/r_reg[udpsrc_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\a9.x[0].r0_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_92__0 
       (.I0(\m100.u0/rxwdata [4]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][36] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][4] ),
        .O(\a9.x[0].r0_i_92__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \a9.x[0].r0_i_93 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][16] ),
        .I1(\m100.u0/ethc0/v[writeok]1 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\a9.x[0].r0_i_94__0_n_0 ),
        .I4(\m100.u0/rxwdata [0]),
        .I5(\m100.u0/ethc0/setmz11_out ),
        .O(\a9.x[0].r0_i_93_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_93__0 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][36] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [4]),
        .O(\a9.x[0].r0_i_93__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_94 
       (.I0(\m100.u0/rxwdata [3]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][35] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][3] ),
        .O(\a9.x[0].r0_i_94_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hED)) 
    \a9.x[0].r0_i_94__0 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .O(\a9.x[0].r0_i_94__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_95 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][35] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [3]),
        .O(\a9.x[0].r0_i_95_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_96 
       (.I0(\m100.u0/rxwdata [2]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][34] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][2] ),
        .O(\a9.x[0].r0_i_96_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_97 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][34] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [2]),
        .O(\a9.x[0].r0_i_97_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \a9.x[0].r0_i_97__0 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/rxwdata [10]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I4(\m100.u0/rxwdata [26]),
        .O(\a9.x[0].r0_i_97__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \a9.x[0].r0_i_98 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/rxwdata [8]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I4(\m100.u0/rxwdata [24]),
        .O(\a9.x[0].r0_i_98_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABAEA8AEABA2A8A2)) 
    \a9.x[0].r0_i_98__0 
       (.I0(\m100.u0/rxwdata [1]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][33] ),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][1] ),
        .O(\a9.x[0].r0_i_98__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB8FF0000B800)) 
    \a9.x[0].r0_i_99 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][33] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/rxwdata [1]),
        .O(\a9.x[0].r0_i_99_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB8BB8888B888)) 
    \a9.x[0].r0_i_9__0 
       (.I0(\m100.u0/rxwdata [24]),
        .I1(\m100.u0/ethc0/swap ),
        .I2(\a9.x[0].r0_i_35_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\a9.x[0].r0_i_36__0_n_0 ),
        .O(\m100.u0/datain [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    \a9.x[0].r0_i_9__1 
       (.I0(\m100.u0/erdata [24]),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\ahbmi[hrdata] [24]),
        .O(\m100.u0/txwdata [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][10]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [10]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [10]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][11]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [11]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [11]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][12]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [12]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [12]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][13]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [13]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [13]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][14]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [14]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [14]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][15]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [15]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [15]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][16]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [16]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [16]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][17]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [17]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [17]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][18]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [18]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [18]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][19]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [19]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [19]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][1]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [1]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [1]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][20]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [20]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [20]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][21]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [21]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [21]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][22]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [22]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [22]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][23]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [23]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [23]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][24]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [24]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [24]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][25]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [25]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [25]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][26]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [26]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [26]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][27]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [27]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [27]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][28]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [28]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [28]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][29]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [29]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [29]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][2]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [2]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [2]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][30]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [30]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [30]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][31]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [31]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [31]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][3]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [3]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [3]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][4]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [4]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [4]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][5]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [5]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [5]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][6]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [6]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [6]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][7]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [7]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [7]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][8]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [8]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [8]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[haddr][9]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [9]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [9]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\^ahbmo[haddr] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \ahbmo[hbusreq]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .O(ahbmo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0404040000040000)) 
    \ahbmo[htrans][0]_INST_0 
       (.I0(\ahbmo[htrans][0]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/ahb0/r_reg ),
        .I2(\m100.u0/ethc0/ahb0/r_reg[bb]__0 ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .O(\ahbmo[htrans] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \ahbmo[htrans][0]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/ahb0/r_reg[error]__0 ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .O(\ahbmo[htrans][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h000E)) 
    \ahbmo[htrans][1]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I2(\m100.u0/ethc0/ahb0/r_reg[error]__0 ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .O(\ahbmo[htrans] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][0]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][0] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][0] ),
        .O(\ahbmo[hwdata] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][10]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][10] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][10] ),
        .O(\ahbmo[hwdata] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][11]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][11] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][11] ),
        .O(\ahbmo[hwdata] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][12]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][12] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][12] ),
        .O(\ahbmo[hwdata] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][13]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][13] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][13] ),
        .O(\ahbmo[hwdata] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][14]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][14] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][14] ),
        .O(\ahbmo[hwdata] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][15]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][15] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][15] ),
        .O(\ahbmo[hwdata] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][16]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][16] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][16] ),
        .O(\ahbmo[hwdata] [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][17]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][17] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][17] ),
        .O(\ahbmo[hwdata] [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][18]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][18] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][18] ),
        .O(\ahbmo[hwdata] [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][19]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][19] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][19] ),
        .O(\ahbmo[hwdata] [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][1]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][1] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][1] ),
        .O(\ahbmo[hwdata] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][20]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][20] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][20] ),
        .O(\ahbmo[hwdata] [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][21]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][21] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][21] ),
        .O(\ahbmo[hwdata] [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][22]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][22] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][22] ),
        .O(\ahbmo[hwdata] [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][23]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][23] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][23] ),
        .O(\ahbmo[hwdata] [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][24]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][24] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][24] ),
        .O(\ahbmo[hwdata] [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][25]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][25] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][25] ),
        .O(\ahbmo[hwdata] [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][26]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][26] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][26] ),
        .O(\ahbmo[hwdata] [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][27]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][27] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][27] ),
        .O(\ahbmo[hwdata] [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][28]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][28] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][28] ),
        .O(\ahbmo[hwdata] [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][29]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][29] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][29] ),
        .O(\ahbmo[hwdata] [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][2]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][2] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][2] ),
        .O(\ahbmo[hwdata] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][30]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][30] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][30] ),
        .O(\ahbmo[hwdata] [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][31]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][31] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][31] ),
        .O(\ahbmo[hwdata] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][3]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][3] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][3] ),
        .O(\ahbmo[hwdata] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][4]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][4] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][4] ),
        .O(\ahbmo[hwdata] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][5]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][5] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][5] ),
        .O(\ahbmo[hwdata] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][6]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][6] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][6] ),
        .O(\ahbmo[hwdata] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][7]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][7] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][7] ),
        .O(\ahbmo[hwdata] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][8]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][8] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][8] ),
        .O(\ahbmo[hwdata] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \ahbmo[hwdata][9]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][9] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][9] ),
        .O(\ahbmo[hwdata] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAACAAACCCCCCCAC)) 
    \ahbmo[hwrite]_INST_0 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][write_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[rmsto][write_n_0_] ),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\ahbmo[hwrite] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF10000000)) 
    \apbo[pirq][12]_INST_0 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\apbo[pirq][12]_INST_0_i_1_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxirq]__0 ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\apbo[pirq][12]_INST_0_i_2_n_0 ),
        .O(\^apbo[pirq] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    \apbo[pirq][12]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_6_in [3]),
        .I1(\m100.u0/ethc0/ahb0/r_reg ),
        .I2(\ahbmi[hready] ),
        .I3(\ahbmi[hresp] [1]),
        .I4(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I5(\ahbmi[hresp] [0]),
        .O(\apbo[pirq][12]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000002)) 
    \apbo[pirq][12]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txirqgen_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\apbo[pirq][12]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][0]_INST_0 
       (.I0(\apbo[prdata][0]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][0]_INST_0_i_2_n_0 ),
        .O(\apbo[prdata] [0]),
        .S(\apbi[paddr] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8380FFFF83800000)) 
    \apbo[prdata][0]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][0] ),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][write]__0 ),
        .I4(\apbi[paddr] [4]),
        .I5(\apbo[prdata][0]_INST_0_i_3_n_0 ),
        .O(\apbo[prdata][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00B00080)) 
    \apbo[prdata][0]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][0] ),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [4]),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][32] ),
        .O(\apbo[prdata][0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][0]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][32] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[status][rx_err_n_0_] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/p_6_in [0]),
        .O(\apbo[prdata][0]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF5410)) 
    \apbo[prdata][10]_INST_0 
       (.I0(\apbo[prdata][10]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][10]_INST_0_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[emacaddr_n_0_][10] ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][42] ),
        .I4(\apbo[prdata][10]_INST_0_i_3_n_0 ),
        .O(\apbo[prdata] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \apbo[prdata][10]_INST_0_i_1 
       (.I0(\apbi[paddr] [5]),
        .I1(\apbi[paddr] [4]),
        .I2(\apbi[paddr] [3]),
        .O(\apbo[prdata][10]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h15)) 
    \apbo[prdata][10]_INST_0_i_2 
       (.I0(\apbi[paddr] [4]),
        .I1(\apbi[paddr] [3]),
        .I2(\apbi[paddr] [2]),
        .O(\apbo[prdata][10]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4FFF44444444444)) 
    \apbo[prdata][10]_INST_0_i_3 
       (.I0(\apbo[prdata][14]_INST_0_i_5_n_0 ),
        .I1(\apbo[prdata][10]_INST_0_i_4_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mac_addr_n_0_][10] ),
        .I3(\apbi[paddr] [2]),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][42] ),
        .I5(\apbo[prdata][10]_INST_0_i_5_n_0 ),
        .O(\apbo[prdata][10]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][10]_INST_0_i_4 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][10] ),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][10] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [0]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [4]),
        .O(\apbo[prdata][10]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \apbo[prdata][10]_INST_0_i_5 
       (.I0(\apbi[paddr] [4]),
        .I1(\apbi[paddr] [5]),
        .I2(\apbi[paddr] [3]),
        .O(\apbo[prdata][10]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][11]_INST_0 
       (.I0(\apbo[prdata][11]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][11]_INST_0_i_2_n_0 ),
        .O(\apbo[prdata] [11]),
        .S(\apbi[paddr] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB888B888888888)) 
    \apbo[prdata][11]_INST_0_i_1 
       (.I0(\apbo[prdata][11]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [4]),
        .I2(\m100.u0/ethc0/r_reg[mac_addr_n_0_][43] ),
        .I3(\apbi[paddr] [2]),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][11] ),
        .I5(\apbi[paddr] [3]),
        .O(\apbo[prdata][11]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00B00080)) 
    \apbo[prdata][11]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][11] ),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [4]),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][43] ),
        .O(\apbo[prdata][11]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][11]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][11] ),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][11] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [1]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][phyadr_n_0_][0] ),
        .O(\apbo[prdata][11]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFEAFFEAFFFFFFEA)) 
    \apbo[prdata][12]_INST_0 
       (.I0(\apbo[prdata][12]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][14]_INST_0_i_2_n_0 ),
        .I2(\m100.u0/ethc0/p_6_in [12]),
        .I3(\apbo[prdata][12]_INST_0_i_2_n_0 ),
        .I4(\apbo[prdata][12]_INST_0_i_3_n_0 ),
        .I5(\apbo[prdata][14]_INST_0_i_5_n_0 ),
        .O(\apbo[prdata] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000CA0000000000)) 
    \apbo[prdata][12]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][44] ),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][12] ),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][12]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0202020000000200)) 
    \apbo[prdata][12]_INST_0_i_2 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[paddr] [5]),
        .I2(\apbi[paddr] [4]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][44] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mac_addr_n_0_][12] ),
        .O(\apbo[prdata][12]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][12]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][12] ),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][12] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [2]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][phyadr_n_0_][1] ),
        .O(\apbo[prdata][12]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][13]_INST_0 
       (.I0(\apbo[prdata][13]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][13]_INST_0_i_2_n_0 ),
        .O(\apbo[prdata] [13]),
        .S(\apbi[paddr] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB888B888888888)) 
    \apbo[prdata][13]_INST_0_i_1 
       (.I0(\apbo[prdata][13]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [4]),
        .I2(\m100.u0/ethc0/r_reg[mac_addr_n_0_][45] ),
        .I3(\apbi[paddr] [2]),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][13] ),
        .I5(\apbi[paddr] [3]),
        .O(\apbo[prdata][13]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00B00080)) 
    \apbo[prdata][13]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][13] ),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [4]),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][45] ),
        .O(\apbo[prdata][13]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][13]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][13] ),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][13] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [3]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/data2 ),
        .O(\apbo[prdata][13]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFEAFFEAFFFFFFEA)) 
    \apbo[prdata][14]_INST_0 
       (.I0(\apbo[prdata][14]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][14]_INST_0_i_2_n_0 ),
        .I2(\m100.u0/ethc0/p_6_in [14]),
        .I3(\apbo[prdata][14]_INST_0_i_3_n_0 ),
        .I4(\apbo[prdata][14]_INST_0_i_4_n_0 ),
        .I5(\apbo[prdata][14]_INST_0_i_5_n_0 ),
        .O(\apbo[prdata] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B0008000000000)) 
    \apbo[prdata][14]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][14] ),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [4]),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][46] ),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][14]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \apbo[prdata][14]_INST_0_i_2 
       (.I0(\apbi[paddr] [4]),
        .I1(\apbi[paddr] [5]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [2]),
        .O(\apbo[prdata][14]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0202020000000200)) 
    \apbo[prdata][14]_INST_0_i_3 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[paddr] [5]),
        .I2(\apbi[paddr] [4]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][46] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mac_addr_n_0_][14] ),
        .O(\apbo[prdata][14]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][14]_INST_0_i_4 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][14] ),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][14] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [4]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/data1 ),
        .O(\apbo[prdata][14]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \apbo[prdata][14]_INST_0_i_5 
       (.I0(\apbi[paddr] [5]),
        .I1(\apbi[paddr] [4]),
        .O(\apbo[prdata][14]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][15]_INST_0 
       (.I0(\apbo[prdata][15]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_2_n_0 ),
        .O(\apbo[prdata] [15]),
        .S(\apbi[paddr] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB888B888888888)) 
    \apbo[prdata][15]_INST_0_i_1 
       (.I0(\apbo[prdata][15]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [4]),
        .I2(\m100.u0/ethc0/r_reg[mac_addr_n_0_][47] ),
        .I3(\apbi[paddr] [2]),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][15] ),
        .I5(\apbi[paddr] [3]),
        .O(\apbo[prdata][15]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00B00080)) 
    \apbo[prdata][15]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][15] ),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [4]),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][47] ),
        .O(\apbo[prdata][15]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][15]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][15] ),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][15] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [5]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][phyadr_n_0_][4] ),
        .O(\apbo[prdata][15]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][16]_INST_0 
       (.I0(\apbo[prdata][16]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][16] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][16] ),
        .O(\apbo[prdata] [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][16]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [0]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][16] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [6]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .O(\apbo[prdata][16]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][17]_INST_0 
       (.I0(\apbo[prdata][17]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][17] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][17] ),
        .O(\apbo[prdata] [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][17]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [1]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][17] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [7]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][1] ),
        .O(\apbo[prdata][17]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][18]_INST_0 
       (.I0(\apbo[prdata][18]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][18] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][18] ),
        .O(\apbo[prdata] [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][18]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [2]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][18] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [8]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][2] ),
        .O(\apbo[prdata][18]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][19]_INST_0 
       (.I0(\apbo[prdata][19]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][19] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][19] ),
        .O(\apbo[prdata] [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][19]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [3]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][19] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [9]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][3] ),
        .O(\apbo[prdata][19]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][1]_INST_0 
       (.I0(\apbo[prdata][1]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][1]_INST_0_i_2_n_0 ),
        .O(\apbo[prdata] [1]),
        .S(\apbi[paddr] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8380FFFF83800000)) 
    \apbo[prdata][1]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][1] ),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I4(\apbi[paddr] [4]),
        .I5(\apbo[prdata][1]_INST_0_i_3_n_0 ),
        .O(\apbo[prdata][1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00B00080)) 
    \apbo[prdata][1]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][1] ),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [4]),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][33] ),
        .O(\apbo[prdata][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][1]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][33] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[status][tx_err_n_0_] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/p_6_in [1]),
        .O(\apbo[prdata][1]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][20]_INST_0 
       (.I0(\apbo[prdata][20]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][20] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][20] ),
        .O(\apbo[prdata] [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][20]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [4]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][20] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [10]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][4] ),
        .O(\apbo[prdata][20]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][21]_INST_0 
       (.I0(\apbo[prdata][21]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][21] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][21] ),
        .O(\apbo[prdata] [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][21]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [5]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][21] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [11]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][5] ),
        .O(\apbo[prdata][21]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][22]_INST_0 
       (.I0(\apbo[prdata][22]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][22] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][22] ),
        .O(\apbo[prdata] [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][22]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [6]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][22] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [12]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][6] ),
        .O(\apbo[prdata][22]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][23]_INST_0 
       (.I0(\apbo[prdata][23]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][23] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][23] ),
        .O(\apbo[prdata] [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][23]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [7]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][23] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [13]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][7] ),
        .O(\apbo[prdata][23]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][24]_INST_0 
       (.I0(\apbo[prdata][24]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][24] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][24] ),
        .O(\apbo[prdata] [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][24]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [8]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][24] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [14]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/p_1_in128_in ),
        .O(\apbo[prdata][24]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][25]_INST_0 
       (.I0(\apbo[prdata][25]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][25] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][25] ),
        .O(\apbo[prdata] [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][25]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [9]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][25] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [15]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][9] ),
        .O(\apbo[prdata][25]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][26]_INST_0 
       (.I0(\apbo[prdata][26]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][26] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][26] ),
        .O(\apbo[prdata] [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][26]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [10]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][26] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [16]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][10] ),
        .O(\apbo[prdata][26]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][27]_INST_0 
       (.I0(\apbo[prdata][27]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][27] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][27] ),
        .O(\apbo[prdata] [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][27]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [11]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][27] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [17]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][11] ),
        .O(\apbo[prdata][27]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF40)) 
    \apbo[prdata][28]_INST_0 
       (.I0(\apbi[paddr] [5]),
        .I1(\apbi[paddr] [4]),
        .I2(\apbo[prdata][28]_INST_0_i_1_n_0 ),
        .I3(\apbo[prdata][28]_INST_0_i_2_n_0 ),
        .O(\apbo[prdata] [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][28]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [12]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][28] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [18]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][12] ),
        .O(\apbo[prdata][28]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000C0000000A00F)) 
    \apbo[prdata][28]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][28] ),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][28] ),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][28]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][29]_INST_0 
       (.I0(\apbo[prdata][29]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][29] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][29] ),
        .O(\apbo[prdata] [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][29]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [13]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][29] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [19]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][13] ),
        .O(\apbo[prdata][29]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][2]_INST_0 
       (.I0(\apbo[prdata][2]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][2]_INST_0_i_2_n_0 ),
        .O(\apbo[prdata] [2]),
        .S(\apbi[paddr] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8380FFFF83800000)) 
    \apbo[prdata][2]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][2] ),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][linkfail_n_0_] ),
        .I4(\apbi[paddr] [4]),
        .I5(\apbo[prdata][2]_INST_0_i_3_n_0 ),
        .O(\apbo[prdata][2]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00B00080)) 
    \apbo[prdata][2]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][2] ),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [4]),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][34] ),
        .O(\apbo[prdata][2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][2]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][34] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[status][rx_int_n_0_] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/p_6_in [2]),
        .O(\apbo[prdata][2]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AAF0C000AA00C0)) 
    \apbo[prdata][30]_INST_0 
       (.I0(\apbo[prdata][30]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][30] ),
        .I2(\apbo[prdata][30]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .I5(\m100.u0/ethc0/r_reg[emacaddr_n_0_][30] ),
        .O(\apbo[prdata] [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][30]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [14]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][30] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [20]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][14] ),
        .O(\apbo[prdata][30]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \apbo[prdata][30]_INST_0_i_2 
       (.I0(\apbi[paddr] [2]),
        .I1(\apbi[paddr] [3]),
        .O(\apbo[prdata][30]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF40)) 
    \apbo[prdata][31]_INST_0 
       (.I0(\apbi[paddr] [5]),
        .I1(\apbi[paddr] [4]),
        .I2(\apbo[prdata][31]_INST_0_i_1_n_0 ),
        .I3(\apbo[prdata][31]_INST_0_i_2_n_0 ),
        .O(\apbo[prdata] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][31]_INST_0_i_1 
       (.I0(\m100.u0/ethc0/p_0_in0_in [15]),
        .I1(\m100.u0/ethc0/r_reg[rxdesc_n_0_][31] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdesc]__0 [21]),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][15] ),
        .O(\apbo[prdata][31]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000C0000000A00F)) 
    \apbo[prdata][31]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][31] ),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][31] ),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][31]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA808FFFFA8080000)) 
    \apbo[prdata][3]_INST_0 
       (.I0(\apbo[prdata][9]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][3] ),
        .I2(\apbo[prdata][10]_INST_0_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][35] ),
        .I4(\apbi[paddr] [5]),
        .I5(\apbo[prdata][3]_INST_0_i_1_n_0 ),
        .O(\apbo[prdata] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][3]_INST_0_i_1 
       (.I0(\apbo[prdata][3]_INST_0_i_2_n_0 ),
        .I1(\apbo[prdata][3]_INST_0_i_3_n_0 ),
        .O(\apbo[prdata][3]_INST_0_i_1_n_0 ),
        .S(\apbi[paddr] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][3]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][35] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[status][tx_int_n_0_] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/p_6_in [3]),
        .O(\apbo[prdata][3]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][3]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][3] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdsel_n_0_][3] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][busy]__0 ),
        .O(\apbo[prdata][3]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA808FFFFA8080000)) 
    \apbo[prdata][4]_INST_0 
       (.I0(\apbo[prdata][9]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][4] ),
        .I2(\apbo[prdata][10]_INST_0_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][36] ),
        .I4(\apbi[paddr] [5]),
        .I5(\apbo[prdata][4]_INST_0_i_1_n_0 ),
        .O(\apbo[prdata] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][4]_INST_0_i_1 
       (.I0(\apbo[prdata][4]_INST_0_i_2_n_0 ),
        .I1(\apbo[prdata][4]_INST_0_i_3_n_0 ),
        .O(\apbo[prdata][4]_INST_0_i_1_n_0 ),
        .S(\apbi[paddr] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][4]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][36] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[status][rxahberr_n_0_] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/p_6_in [4]),
        .O(\apbo[prdata][4]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \apbo[prdata][4]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][4] ),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [2]),
        .I4(\m100.u0/ethc0/r_reg[txdsel_n_0_][4] ),
        .O(\apbo[prdata][4]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA808FFFFA8080000)) 
    \apbo[prdata][5]_INST_0 
       (.I0(\apbo[prdata][9]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][5] ),
        .I2(\apbo[prdata][10]_INST_0_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][37] ),
        .I4(\apbi[paddr] [5]),
        .I5(\apbo[prdata][5]_INST_0_i_1_n_0 ),
        .O(\apbo[prdata] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][5]_INST_0_i_1 
       (.I0(\apbo[prdata][5]_INST_0_i_2_n_0 ),
        .I1(\apbo[prdata][5]_INST_0_i_3_n_0 ),
        .O(\apbo[prdata][5]_INST_0_i_1_n_0 ),
        .S(\apbi[paddr] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][5]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][37] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[status][txahberr_n_0_] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/p_6_in [5]),
        .O(\apbo[prdata][5]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFC0A0C0)) 
    \apbo[prdata][5]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][5] ),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [2]),
        .I4(\m100.u0/ethc0/r_reg[txdsel_n_0_][5] ),
        .O(\apbo[prdata][5]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA808FFFFA8080000)) 
    \apbo[prdata][6]_INST_0 
       (.I0(\apbo[prdata][9]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][6] ),
        .I2(\apbo[prdata][10]_INST_0_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][38] ),
        .I4(\apbi[paddr] [5]),
        .I5(\apbo[prdata][6]_INST_0_i_1_n_0 ),
        .O(\apbo[prdata] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][6]_INST_0_i_1 
       (.I0(\apbo[prdata][6]_INST_0_i_2_n_0 ),
        .I1(\apbo[prdata][6]_INST_0_i_3_n_0 ),
        .O(\apbo[prdata][6]_INST_0_i_1_n_0 ),
        .S(\apbi[paddr] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][6]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][6] ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][38] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[status][toosmall_n_0_] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/p_6_in [6]),
        .O(\apbo[prdata][6]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][6]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][6] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][6] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdsel_n_0_][6] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [0]),
        .O(\apbo[prdata][6]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA808FFFFA8080000)) 
    \apbo[prdata][7]_INST_0 
       (.I0(\apbo[prdata][9]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][7] ),
        .I2(\apbo[prdata][10]_INST_0_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][39] ),
        .I4(\apbi[paddr] [5]),
        .I5(\apbo[prdata][7]_INST_0_i_1_n_0 ),
        .O(\apbo[prdata] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][7]_INST_0_i_1 
       (.I0(\apbo[prdata][7]_INST_0_i_2_n_0 ),
        .I1(\apbo[prdata][7]_INST_0_i_3_n_0 ),
        .O(\apbo[prdata][7]_INST_0_i_1_n_0 ),
        .S(\apbi[paddr] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][7]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][39] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[status][invaddr_n_0_] ),
        .I4(\apbi[paddr] [2]),
        .I5(\etho[speed] ),
        .O(\apbo[prdata][7]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][7]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][7] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdsel_n_0_][7] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [1]),
        .O(\apbo[prdata][7]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][8]_INST_0 
       (.I0(\apbo[prdata][8]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][8]_INST_0_i_2_n_0 ),
        .O(\apbo[prdata] [8]),
        .S(\apbi[paddr] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB888B888888888)) 
    \apbo[prdata][8]_INST_0_i_1 
       (.I0(\apbo[prdata][8]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [4]),
        .I2(\m100.u0/ethc0/r_reg[mac_addr_n_0_][40] ),
        .I3(\apbi[paddr] [2]),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][8] ),
        .I5(\apbi[paddr] [3]),
        .O(\apbo[prdata][8]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00B00080)) 
    \apbo[prdata][8]_INST_0_i_2 
       (.I0(\m100.u0/ethc0/r_reg[emacaddr_n_0_][8] ),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [4]),
        .I4(\m100.u0/ethc0/r_reg[emacaddr_n_0_][40] ),
        .O(\apbo[prdata][8]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][8]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][8] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][8] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdsel_n_0_][8] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [2]),
        .O(\apbo[prdata][8]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA808FFFFA8080000)) 
    \apbo[prdata][9]_INST_0 
       (.I0(\apbo[prdata][9]_INST_0_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[emacaddr_n_0_][9] ),
        .I2(\apbo[prdata][10]_INST_0_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[emacaddr_n_0_][41] ),
        .I4(\apbi[paddr] [5]),
        .I5(\apbo[prdata][9]_INST_0_i_2_n_0 ),
        .O(\apbo[prdata] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \apbo[prdata][9]_INST_0_i_1 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[paddr] [4]),
        .O(\apbo[prdata][9]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][9]_INST_0_i_2 
       (.I0(\apbo[prdata][9]_INST_0_i_3_n_0 ),
        .I1(\apbo[prdata][9]_INST_0_i_4_n_0 ),
        .O(\apbo[prdata][9]_INST_0_i_2_n_0 ),
        .S(\apbi[paddr] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF101F0F0F1010000)) 
    \apbo[prdata][9]_INST_0_i_3 
       (.I0(\m100.u0/ethc0/r_reg[etxidle]__0 ),
        .I1(\m100.u0/ethc0/r_reg[erxidle]__0 ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][9] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mac_addr_n_0_][41] ),
        .O(\apbo[prdata][9]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \apbo[prdata][9]_INST_0_i_4 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][9] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][9] ),
        .I2(\apbi[paddr] [3]),
        .I3(\m100.u0/ethc0/r_reg[txdsel_n_0_][9] ),
        .I4(\apbi[paddr] [2]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [3]),
        .O(\apbo[prdata][9]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \etho[reset]_INST_0 
       (.I0(rst),
        .I1(\m100.u0/ethc0/p_6_in [6]),
        .O(\etho[reset] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFA8A8A8AA)) 
    \gmiimode0.r[act]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[en]__0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[enold]__0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero]__0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/v ),
        .O(\gmiimode0.r ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB08080B0B08080)) 
    \gmiimode0.r[byte_count][0]_i_1 
       (.I0(\gmiimode0.r_reg[byte_count][3]_i_2_n_7 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \gmiimode0.r[byte_count][0]_i_1__0 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .O(\gmiimode0.r[byte_count][0]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000033335115)) 
    \gmiimode0.r[byte_count][10]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I2(\m100.u0/ethc0/rxo[write] ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[write_ack] ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\gmiimode0.r[byte_count][10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000028)) 
    \gmiimode0.r[byte_count][10]_i_1__0 
       (.I0(\gmiimode0.r[byte_count][10]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[deferring_n_0_] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .O(\gmiimode0.r[byte_count][10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000C0F0200000002)) 
    \gmiimode0.r[byte_count][10]_i_2 
       (.I0(\gmiimode0.r[byte_count][10]_i_4__0_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I5(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .O(\gmiimode0.r[byte_count][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFB800)) 
    \gmiimode0.r[byte_count][10]_i_2__0 
       (.I0(\gmiimode0.r_reg [2]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [10]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\gmiimode0.r[byte_count][10]_i_4_n_0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \gmiimode0.r[byte_count][10]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\gmiimode0.r[byte_count][10]_i_5_n_0 ),
        .O(\gmiimode0.r[byte_count][10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8888828800000000)) 
    \gmiimode0.r[byte_count][10]_i_4 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [10]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [9]),
        .I3(\gmiimode0.r[byte_count][10]_i_8_n_0 ),
        .I4(\m100.u0/ethc0/rxo[byte_count] [8]),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .O(\gmiimode0.r[byte_count][10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \gmiimode0.r[byte_count][10]_i_4__0 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[deferring_n_0_] ),
        .O(\gmiimode0.r[byte_count][10]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9555555555555555)) 
    \gmiimode0.r[byte_count][10]_i_5 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][10] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][8] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][6] ),
        .I3(\gmiimode0.r[byte_count][10]_i_6_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][7] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][9] ),
        .O(\gmiimode0.r[byte_count][10]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \gmiimode0.r[byte_count][10]_i_6 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][5] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .O(\gmiimode0.r[byte_count][10]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \gmiimode0.r[byte_count][10]_i_8 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [4]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [5]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [7]),
        .I5(\m100.u0/ethc0/rxo[byte_count] [6]),
        .O(\gmiimode0.r[byte_count][10]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0440)) 
    \gmiimode0.r[byte_count][1]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .O(\gmiimode0.r[byte_count][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB08080B0B08080)) 
    \gmiimode0.r[byte_count][1]_i_1__0 
       (.I0(\gmiimode0.r_reg[byte_count][3]_i_2_n_6 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h04404040)) 
    \gmiimode0.r[byte_count][2]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .O(\gmiimode0.r[byte_count][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF8BB80000)) 
    \gmiimode0.r[byte_count][2]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_1_in6_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I3(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I5(\gmiimode0.r[byte_count][2]_i_2_n_0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \gmiimode0.r[byte_count][2]_i_2 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .O(\gmiimode0.r[byte_count][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFCFFB800)) 
    \gmiimode0.r[byte_count][3]_i_1 
       (.I0(\gmiimode0.r_reg[byte_count][3]_i_2_n_4 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\gmiimode0.r[byte_count][3]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\gmiimode0.r[byte_count][3]_i_4_n_0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0444444440000000)) 
    \gmiimode0.r[byte_count][3]_i_1__0 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .O(\gmiimode0.r[byte_count][3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0F00FF8)) 
    \gmiimode0.r[byte_count][3]_i_3 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I4(\m100.u0/ethc0/rxo[byte_count] [2]),
        .O(\gmiimode0.r[byte_count][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8200)) 
    \gmiimode0.r[byte_count][3]_i_4 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .O(\gmiimode0.r[byte_count][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6AAA6AAA6AAAAAAA)) 
    \gmiimode0.r[byte_count][3]_i_8 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dv]__0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[en]__0 ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero]__0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .O(\gmiimode0.r[byte_count][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    \gmiimode0.r[byte_count][4]_i_1 
       (.I0(\gmiimode0.r[byte_count][6]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ),
        .O(\gmiimode0.r[byte_count][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFCFFB800)) 
    \gmiimode0.r[byte_count][4]_i_1__0 
       (.I0(\gmiimode0.r_reg[byte_count][7]_i_2_n_7 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\gmiimode0.r[byte_count][4]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\gmiimode0.r[byte_count][4]_i_3_n_0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFF55000000EA)) 
    \gmiimode0.r[byte_count][4]_i_2 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I5(\m100.u0/ethc0/rxo[byte_count] [4]),
        .O(\gmiimode0.r[byte_count][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88820000)) 
    \gmiimode0.r[byte_count][4]_i_3 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [4]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .O(\gmiimode0.r[byte_count][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \gmiimode0.r[byte_count][5]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [5]),
        .O(\gmiimode0.r[byte_count][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFB800)) 
    \gmiimode0.r[byte_count][5]_i_1__0 
       (.I0(\gmiimode0.r_reg[byte_count][7]_i_2_n_6 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\gmiimode0.r[byte_count][5]_i_2__0_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\gmiimode0.r[byte_count][5]_i_3_n_0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    \gmiimode0.r[byte_count][5]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][5] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFD0002)) 
    \gmiimode0.r[byte_count][5]_i_2__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I1(\m100.u0/ethc0/rxo[byte_count] [4]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [5]),
        .O(\gmiimode0.r[byte_count][5]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAA8000200000000)) 
    \gmiimode0.r[byte_count][5]_i_3 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [4]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [5]),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .O(\gmiimode0.r[byte_count][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    \gmiimode0.r[byte_count][6]_i_1 
       (.I0(\gmiimode0.r[byte_count][6]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][5] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ),
        .I4(\gmiimode0.r[byte_count][6]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][6] ),
        .O(\gmiimode0.r[byte_count][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFB800)) 
    \gmiimode0.r[byte_count][6]_i_1__0 
       (.I0(\gmiimode0.r_reg[byte_count][7]_i_2_n_5 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\gmiimode0.r[byte_count][6]_i_2__0_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\gmiimode0.r[byte_count][6]_i_3__0_n_0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \gmiimode0.r[byte_count][6]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .O(\gmiimode0.r[byte_count][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCCCCCCCCCCCCC6)) 
    \gmiimode0.r[byte_count][6]_i_2__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I1(\m100.u0/ethc0/rxo[byte_count] [6]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [4]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I5(\m100.u0/ethc0/rxo[byte_count] [5]),
        .O(\gmiimode0.r[byte_count][6]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \gmiimode0.r[byte_count][6]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .O(\gmiimode0.r[byte_count][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2800)) 
    \gmiimode0.r[byte_count][6]_i_3__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [6]),
        .I2(\gmiimode0.r[byte_count][9]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .O(\gmiimode0.r[byte_count][6]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \gmiimode0.r[byte_count][7]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [7]),
        .O(\gmiimode0.r[byte_count][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFCFFB800)) 
    \gmiimode0.r[byte_count][7]_i_1__0 
       (.I0(\gmiimode0.r_reg[byte_count][7]_i_2_n_4 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\gmiimode0.r[byte_count][7]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\gmiimode0.r[byte_count][7]_i_4_n_0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    \gmiimode0.r[byte_count][7]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][7] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][5] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ),
        .I4(\gmiimode0.r[byte_count][6]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][6] ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF0FFFFF00F80000)) 
    \gmiimode0.r[byte_count][7]_i_3 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I3(\m100.u0/ethc0/rxo[byte_count] [6]),
        .I4(\gmiimode0.r[byte_count][9]_i_4_n_0 ),
        .I5(\m100.u0/ethc0/rxo[byte_count] [7]),
        .O(\gmiimode0.r[byte_count][7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88280000)) 
    \gmiimode0.r[byte_count][7]_i_4 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [7]),
        .I2(\gmiimode0.r[byte_count][9]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/rxo[byte_count] [6]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .O(\gmiimode0.r[byte_count][7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \gmiimode0.r[byte_count][8]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [8]),
        .O(\gmiimode0.r[byte_count][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFB800)) 
    \gmiimode0.r[byte_count][8]_i_1__0 
       (.I0(\gmiimode0.r_reg [0]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\gmiimode0.r[byte_count][8]_i_2__0_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\gmiimode0.r[byte_count][8]_i_3_n_0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \gmiimode0.r[byte_count][8]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][8] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][6] ),
        .I2(\gmiimode0.r[byte_count][10]_i_6_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][7] ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCC6CCCC)) 
    \gmiimode0.r[byte_count][8]_i_2__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I1(\m100.u0/ethc0/rxo[byte_count] [8]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [6]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [7]),
        .I4(\gmiimode0.r[byte_count][9]_i_4_n_0 ),
        .O(\gmiimode0.r[byte_count][8]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8882888800000000)) 
    \gmiimode0.r[byte_count][8]_i_3 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [8]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [6]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [7]),
        .I4(\gmiimode0.r[byte_count][9]_i_4_n_0 ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .O(\gmiimode0.r[byte_count][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \gmiimode0.r[byte_count][9]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [9]),
        .O(\gmiimode0.r[byte_count][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFB800)) 
    \gmiimode0.r[byte_count][9]_i_1__0 
       (.I0(\gmiimode0.r_reg [1]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\gmiimode0.r[byte_count][9]_i_2__0_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\gmiimode0.r[byte_count][9]_i_3_n_0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \gmiimode0.r[byte_count][9]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][9] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][7] ),
        .I2(\gmiimode0.r[byte_count][10]_i_6_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][6] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][8] ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCCCCCCCCCCC6CC)) 
    \gmiimode0.r[byte_count][9]_i_2__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I1(\m100.u0/ethc0/rxo[byte_count] [9]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [8]),
        .I3(\gmiimode0.r[byte_count][9]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/rxo[byte_count] [7]),
        .I5(\m100.u0/ethc0/rxo[byte_count] [6]),
        .O(\gmiimode0.r[byte_count][9]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h82880000)) 
    \gmiimode0.r[byte_count][9]_i_3 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [9]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [8]),
        .I3(\gmiimode0.r[byte_count][10]_i_8_n_0 ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .O(\gmiimode0.r[byte_count][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \gmiimode0.r[byte_count][9]_i_4 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [5]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [4]),
        .O(\gmiimode0.r[byte_count][9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00005502)) 
    \gmiimode0.r[cnt][0]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[cnt] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \gmiimode0.r[cnt][0]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[cnt] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0069FFFF006941FF)) 
    \gmiimode0.r[cnt][1]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[cnt] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT4 #(
    .INIT(16'hF00E)) 
    \gmiimode0.r[cnt][1]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[cnt] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0CFF0C4F)) 
    \gmiimode0.r[cnt][2]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I1(\gmiimode0.r[cnt][2]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[cnt] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT4 #(
    .INIT(16'hFC02)) 
    \gmiimode0.r[cnt][2]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[cnt] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF8F007070FF8F00)) 
    \gmiimode0.r[cnt][2]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I3(\gmiimode0.r[cnt][3]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .O(\gmiimode0.r[cnt][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF290100002901)) 
    \gmiimode0.r[cnt][3]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I3(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[cnt][3]_i_3_n_0 ),
        .O(\gmiimode0.r[cnt][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000001)) 
    \gmiimode0.r[cnt][3]_i_10 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][10] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][8] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][6] ),
        .I3(\gmiimode0.r[byte_count][10]_i_6_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][7] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][9] ),
        .O(\gmiimode0.r[cnt][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \gmiimode0.r[cnt][3]_i_11 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .O(\gmiimode0.r[cnt][3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT4 #(
    .INIT(16'hAAA9)) 
    \gmiimode0.r[cnt][3]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[cnt] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2802)) 
    \gmiimode0.r[cnt][3]_i_2 
       (.I0(\gmiimode0.r[cnt][3]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[cnt] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBAAAAAAAAAAAAAAA)) 
    \gmiimode0.r[cnt][3]_i_3 
       (.I0(\gmiimode0.r[cnt][3]_i_5_n_0 ),
        .I1(\gmiimode0.r[tx_en]_i_5_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I4(\gmiimode0.r_reg[tx_en]_i_7_n_0 ),
        .I5(\gmiimode0.r[cnt][3]_i_6_n_0 ),
        .O(\gmiimode0.r[cnt][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFDC002FFFFFFFF)) 
    \gmiimode0.r[cnt][3]_i_4 
       (.I0(\gmiimode0.r[cnt][3]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I2(\gmiimode0.r[cnt][3]_i_8_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][3] ),
        .I5(\gmiimode0.r[start][1]_i_2_n_0 ),
        .O(\gmiimode0.r[cnt][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000004040000FF00)) 
    \gmiimode0.r[cnt][3]_i_5 
       (.I0(\gmiimode0.r[cnt][3]_i_9_n_0 ),
        .I1(\gmiimode0.r[cnt][3]_i_10_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I3(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .O(\gmiimode0.r[cnt][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h80080000FFFFFFFF)) 
    \gmiimode0.r[cnt][3]_i_6 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .I3(\gmiimode0.r[cnt][3]_i_11_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][5] ),
        .I5(\gmiimode0.r[cnt][3]_i_10_n_0 ),
        .O(\gmiimode0.r[cnt][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \gmiimode0.r[cnt][3]_i_7 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .O(\gmiimode0.r[cnt][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7000000070707070)) 
    \gmiimode0.r[cnt][3]_i_8 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .O(\gmiimode0.r[cnt][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFF7FFFFFFFFF)) 
    \gmiimode0.r[cnt][3]_i_9 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .I4(\gmiimode0.r[cnt][3]_i_11_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][5] ),
        .O(\gmiimode0.r[cnt][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F203F3F3F202020)) 
    \gmiimode0.r[crc][0]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\gmiimode0.r[crc][31]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][0] ),
        .I4(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I5(\gmiimode0.r[crc][0]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT4 #(
    .INIT(16'h6F60)) 
    \gmiimode0.r[crc][0]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \gmiimode0.r[crc][0]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ),
        .I1(\^etho[txd] [3]),
        .O(\gmiimode0.r[crc][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][10]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][10]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \gmiimode0.r[crc][10]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][6] ),
        .I1(\gmiimode0.r[crc][13]_i_2__0_n_0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \gmiimode0.r[crc][10]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][10] ),
        .I1(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_12_in ),
        .I3(\gmiimode0.r[crc][13]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ),
        .I5(\^etho[txd] [3]),
        .O(\gmiimode0.r[crc][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][11]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][11]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT4 #(
    .INIT(16'h6F60)) 
    \gmiimode0.r[crc][11]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_13_in ),
        .I1(\gmiimode0.r[crc][11]_i_2__0_n_0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h2AEAEA2A)) 
    \gmiimode0.r[crc][11]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_17_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_13_in ),
        .I4(\gmiimode0.r[crc][11]_i_3_n_0 ),
        .O(\gmiimode0.r[crc][11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \gmiimode0.r[crc][11]_i_2__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in10_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in15_in ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .O(\gmiimode0.r[crc][11]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \gmiimode0.r[crc][11]_i_3 
       (.I0(\^etho[txd] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in10_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ),
        .I3(\^etho[txd] [3]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ),
        .I5(\^etho[txd] [2]),
        .O(\gmiimode0.r[crc][11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][12]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][12]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \gmiimode0.r[crc][12]_i_1__0 
       (.I0(\gmiimode0.r[crc][24]_i_2__0_n_0 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_14_in ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \gmiimode0.r[crc][12]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][12] ),
        .I1(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_14_in ),
        .I3(\gmiimode0.r[crc][12]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ),
        .I5(\^etho[txd] [3]),
        .O(\gmiimode0.r[crc][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \gmiimode0.r[crc][12]_i_3 
       (.I0(\^etho[txd] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .I2(\^etho[txd] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ),
        .O(\gmiimode0.r[crc][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][13]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][13]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \gmiimode0.r[crc][13]_i_1__0 
       (.I0(\gmiimode0.r[crc][13]_i_2__0_n_0 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in15_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_15_in ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \gmiimode0.r[crc][13]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][13] ),
        .I1(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][9] ),
        .I3(\gmiimode0.r[crc][13]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ),
        .I5(\^etho[txd] [2]),
        .O(\gmiimode0.r[crc][13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \gmiimode0.r[crc][13]_i_2__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in10_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in12_in ),
        .O(\gmiimode0.r[crc][13]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \gmiimode0.r[crc][13]_i_3 
       (.I0(\^etho[txd] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .I2(\^etho[txd] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in10_in ),
        .O(\gmiimode0.r[crc][13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][14]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][14]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \gmiimode0.r[crc][14]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_16_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in12_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .I3(\gmiimode0.r[crc][25]_i_2__0_n_0 ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \gmiimode0.r[crc][14]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][14] ),
        .I1(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][10] ),
        .I3(\gmiimode0.r[crc][25]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .I5(\^etho[txd] [1]),
        .O(\gmiimode0.r[crc][14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][15]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][15]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \gmiimode0.r[crc][15]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_17_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in10_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEA2A2AEA2AEAEA2A)) 
    \gmiimode0.r[crc][15]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_22_in55_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_17_in ),
        .I4(\^etho[txd] [0]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in10_in ),
        .O(\gmiimode0.r[crc][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][16]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][16]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \gmiimode0.r[crc][16]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_18_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEA2A2AEA2AEAEA2A)) 
    \gmiimode0.r[crc][16]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_31_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][12] ),
        .I4(\^etho[txd] [3]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ),
        .O(\gmiimode0.r[crc][16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][17]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][17]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \gmiimode0.r[crc][17]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_19_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in15_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEA2A2AEA2AEAEA2A)) 
    \gmiimode0.r[crc][17]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_32_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][13] ),
        .I4(\^etho[txd] [2]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ),
        .O(\gmiimode0.r[crc][17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][18]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][18]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \gmiimode0.r[crc][18]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_20_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in12_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEA2A2AEA2AEAEA2A)) 
    \gmiimode0.r[crc][18]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_23_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][14] ),
        .I4(\^etho[txd] [1]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .O(\gmiimode0.r[crc][18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][19]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][19]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \gmiimode0.r[crc][19]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_22_in55_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in10_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEA2A2AEA2AEAEA2A)) 
    \gmiimode0.r[crc][19]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_24_in59_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_22_in55_in ),
        .I4(\^etho[txd] [0]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in10_in ),
        .O(\gmiimode0.r[crc][19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F203F3F3F202020)) 
    \gmiimode0.r[crc][1]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\gmiimode0.r[crc][31]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][1] ),
        .I4(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I5(\gmiimode0.r[crc][1]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \gmiimode0.r[crc][1]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in15_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \gmiimode0.r[crc][1]_i_2 
       (.I0(\^etho[txd] [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ),
        .I2(\^etho[txd] [3]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ),
        .O(\gmiimode0.r[crc][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F203F3F3F202020)) 
    \gmiimode0.r[crc][20]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\gmiimode0.r[crc][31]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_25_in ),
        .I4(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_31_in ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF00FF00BF00)) 
    \gmiimode0.r[crc][20]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_31_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F203F3F3F202020)) 
    \gmiimode0.r[crc][21]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\gmiimode0.r[crc][31]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_26_in64_in ),
        .I4(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_32_in ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF00FF00BF00)) 
    \gmiimode0.r[crc][21]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_32_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][22]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][22]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \gmiimode0.r[crc][22]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_23_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEA2A2AEA2AEAEA2A)) 
    \gmiimode0.r[crc][22]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_27_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_23_in ),
        .I4(\^etho[txd] [3]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ),
        .O(\gmiimode0.r[crc][22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][23]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][23]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \gmiimode0.r[crc][23]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in15_in ),
        .I2(\gmiimode0.r[crc][26]_i_2__0_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_24_in59_in ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \gmiimode0.r[crc][23]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_28_in69_in ),
        .I1(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_24_in59_in ),
        .I3(\gmiimode0.r[crc][0]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ),
        .I5(\^etho[txd] [2]),
        .O(\gmiimode0.r[crc][23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][24]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][24]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT4 #(
    .INIT(16'h6F60)) 
    \gmiimode0.r[crc][24]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_25_in ),
        .I1(\gmiimode0.r[crc][24]_i_2__0_n_0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \gmiimode0.r[crc][24]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][24] ),
        .I1(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_25_in ),
        .I3(\gmiimode0.r[crc][24]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .I5(\^etho[txd] [1]),
        .O(\gmiimode0.r[crc][24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \gmiimode0.r[crc][24]_i_2__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in12_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in15_in ),
        .O(\gmiimode0.r[crc][24]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \gmiimode0.r[crc][24]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ),
        .I1(\^etho[txd] [2]),
        .O(\gmiimode0.r[crc][24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][25]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][25]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \gmiimode0.r[crc][25]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_26_in64_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in12_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .I3(\gmiimode0.r[crc][25]_i_2__0_n_0 ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \gmiimode0.r[crc][25]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_30_in72_in ),
        .I1(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_26_in64_in ),
        .I3(\gmiimode0.r[crc][25]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .I5(\^etho[txd] [1]),
        .O(\gmiimode0.r[crc][25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \gmiimode0.r[crc][25]_i_2__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in10_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .O(\gmiimode0.r[crc][25]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \gmiimode0.r[crc][25]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in10_in ),
        .I1(\^etho[txd] [0]),
        .O(\gmiimode0.r[crc][25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][26]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][26]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \gmiimode0.r[crc][26]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in10_in ),
        .I2(\gmiimode0.r[crc][26]_i_2__0_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_27_in ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \gmiimode0.r[crc][26]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_33_in ),
        .I1(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I2(\^etho[txd] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in10_in ),
        .I4(\gmiimode0.r[crc][0]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_27_in ),
        .O(\gmiimode0.r[crc][26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \gmiimode0.r[crc][26]_i_2__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .O(\gmiimode0.r[crc][26]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][27]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][27]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \gmiimode0.r[crc][27]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_28_in69_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in15_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEA2A2AEA2AEAEA2A)) 
    \gmiimode0.r[crc][27]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][27] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_28_in69_in ),
        .I4(\^etho[txd] [2]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ),
        .O(\gmiimode0.r[crc][27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000002003FFFFFFF)) 
    \gmiimode0.r[crc][28]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][28]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \gmiimode0.r[crc][28]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_29_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in12_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3CC3555555555555)) 
    \gmiimode0.r[crc][28]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][24] ),
        .I2(\^etho[txd] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .O(\gmiimode0.r[crc][28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000002003FFFFFFF)) 
    \gmiimode0.r[crc][29]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][29]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \gmiimode0.r[crc][29]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_30_in72_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in10_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3CC3555555555555)) 
    \gmiimode0.r[crc][29]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_30_in72_in ),
        .I2(\^etho[txd] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in10_in ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .O(\gmiimode0.r[crc][29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000080)) 
    \gmiimode0.r[crc][29]_i_2__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F2020203F203F3F)) 
    \gmiimode0.r[crc][2]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\gmiimode0.r[crc][31]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_8_in ),
        .I4(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I5(\gmiimode0.r[crc][2]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \gmiimode0.r[crc][2]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .I2(\gmiimode0.r[crc][24]_i_2__0_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9669699669969669)) 
    \gmiimode0.r[crc][2]_i_2 
       (.I0(\^etho[txd] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ),
        .I3(\^etho[txd] [2]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .I5(\^etho[txd] [1]),
        .O(\gmiimode0.r[crc][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F203F3F3F202020)) 
    \gmiimode0.r[crc][30]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\gmiimode0.r[crc][31]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .I4(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_33_in ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF00FF00BF00)) 
    \gmiimode0.r[crc][30]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_33_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F203F3F3F202020)) 
    \gmiimode0.r[crc][31]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\gmiimode0.r[crc][31]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in10_in ),
        .I4(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][27] ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000001000100)) 
    \gmiimode0.r[crc][31]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .O(\gmiimode0.r[crc][31]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8010)) 
    \gmiimode0.r[crc][31]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\gmiimode0.r[crc][31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF00FF00BF00)) 
    \gmiimode0.r[crc][31]_i_2__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][27] ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \gmiimode0.r[crc][31]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .O(\gmiimode0.r[crc][31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F203F3F3F202020)) 
    \gmiimode0.r[crc][3]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\gmiimode0.r[crc][31]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_9_in ),
        .I4(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I5(\gmiimode0.r[crc][3]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96FF9600)) 
    \gmiimode0.r[crc][3]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in10_in ),
        .I2(\gmiimode0.r[crc][24]_i_2__0_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996966996696996)) 
    \gmiimode0.r[crc][3]_i_2 
       (.I0(\^etho[txd] [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in10_in ),
        .I3(\^etho[txd] [0]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .I5(\^etho[txd] [1]),
        .O(\gmiimode0.r[crc][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][4]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][4]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \gmiimode0.r[crc][4]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][0] ),
        .I1(\gmiimode0.r[crc][13]_i_2__0_n_0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \gmiimode0.r[crc][4]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_10_in ),
        .I1(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][0] ),
        .I3(\gmiimode0.r[crc][13]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ),
        .I5(\^etho[txd] [3]),
        .O(\gmiimode0.r[crc][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][5]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][5]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT4 #(
    .INIT(16'h6F60)) 
    \gmiimode0.r[crc][5]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][1] ),
        .I1(\gmiimode0.r[crc][11]_i_2__0_n_0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h2AEAEA2A)) 
    \gmiimode0.r[crc][5]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_11_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][1] ),
        .I4(\gmiimode0.r[crc][11]_i_3_n_0 ),
        .O(\gmiimode0.r[crc][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][6]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][6]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT4 #(
    .INIT(16'h6F60)) 
    \gmiimode0.r[crc][6]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][2] ),
        .I1(\gmiimode0.r[crc][24]_i_2__0_n_0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \gmiimode0.r[crc][6]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_12_in ),
        .I1(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_8_in ),
        .I3(\gmiimode0.r[crc][24]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .I5(\^etho[txd] [1]),
        .O(\gmiimode0.r[crc][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][7]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][7]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6996FFFF69960000)) 
    \gmiimode0.r[crc][7]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_9_in ),
        .I1(\gmiimode0.r[crc][13]_i_2__0_n_0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \gmiimode0.r[crc][7]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_13_in ),
        .I1(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_9_in ),
        .I3(\gmiimode0.r[crc][13]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ),
        .I5(\^etho[txd] [3]),
        .O(\gmiimode0.r[crc][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][8]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][8]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6F60)) 
    \gmiimode0.r[crc][8]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_10_in ),
        .I1(\gmiimode0.r[crc][11]_i_2__0_n_0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h2AEAEA2A)) 
    \gmiimode0.r[crc][8]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_14_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_10_in ),
        .I4(\gmiimode0.r[crc][11]_i_3_n_0 ),
        .O(\gmiimode0.r[crc][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFF00000200)) 
    \gmiimode0.r[crc][9]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I5(\gmiimode0.r[crc][9]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6F60)) 
    \gmiimode0.r[crc][9]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_11_in ),
        .I1(\gmiimode0.r[crc][24]_i_2__0_n_0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/crc_en ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BB8B88BB88B8BB8)) 
    \gmiimode0.r[crc][9]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][9] ),
        .I1(\gmiimode0.r[crc][31]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_11_in ),
        .I3(\gmiimode0.r[crc][24]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .I5(\^etho[txd] [1]),
        .O(\gmiimode0.r[crc][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFDBFFFFF00040000)) 
    \gmiimode0.r[crc_en]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I4(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .O(\gmiimode0.r[crc_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hC8C0)) 
    \gmiimode0.r[crs_act]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_act]__1 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/txrst ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/rin ),
        .O(\gmiimode0.r[crs_act]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \gmiimode0.r[data][11]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I2(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I4(\gmiimode0.r[data][27]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \gmiimode0.r[data][15]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I2(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I4(\gmiimode0.r[data][31]_i_2__0_n_0 ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \gmiimode0.r[data][19]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I4(\gmiimode0.r[data][27]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \gmiimode0.r[data][23]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I4(\gmiimode0.r[data][31]_i_2__0_n_0 ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    \gmiimode0.r[data][27]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I4(\gmiimode0.r[data][27]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \gmiimode0.r[data][27]_i_2 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .O(\gmiimode0.r[data][27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000004000C000)) 
    \gmiimode0.r[data][31]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_28_out ),
        .I3(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I4(\gmiimode0.r[data][31]_i_2_n_0 ),
        .I5(\gmiimode0.r[tx_en]_i_5_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    \gmiimode0.r[data][31]_i_1__0 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I4(\gmiimode0.r[data][31]_i_2__0_n_0 ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \gmiimode0.r[data][31]_i_2 
       (.I0(\gmiimode0.r_reg[tx_en]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .O(\gmiimode0.r[data][31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \gmiimode0.r[data][31]_i_2__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .O(\gmiimode0.r[data][31]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \gmiimode0.r[data][3]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I2(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I4(\gmiimode0.r[data][27]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \gmiimode0.r[data][7]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I2(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I4(\gmiimode0.r[data][31]_i_2__0_n_0 ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0082)) 
    \gmiimode0.r[dataout][31]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/write_req ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[write_ack] ),
        .I2(\m100.u0/ethc0/rxo[write] ),
        .I3(\m100.u0/ethc0/rxo[status] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFBBFF00000030)) 
    \gmiimode0.r[deferring]_i_1 
       (.I0(\gmiimode0.r[ifg_cycls][7]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_5_out ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [2]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[deferring_n_0_] ),
        .O(\gmiimode0.r[deferring]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB888B8B8)) 
    \gmiimode0.r[deferring]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[transmitting]__0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in38_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/rin ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_prev_n_0_] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_act]__1 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/p_5_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \gmiimode0.r[delay_val][0]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/v [0]),
        .O(\gmiimode0.r[delay_val][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h009F0090)) 
    \gmiimode0.r[delay_val][1]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/v [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\gmiimode0.r[delay_val][1]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFE00000000)) 
    \gmiimode0.r[delay_val][1]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][1] ),
        .O(\gmiimode0.r[delay_val][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000A9FF0000A900)) 
    \gmiimode0.r[delay_val][2]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/v [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/v [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I5(\gmiimode0.r[delay_val][2]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFE0000)) 
    \gmiimode0.r[delay_val][2]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_1_in75_in ),
        .O(\gmiimode0.r[delay_val][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h009F0090)) 
    \gmiimode0.r[delay_val][3]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [3]),
        .I1(\gmiimode0.r[delay_val][3]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\gmiimode0.r[delay_val][3]_i_3_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \gmiimode0.r[delay_val][3]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/v [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/v [2]),
        .O(\gmiimode0.r[delay_val][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEEE00000000)) 
    \gmiimode0.r[delay_val][3]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_5_in ),
        .O(\gmiimode0.r[delay_val][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h009F0090)) 
    \gmiimode0.r[delay_val][4]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [4]),
        .I1(\gmiimode0.r[delay_val][4]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\gmiimode0.r[delay_val][4]_i_3_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \gmiimode0.r[delay_val][4]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/v [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/v [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/v [3]),
        .O(\gmiimode0.r[delay_val][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \gmiimode0.r[delay_val][4]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_7_in ),
        .O(\gmiimode0.r[delay_val][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h009F0090)) 
    \gmiimode0.r[delay_val][5]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [5]),
        .I1(\gmiimode0.r[delay_val][5]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\gmiimode0.r[delay_val][5]_i_3_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \gmiimode0.r[delay_val][5]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/v [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/v [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/v [2]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/v [4]),
        .O(\gmiimode0.r[delay_val][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFEEEA00000000)) 
    \gmiimode0.r[delay_val][5]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][5] ),
        .O(\gmiimode0.r[delay_val][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h009F0090)) 
    \gmiimode0.r[delay_val][6]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [6]),
        .I1(\gmiimode0.r[delay_val][7]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\gmiimode0.r[delay_val][6]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEA0000)) 
    \gmiimode0.r[delay_val][6]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][6] ),
        .O(\gmiimode0.r[delay_val][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000A9FF0000A900)) 
    \gmiimode0.r[delay_val][7]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [7]),
        .I1(\gmiimode0.r[delay_val][7]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/v [6]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I5(\gmiimode0.r[delay_val][7]_i_3_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \gmiimode0.r[delay_val][7]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [4]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/v [2]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/v [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/v [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/v [3]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/v [5]),
        .O(\gmiimode0.r[delay_val][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFEAAA00000000)) 
    \gmiimode0.r[delay_val][7]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][7] ),
        .O(\gmiimode0.r[delay_val][7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h009F0090)) 
    \gmiimode0.r[delay_val][8]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [8]),
        .I1(\gmiimode0.r[delay_val][8]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\gmiimode0.r[delay_val][8]_i_3_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \gmiimode0.r[delay_val][8]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [6]),
        .I1(\gmiimode0.r[delay_val][7]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/v [7]),
        .O(\gmiimode0.r[delay_val][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE0)) 
    \gmiimode0.r[delay_val][8]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][8] ),
        .O(\gmiimode0.r[delay_val][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040004000404040)) 
    \gmiimode0.r[delay_val][9]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][6] ),
        .I5(\gmiimode0.r[delay_val][9]_i_3_n_0 ),
        .O(\gmiimode0.r[delay_val][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h009F0090)) 
    \gmiimode0.r[delay_val][9]_i_2 
       (.I0(\gmiimode0.r[delay_val][9]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/v [9]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\gmiimode0.r[delay_val][9]_i_5_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \gmiimode0.r[delay_val][9]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][2] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][3] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][5] ),
        .O(\gmiimode0.r[delay_val][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \gmiimode0.r[delay_val][9]_i_4 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v [7]),
        .I1(\gmiimode0.r[delay_val][7]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/v [6]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/v [8]),
        .O(\gmiimode0.r[delay_val][9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFEAAAA00000000)) 
    \gmiimode0.r[delay_val][9]_i_5 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in74_in ),
        .O(\gmiimode0.r[delay_val][9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF7F0080)) 
    \gmiimode0.r[done]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I4(\m100.u0/ethc0/txo ),
        .O(\gmiimode0.r[done]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBAAFBFF04550400)) 
    \gmiimode0.r[done]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\gmiimode0.r[done]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/rxo ),
        .O(\gmiimode0.r[done]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3404043404040404)) 
    \gmiimode0.r[done]_i_2 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[write_ack] ),
        .I4(\m100.u0/ethc0/rxo[write] ),
        .I5(\FSM_sequential_gmiimode0.r[rx_state][0]_i_3_n_0 ),
        .O(\gmiimode0.r[done]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000444A0000)) 
    \gmiimode0.r[dv]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dv]__0 ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero]__0 ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/rxrst ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/v ),
        .O(\gmiimode0.r[dv]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \gmiimode0.r[enold]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[en]__0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero]__0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[enold]__0 ),
        .O(\gmiimode0.r[enold]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFAFE00000A02)) 
    \gmiimode0.r[got4b]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/v[got4b] ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .O(\gmiimode0.r[got4b]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF6F0F600000000)) 
    \gmiimode0.r[got4b]_i_2 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/p_1_in6_in ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[got4b] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEE00002204)) 
    \gmiimode0.r[gotframe]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .I5(\m100.u0/ethc0/rxo[gotframe] ),
        .O(\gmiimode0.r[gotframe]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFFFFFF02000000)) 
    \gmiimode0.r[icnt][0]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .O(\gmiimode0.r[icnt][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF2FFFFFF08000000)) 
    \gmiimode0.r[icnt][1]_i_1 
       (.I0(\gmiimode0.r[byte_count][6]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .I2(\gmiimode0.r[tx_en]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .O(\gmiimode0.r[icnt][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0A02)) 
    \gmiimode0.r[ifg_cycls][0]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .I1(\gmiimode0.r[ifg_cycls][3]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/d [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .O(\gmiimode0.r[ifg_cycls][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA00A2002)) 
    \gmiimode0.r[ifg_cycls][1]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .I1(\gmiimode0.r[ifg_cycls][3]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/d [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/d [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .O(\gmiimode0.r[ifg_cycls][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAA0000A22200002)) 
    \gmiimode0.r[ifg_cycls][2]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .I1(\gmiimode0.r[ifg_cycls][3]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/d [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/d [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/d [2]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .O(\gmiimode0.r[ifg_cycls][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA00A2002)) 
    \gmiimode0.r[ifg_cycls][3]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .I1(\gmiimode0.r[ifg_cycls][3]_i_2_n_0 ),
        .I2(\gmiimode0.r[ifg_cycls][3]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/d [3]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .O(\gmiimode0.r[ifg_cycls][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4044FFFF)) 
    \gmiimode0.r[ifg_cycls][3]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in38_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/rin ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_prev_n_0_] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_act]__1 ),
        .I4(\gmiimode0.r[ifg_cycls][7]_i_2_n_0 ),
        .O(\gmiimode0.r[ifg_cycls][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \gmiimode0.r[ifg_cycls][3]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/d [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/d [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/d [0]),
        .O(\gmiimode0.r[ifg_cycls][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4E0E0A0EFFFF0000)) 
    \gmiimode0.r[ifg_cycls][4]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .I1(\gmiimode0.r[ifg_cycls][7]_i_2_n_0 ),
        .I2(\gmiimode0.r[ifg_cycls][4]_i_2_n_0 ),
        .I3(\gmiimode0.r[ifg_cycls][8]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .O(\gmiimode0.r[ifg_cycls][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55555556)) 
    \gmiimode0.r[ifg_cycls][4]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/d [4]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/d [2]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/d [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/d [0]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/d [3]),
        .O(\gmiimode0.r[ifg_cycls][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB0F5F4A00000FFFF)) 
    \gmiimode0.r[ifg_cycls][5]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .I1(\gmiimode0.r[ifg_cycls][8]_i_5_n_0 ),
        .I2(\gmiimode0.r[ifg_cycls][5]_i_2_n_0 ),
        .I3(\gmiimode0.r[ifg_cycls][7]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .O(\gmiimode0.r[ifg_cycls][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA9)) 
    \gmiimode0.r[ifg_cycls][5]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/d [5]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/d [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/d [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/d [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/d [2]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/d [4]),
        .O(\gmiimode0.r[ifg_cycls][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8888888800800A8A)) 
    \gmiimode0.r[ifg_cycls][6]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .I1(\gmiimode0.r[ifg_cycls][6]_i_2_n_0 ),
        .I2(\gmiimode0.r[ifg_cycls][7]_i_2_n_0 ),
        .I3(\gmiimode0.r[ifg_cycls][8]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .O(\gmiimode0.r[ifg_cycls][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE01)) 
    \gmiimode0.r[ifg_cycls][6]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/d [5]),
        .I1(\gmiimode0.r[ifg_cycls][8]_i_6_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/d [4]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/d [6]),
        .O(\gmiimode0.r[ifg_cycls][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0A0E4E0E0000FFFF)) 
    \gmiimode0.r[ifg_cycls][7]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .I1(\gmiimode0.r[ifg_cycls][7]_i_2_n_0 ),
        .I2(\gmiimode0.r[ifg_cycls][7]_i_3_n_0 ),
        .I3(\gmiimode0.r[ifg_cycls][8]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .O(\gmiimode0.r[ifg_cycls][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \gmiimode0.r[ifg_cycls][7]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/d [8]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/d [6]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/d [4]),
        .I3(\gmiimode0.r[ifg_cycls][8]_i_6_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/d [5]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/d [7]),
        .O(\gmiimode0.r[ifg_cycls][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55555556)) 
    \gmiimode0.r[ifg_cycls][7]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/d [7]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/d [5]),
        .I2(\gmiimode0.r[ifg_cycls][8]_i_6_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/d [4]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/d [6]),
        .O(\gmiimode0.r[ifg_cycls][7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555555544440004)) 
    \gmiimode0.r[ifg_cycls][8]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[transmitting]__0 ),
        .I3(\gmiimode0.r[ifg_cycls][8]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in38_in ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[ifg_cycls] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA00AA00A0002A002)) 
    \gmiimode0.r[ifg_cycls][8]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\gmiimode0.r[ifg_cycls][8]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/d [8]),
        .I4(\gmiimode0.r[ifg_cycls][8]_i_5_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .O(\gmiimode0.r[ifg_cycls][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \gmiimode0.r[ifg_cycls][8]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/rin ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_prev_n_0_] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_act]__1 ),
        .O(\gmiimode0.r[ifg_cycls][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \gmiimode0.r[ifg_cycls][8]_i_4 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/d [7]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/d [5]),
        .I2(\gmiimode0.r[ifg_cycls][8]_i_6_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/d [4]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/d [6]),
        .O(\gmiimode0.r[ifg_cycls][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00D0)) 
    \gmiimode0.r[ifg_cycls][8]_i_5 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_act]__1 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_prev_n_0_] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/rin ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in38_in ),
        .O(\gmiimode0.r[ifg_cycls][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \gmiimode0.r[ifg_cycls][8]_i_6 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/d [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/d [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/d [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/d [2]),
        .O(\gmiimode0.r[ifg_cycls][8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00001000)) 
    \gmiimode0.r[lentype][15]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [4]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/write_req ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[ltfound_n_0_] ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFF0000)) 
    \gmiimode0.r[ltfound]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[ltfound_n_0_] ),
        .O(\gmiimode0.r[ltfound]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFCEFE00003000)) 
    \gmiimode0.r[odd_nibble]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I3(\gmiimode0.r[odd_nibble]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[odd_nibble_n_0_] ),
        .O(\gmiimode0.r[odd_nibble]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hE0000000)) 
    \gmiimode0.r[odd_nibble]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero]__0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[en]__0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dv]__0 ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .O(\gmiimode0.r[odd_nibble]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \gmiimode0.r[random][0]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_1_in75_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in74_in ),
        .O(\gmiimode0.r[random][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0BBBBBBBBBBBBBBF)) 
    \gmiimode0.r[rcnt][0]_i_1 
       (.I0(\gmiimode0.r[rcnt][0]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[rcnt] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \gmiimode0.r[rcnt][0]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .O(\gmiimode0.r[rcnt][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99090000)) 
    \gmiimode0.r[rcnt][1]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I4(\gmiimode0.r[rcnt][2]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[rcnt] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD0D0D00D00000000)) 
    \gmiimode0.r[rcnt][2]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][0] ),
        .I5(\gmiimode0.r[rcnt][2]_i_2_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[rcnt] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFE)) 
    \gmiimode0.r[rcnt][2]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .O(\gmiimode0.r[rcnt][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h2AAAAAAB)) 
    \gmiimode0.r[rcnt][3]_i_1 
       (.I0(\etho[tx_en] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .O(\gmiimode0.r[rcnt][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h2AAAAAAB)) 
    \gmiimode0.r[rcnt][3]_i_2 
       (.I0(\gmiimode0.r[rcnt][3]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[rcnt] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFF44444444F)) 
    \gmiimode0.r[rcnt][3]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][3] ),
        .O(\gmiimode0.r[rcnt][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEFEEEF10101110)) 
    \gmiimode0.r[read]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\gmiimode0.r[read]_i_2_n_0 ),
        .I3(\gmiimode0.r[byte_count][10]_i_4__0_n_0 ),
        .I4(\gmiimode0.r[start][1]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/txo[read] ),
        .O(\gmiimode0.r[read]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h10000000F0000000)) 
    \gmiimode0.r[read]_i_2 
       (.I0(\gmiimode0.r[read]_i_3_n_0 ),
        .I1(\gmiimode0.r_reg[tx_en]_i_7_n_0 ),
        .I2(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_28_out ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\gmiimode0.r[read]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \gmiimode0.r[read]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .O(\gmiimode0.r[read]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF7FFFFFF08000000)) 
    \gmiimode0.r[restart]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I4(\gmiimode0.r[restart]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/txo[restart] ),
        .O(\gmiimode0.r[restart]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFD)) 
    \gmiimode0.r[restart]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .O(\gmiimode0.r[restart]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \gmiimode0.r[retry_cnt][0]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .O(\gmiimode0.r[retry_cnt][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \gmiimode0.r[retry_cnt][1]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[retry_cnt] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h006A)) 
    \gmiimode0.r[retry_cnt][2]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[retry_cnt] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00006AAA)) 
    \gmiimode0.r[retry_cnt][3]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[retry_cnt] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40404000)) 
    \gmiimode0.r[retry_cnt][4]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]14_out ),
        .O(\gmiimode0.r[retry_cnt][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000006AAAAAAA)) 
    \gmiimode0.r[retry_cnt][4]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[retry_cnt] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000002)) 
    \gmiimode0.r[retry_cnt][4]_i_3 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]14_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE000)) 
    \gmiimode0.r[rmii_crc_en]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I2(\etho[tx_en] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch]__0 ),
        .O(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBABB8A88)) 
    \gmiimode0.r[rxd2][0]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dv]__0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero]__0 ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .O(\gmiimode0.r[rxd2][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBABB8A88)) 
    \gmiimode0.r[rxd2][1]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dv]__0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero]__0 ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .O(\gmiimode0.r[rxd2][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFEAAAAAA)) 
    \gmiimode0.r[rxdp][3]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/v ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero]__0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[en]__0 ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dv]__0 ),
        .O(\gmiimode0.r[rxdp][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \gmiimode0.r[rxdp][3]_i_2 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .I5(\gmiimode0.r[rxdp][3]_i_3_n_0 ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/v ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h1F)) 
    \gmiimode0.r[rxdp][3]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero]__0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[en]__0 ),
        .O(\gmiimode0.r[rxdp][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h13)) 
    \gmiimode0.r[slot_count][0]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][0] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h090F)) 
    \gmiimode0.r[slot_count][1]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][1] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][0] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00A900FF)) 
    \gmiimode0.r[slot_count][2]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][2] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][0] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000AAA90000FFFF)) 
    \gmiimode0.r[slot_count][3]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][3] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][1] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][2] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h090F)) 
    \gmiimode0.r[slot_count][4]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][4] ),
        .I1(\gmiimode0.r[slot_count][4]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \gmiimode0.r[slot_count][4]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][2] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][0] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][3] ),
        .O(\gmiimode0.r[slot_count][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h090F)) 
    \gmiimode0.r[slot_count][5]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][5] ),
        .I1(\gmiimode0.r[slot_count][5]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \gmiimode0.r[slot_count][5]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][3] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][1] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][2] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][4] ),
        .O(\gmiimode0.r[slot_count][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \gmiimode0.r[slot_count][6]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .O(\gmiimode0.r[slot_count][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h090F)) 
    \gmiimode0.r[slot_count][6]_i_2 
       (.I0(\gmiimode0.r[delay_val][9]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][6] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCCCCCCCCCCCCD8)) 
    \gmiimode0.r[start][1]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[deferring_n_0_] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [0]),
        .I3(\gmiimode0.r[start][1]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .O(\gmiimode0.r[start][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \gmiimode0.r[start][1]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .O(\gmiimode0.r[start][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80FF8000)) 
    \gmiimode0.r[start]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I3(\gmiimode0.r[start]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[start]__0 ),
        .O(\gmiimode0.r[start]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000008040004)) 
    \gmiimode0.r[start]_i_2 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\gmiimode0.r[start]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F00FFFF2F000000)) 
    \gmiimode0.r[status][0]_i_1 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\gmiimode0.r[status][0]_i_2_n_0 ),
        .I4(\gmiimode0.r[status][0]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/txo[status] [0]),
        .O(\gmiimode0.r[status][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAABAFFBFAA8A0080)) 
    \gmiimode0.r[status][0]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\gmiimode0.r[status][2]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[odd_nibble_n_0_] ),
        .I3(\gmiimode0.r[status][2]_i_3_n_0 ),
        .I4(\gmiimode0.r[status][3]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/rxo[status] [0]),
        .O(\gmiimode0.r[status][0]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \gmiimode0.r[status][0]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .O(\gmiimode0.r[status][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000003B112A00)) 
    \gmiimode0.r[status][0]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\gmiimode0.r[data][31]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]9_out ),
        .I4(\gmiimode0.r[byte_count][10]_i_4__0_n_0 ),
        .I5(\gmiimode0.r[tx_en]_i_5_n_0 ),
        .O(\gmiimode0.r[status][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFF800000008)) 
    \gmiimode0.r[status][1]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\gmiimode0.r[status][1]_i_2_n_0 ),
        .I4(\gmiimode0.r[status][1]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/txo[status] [1]),
        .O(\gmiimode0.r[status][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEFE00001000)) 
    \gmiimode0.r[status][1]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/v[status] ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .I5(\m100.u0/ethc0/rxo[status] [1]),
        .O(\gmiimode0.r[status][1]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAA8AAAAAAAA)) 
    \gmiimode0.r[status][1]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .O(\gmiimode0.r[status][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFFFFFFFFF9)) 
    \gmiimode0.r[status][1]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[deferring_n_0_] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .O(\gmiimode0.r[status][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAABFFFBAAA80008)) 
    \gmiimode0.r[status][2]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I1(\gmiimode0.r[status][2]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[odd_nibble_n_0_] ),
        .I3(\gmiimode0.r[status][2]_i_3_n_0 ),
        .I4(\gmiimode0.r[status][3]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/rxo[status] [2]),
        .O(\gmiimode0.r[status][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \gmiimode0.r[status][2]_i_10 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_10_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_9_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][1] ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][0] ),
        .O(\gmiimode0.r[status][2]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \gmiimode0.r[status][2]_i_11 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_29_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_23_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_33_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_30_in72_in ),
        .O(\gmiimode0.r[status][2]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \gmiimode0.r[status][2]_i_2 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\gmiimode0.r[status][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \gmiimode0.r[status][2]_i_3 
       (.I0(\gmiimode0.r[status][2]_i_4_n_0 ),
        .I1(\gmiimode0.r[status][2]_i_5_n_0 ),
        .I2(\gmiimode0.r[status][2]_i_6_n_0 ),
        .I3(\gmiimode0.r[status][2]_i_7_n_0 ),
        .O(\gmiimode0.r[status][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \gmiimode0.r[status][2]_i_4 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_26_in64_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_27_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_24_in59_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_25_in ),
        .I4(\gmiimode0.r[status][2]_i_8_n_0 ),
        .O(\gmiimode0.r[status][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \gmiimode0.r[status][2]_i_5 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_15_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_32_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_19_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_31_in ),
        .I4(\gmiimode0.r[status][2]_i_9_n_0 ),
        .O(\gmiimode0.r[status][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    \gmiimode0.r[status][2]_i_6 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_11_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_16_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][6] ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_14_in ),
        .I4(\gmiimode0.r[status][2]_i_10_n_0 ),
        .O(\gmiimode0.r[status][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    \gmiimode0.r[status][2]_i_7 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_20_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_22_in55_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_17_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_18_in ),
        .I4(\gmiimode0.r[status][2]_i_11_n_0 ),
        .O(\gmiimode0.r[status][2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \gmiimode0.r[status][2]_i_8 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][27] ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_28_in69_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in15_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .O(\gmiimode0.r[status][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF7)) 
    \gmiimode0.r[status][2]_i_9 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in12_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in10_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_13_in ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][2] ),
        .O(\gmiimode0.r[status][2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8CAEAE8CFFAEAEFF)) 
    \gmiimode0.r[status][3]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/write_req ),
        .I1(\m100.u0/ethc0/rxo[status] [3]),
        .I2(\gmiimode0.r[status][3]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[write_ack] ),
        .I4(\m100.u0/ethc0/rxo[write] ),
        .I5(\m100.u0/ethc0/r_reg[writeok_n_0_] ),
        .O(\gmiimode0.r[status][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000002000000)) 
    \gmiimode0.r[status][3]_i_2 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I3(\gmiimode0.r[status][3]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[start]__0 ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/write_req ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \gmiimode0.r[status][3]_i_3 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .O(\gmiimode0.r[status][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \gmiimode0.r[status][3]_i_4 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .I3(\m100.u0/ethc0/rxo[byte_count] [1]),
        .O(\gmiimode0.r[status][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD55555542AAAAAA8)) 
    \gmiimode0.r[switch]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v[switch]3_out ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch]__0 ),
        .O(\gmiimode0.r[switch]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA8)) 
    \gmiimode0.r[switch]_i_2 
       (.I0(\etho[tx_en] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[switch]3_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEF00000010)) 
    \gmiimode0.r[sync_start]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .I2(\gmiimode0.r[sync_start]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .I5(\m100.u0/ethc0/rxo[start] ),
        .O(\gmiimode0.r[sync_start]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \gmiimode0.r[sync_start]_i_2 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/dv17_in ),
        .I1(\gmiimode0.r[sync_start]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp_n_0_][1] ),
        .I4(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp_n_0_][0] ),
        .I5(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp_n_0_][3] ),
        .O(\gmiimode0.r[sync_start]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF7F)) 
    \gmiimode0.r[sync_start]_i_3 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp_n_0_][2] ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .O(\gmiimode0.r[sync_start]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF33FFFFE00000002)) 
    \gmiimode0.r[transmitting]_i_1 
       (.I0(\gmiimode0.r[byte_count][10]_i_4__0_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[transmitting]__0 ),
        .O(\gmiimode0.r[transmitting]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \gmiimode0.r[tx_en]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/txrst ),
        .O(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0990909060090909)) 
    \gmiimode0.r[tx_en]_i_10 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][10] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][10] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][9] ),
        .I3(\gmiimode0.r[tx_en]_i_14_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][8] ),
        .I5(\m100.u0/ethc0/r_reg[txlength_n_0_][9] ),
        .O(\gmiimode0.r[tx_en]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \gmiimode0.r[tx_en]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][7] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [7]),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][6] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [6]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [8]),
        .I5(\m100.u0/ethc0/r_reg[txlength_n_0_][8] ),
        .O(\gmiimode0.r[tx_en]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0990000000000990)) 
    \gmiimode0.r[tx_en]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [4]),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][3] ),
        .I3(\gmiimode0.r[tx_en]_i_17_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [5]),
        .I5(\m100.u0/ethc0/r_reg[txlength_n_0_][5] ),
        .O(\gmiimode0.r[tx_en]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0041820014000082)) 
    \gmiimode0.r[tx_en]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][2] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .I5(\m100.u0/ethc0/r_reg[txlength_n_0_][1] ),
        .O(\gmiimode0.r[tx_en]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \gmiimode0.r[tx_en]_i_14 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][7] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][5] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ),
        .I4(\gmiimode0.r[byte_count][6]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][6] ),
        .O(\gmiimode0.r[tx_en]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \gmiimode0.r[tx_en]_i_15 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][6] ),
        .I1(\gmiimode0.r[byte_count][6]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][5] ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \gmiimode0.r[tx_en]_i_16 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/conv_integer [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9555)) 
    \gmiimode0.r[tx_en]_i_17 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .O(\gmiimode0.r[tx_en]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFBFBFAA808080AA)) 
    \gmiimode0.r[tx_en]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I2(\gmiimode0.r[tx_en]_i_4_n_0 ),
        .I3(\gmiimode0.r[tx_en]_i_5_n_0 ),
        .I4(\gmiimode0.r[tx_en]_i_6_n_0 ),
        .I5(\etho[tx_en] ),
        .O(\gmiimode0.r[tx_en]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD5AA80)) 
    \gmiimode0.r[tx_en]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\gmiimode0.r_reg[tx_en]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_28_out ),
        .I4(\gmiimode0.r[byte_count][10]_i_4__0_n_0 ),
        .I5(\gmiimode0.r[tx_en]_i_5_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBFF88B8BB8888B8)) 
    \gmiimode0.r[tx_en]_i_4 
       (.I0(\gmiimode0.r[tx_en]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]9_out ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]14_out ),
        .O(\gmiimode0.r[tx_en]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \gmiimode0.r[tx_en]_i_5 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .O(\gmiimode0.r[tx_en]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFEFF)) 
    \gmiimode0.r[tx_en]_i_6 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[deferring_n_0_] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [0]),
        .O(\gmiimode0.r[tx_en]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF00FFFFF10000)) 
    \gmiimode0.r[tx_en]_i_8 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_28_out ),
        .I1(\gmiimode0.r[read]_i_3_n_0 ),
        .I2(\gmiimode0.r_reg[tx_en]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I4(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .O(\gmiimode0.r[tx_en]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h28AA)) 
    \gmiimode0.r[tx_en]_i_9 
       (.I0(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[read_ack] ),
        .I2(\m100.u0/ethc0/txo[read] ),
        .I3(\m100.u0/ethc0/r_reg[txvalid_n_0_] ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]9_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \gmiimode0.r[txd][0]_i_10 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_18_in [0]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_20_in [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_19_in [0]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][28] ),
        .O(\gmiimode0.r[txd][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \gmiimode0.r[txd][0]_i_11 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_24_in59_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_28_in69_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][27] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I4(\gmiimode0.r[txd][0]_i_13_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .O(\gmiimode0.r[txd][0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \gmiimode0.r[txd][0]_i_12 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_9_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_13_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/p_17_in ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/p_22_in55_in ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .O(\gmiimode0.r[txd][0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEA2A)) 
    \gmiimode0.r[txd][0]_i_13 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in10_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][27] ),
        .O(\gmiimode0.r[txd][0]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00004700)) 
    \gmiimode0.r[txd][0]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdata_n_0_][24] ),
        .I1(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I2(\gmiimode0.r[txd][0]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I4(\gmiimode0.r[tx_en]_i_5_n_0 ),
        .I5(\gmiimode0.r[txd][2]_i_5_n_0 ),
        .O(\gmiimode0.r[txd][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFBFFFB15110501)) 
    \gmiimode0.r[txd][0]_i_3 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\gmiimode0.r[txd][0]_i_6_n_0 ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]14_out ),
        .I5(\gmiimode0.r[txd][0]_i_5_n_0 ),
        .O(\gmiimode0.r[txd][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAEEEAAAEA)) 
    \gmiimode0.r[txd][0]_i_4 
       (.I0(\gmiimode0.r[txd][0]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\gmiimode0.r[txd][0]_i_5_n_0 ),
        .I3(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I4(\gmiimode0.r_reg[txd][0]_i_8_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .O(\gmiimode0.r[txd][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFABFF0000A800)) 
    \gmiimode0.r[txd][0]_i_5 
       (.I0(\^etho[txd] [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I3(\etho[tx_en] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch]__0 ),
        .I5(\^etho[txd] [0]),
        .O(\gmiimode0.r[txd][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFFFFFFA8000000)) 
    \gmiimode0.r[txd][0]_i_6 
       (.I0(\gmiimode0.r[txd][0]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I3(\etho[tx_en] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch]__0 ),
        .I5(\gmiimode0.r[txd][0]_i_5_n_0 ),
        .O(\gmiimode0.r[txd][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3330203020202020)) 
    \gmiimode0.r[txd][0]_i_7 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\gmiimode0.r[txd][0]_i_5_n_0 ),
        .I3(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I4(\gmiimode0.r[txd][0]_i_10_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\gmiimode0.r[txd][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \gmiimode0.r[txd][0]_i_9 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][0] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_16_in [0]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_15_in [0]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][24] ),
        .O(\gmiimode0.r[txd][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \gmiimode0.r[txd][1]_i_10 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_18_in [1]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_20_in [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_19_in [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][29] ),
        .O(\gmiimode0.r[txd][1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \gmiimode0.r[txd][1]_i_11 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_8_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_12_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][10] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][14] ),
        .O(\gmiimode0.r[txd][1]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \gmiimode0.r[txd][1]_i_12 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_23_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_27_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_33_in ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I5(\gmiimode0.r[txd][1]_i_13_n_0 ),
        .O(\gmiimode0.r[txd][1]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEA2A)) 
    \gmiimode0.r[txd][1]_i_13 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_33_in ),
        .O(\gmiimode0.r[txd][1]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F000F0EECC2200)) 
    \gmiimode0.r[txd][1]_i_2 
       (.I0(\gmiimode0.r[txd][1]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\gmiimode0.r[txd][1]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I4(\gmiimode0.r[txd][1]_i_6_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .O(\gmiimode0.r[txd][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0AAAAAF20AAAAA02)) 
    \gmiimode0.r[txd][1]_i_3 
       (.I0(\gmiimode0.r[txd][1]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]14_out ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I5(\gmiimode0.r[txd][1]_i_7_n_0 ),
        .O(\gmiimode0.r[txd][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFFFFFFA8000000)) 
    \gmiimode0.r[txd][1]_i_4 
       (.I0(\gmiimode0.r[txd][1]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I3(\etho[tx_en] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch]__0 ),
        .I5(\gmiimode0.r[txd][1]_i_6_n_0 ),
        .O(\gmiimode0.r[txd][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEAEFFFFFEAEAAAA)) 
    \gmiimode0.r[txd][1]_i_5 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/r_reg[txdata_n_0_][25] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\gmiimode0.r[txd][1]_i_9_n_0 ),
        .I4(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I5(\gmiimode0.r[txd][1]_i_6_n_0 ),
        .O(\gmiimode0.r[txd][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFABFF0000A800)) 
    \gmiimode0.r[txd][1]_i_6 
       (.I0(\^etho[txd] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I3(\etho[tx_en] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch]__0 ),
        .I5(\^etho[txd] [1]),
        .O(\gmiimode0.r[txd][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFFFFFFA8000000)) 
    \gmiimode0.r[txd][1]_i_7 
       (.I0(\gmiimode0.r[txd][1]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I3(\etho[tx_en] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch]__0 ),
        .I5(\gmiimode0.r[txd][1]_i_6_n_0 ),
        .O(\gmiimode0.r[txd][1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \gmiimode0.r[txd][1]_i_8 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][1] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_16_in [1]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_15_in [1]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][25] ),
        .O(\gmiimode0.r[txd][1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \gmiimode0.r[txd][1]_i_9 
       (.I0(\gmiimode0.r[txd][1]_i_11_n_0 ),
        .I1(\gmiimode0.r[txd][1]_i_12_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .O(\gmiimode0.r[txd][1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAEAEAFFEAEAEA00)) 
    \gmiimode0.r[txd][2]_i_1 
       (.I0(\gmiimode0.r[txd][2]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\gmiimode0.r[txd][2]_i_3_n_0 ),
        .I3(\gmiimode0.r[txd][2]_i_4_n_0 ),
        .I4(\gmiimode0.r[txd][2]_i_5_n_0 ),
        .I5(\gmiimode0.r[txd][2]_i_6_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/rin[txd_msb] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFFFFFFA8000000)) 
    \gmiimode0.r[txd][2]_i_10 
       (.I0(\gmiimode0.r[txd][2]_i_11_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I3(\etho[tx_en] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch]__0 ),
        .I5(\^etho[txd] [2]),
        .O(\gmiimode0.r[txd][2]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \gmiimode0.r[txd][2]_i_11 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][2] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_16_in [2]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_15_in [2]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][26] ),
        .O(\gmiimode0.r[txd][2]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3330203020202020)) 
    \gmiimode0.r[txd][2]_i_2 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\^etho[txd] [2]),
        .I3(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I4(\gmiimode0.r[txd][2]_i_7_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .O(\gmiimode0.r[txd][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000222EE2EE)) 
    \gmiimode0.r[txd][2]_i_3 
       (.I0(\^etho[txd] [2]),
        .I1(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .I3(\gmiimode0.r[txd][2]_i_8_n_0 ),
        .I4(\gmiimode0.r[txd][2]_i_9_n_0 ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .O(\gmiimode0.r[txd][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000001010100010)) 
    \gmiimode0.r[txd][2]_i_4 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\^etho[txd] [2]),
        .I4(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txdata_n_0_][26] ),
        .O(\gmiimode0.r[txd][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9600)) 
    \gmiimode0.r[txd][2]_i_5 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .O(\gmiimode0.r[txd][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFB1511FFFB0501)) 
    \gmiimode0.r[txd][2]_i_6 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .I3(\gmiimode0.r[txd][2]_i_10_n_0 ),
        .I4(\^etho[txd] [2]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]14_out ),
        .O(\gmiimode0.r[txd][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \gmiimode0.r[txd][2]_i_7 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_18_in [2]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_20_in [2]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_19_in [2]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][30] ),
        .O(\gmiimode0.r[txd][2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0C0C0AFA0CFCF)) 
    \gmiimode0.r[txd][2]_i_8 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_32_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_26_in64_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_30_in72_in ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I5(\gmiimode0.r[crc][29]_i_2_n_0 ),
        .O(\gmiimode0.r[txd][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \gmiimode0.r[txd][2]_i_9 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][1] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_11_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][9] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][13] ),
        .O(\gmiimode0.r[txd][2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \gmiimode0.r[txd][3]_i_10 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][0] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_10_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_14_in ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][12] ),
        .O(\gmiimode0.r[txd][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0C0C0AFA0CFCF)) 
    \gmiimode0.r[txd][3]_i_11 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_31_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_25_in ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][24] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I5(\gmiimode0.r[crc][28]_i_2_n_0 ),
        .O(\gmiimode0.r[txd][3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F000F0EECC2200)) 
    \gmiimode0.r[txd][3]_i_2 
       (.I0(\gmiimode0.r[txd][3]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I2(\gmiimode0.r[txd][3]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I4(\^etho[txd] [3]),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .O(\gmiimode0.r[txd][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0AAAAAFE0AAAAA0E)) 
    \gmiimode0.r[txd][3]_i_3 
       (.I0(\^etho[txd] [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/v[tx_en]14_out ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I5(\gmiimode0.r[txd][3]_i_6_n_0 ),
        .O(\gmiimode0.r[txd][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFFFFFFA8000000)) 
    \gmiimode0.r[txd][3]_i_4 
       (.I0(\gmiimode0.r[txd][3]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I3(\etho[tx_en] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch]__0 ),
        .I5(\^etho[txd] [3]),
        .O(\gmiimode0.r[txd][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEAEFFFFFEAEAAAA)) 
    \gmiimode0.r[txd][3]_i_5 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .I1(\m100.u0/ethc0/r_reg[txdata_n_0_][27] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .I3(\gmiimode0.r[txd][3]_i_8_n_0 ),
        .I4(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .I5(\^etho[txd] [3]),
        .O(\gmiimode0.r[txd][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFFFFFFA8000000)) 
    \gmiimode0.r[txd][3]_i_6 
       (.I0(\gmiimode0.r[txd][3]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I3(\etho[tx_en] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch]__0 ),
        .I5(\^etho[txd] [3]),
        .O(\gmiimode0.r[txd][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \gmiimode0.r[txd][3]_i_7 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][3] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_16_in [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_15_in [3]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][27] ),
        .O(\gmiimode0.r[txd][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \gmiimode0.r[txd][3]_i_8 
       (.I0(\gmiimode0.r[txd][3]_i_10_n_0 ),
        .I1(\gmiimode0.r[txd][3]_i_11_n_0 ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .O(\gmiimode0.r[txd][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \gmiimode0.r[txd][3]_i_9 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/p_18_in [3]),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/p_20_in [3]),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/p_19_in [3]),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][31] ),
        .O(\gmiimode0.r[txd][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF072)) 
    \gmiimode0.r[write]_i_1 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/write_req ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[write_ack] ),
        .I2(\m100.u0/ethc0/rxo[write] ),
        .I3(\m100.u0/ethc0/rxo[status] [3]),
        .O(\gmiimode0.r[write]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000CAAAAAAAA)) 
    \gmiimode0.r[zero]_i_1 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][3] ),
        .I5(\m100.u0/ethc0/tx_rmii1.tx0/v[zero]7_out ),
        .O(\gmiimode0.r[zero]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \gmiimode0.r[zero]_i_1__0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][3] ),
        .O(\gmiimode0.r[zero]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \gmiimode0.r[zero]_i_2 
       (.I0(\etho[tx_en] ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/v[zero]7_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \gmiimode0.r_reg[byte_count][10]_i_3 
       (.CI(\gmiimode0.r_reg[byte_count][7]_i_2_n_0 ),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O(\gmiimode0.r_reg ),
        .S({etho,\m100.u0/ethc0/rxo[byte_count] [10:8]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \gmiimode0.r_reg[byte_count][3]_i_2 
       (.CI(etho),
        .CO({\gmiimode0.r_reg[byte_count][3]_i_2_n_0 ,\gmiimode0.r_reg[byte_count][3]_i_2_n_1 ,\gmiimode0.r_reg[byte_count][3]_i_2_n_2 ,\gmiimode0.r_reg[byte_count][3]_i_2_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,\m100.u0/ethc0/rxo[byte_count] [0]}),
        .O({\gmiimode0.r_reg[byte_count][3]_i_2_n_4 ,\m100.u0/ethc0/rx_rmii1.rx0/p_1_in6_in ,\gmiimode0.r_reg[byte_count][3]_i_2_n_6 ,\gmiimode0.r_reg[byte_count][3]_i_2_n_7 }),
        .S({\m100.u0/ethc0/rxo[byte_count] [3:1],\gmiimode0.r[byte_count][3]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \gmiimode0.r_reg[byte_count][7]_i_2 
       (.CI(\gmiimode0.r_reg[byte_count][3]_i_2_n_0 ),
        .CO({\gmiimode0.r_reg[byte_count][7]_i_2_n_0 ,\gmiimode0.r_reg[byte_count][7]_i_2_n_1 ,\gmiimode0.r_reg[byte_count][7]_i_2_n_2 ,\gmiimode0.r_reg[byte_count][7]_i_2_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\gmiimode0.r_reg[byte_count][7]_i_2_n_4 ,\gmiimode0.r_reg[byte_count][7]_i_2_n_5 ,\gmiimode0.r_reg[byte_count][7]_i_2_n_6 ,\gmiimode0.r_reg[byte_count][7]_i_2_n_7 }),
        .S(\m100.u0/ethc0/rxo[byte_count] [7:4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \gmiimode0.r_reg[tx_en]_i_7 
       (.CI(etho),
        .CO({\gmiimode0.r_reg[tx_en]_i_7_n_0 ,\gmiimode0.r_reg[tx_en]_i_7_n_1 ,\gmiimode0.r_reg[tx_en]_i_7_n_2 ,\gmiimode0.r_reg[tx_en]_i_7_n_3 }),
        .CYINIT(apbo),
        .DI({etho,etho,etho,etho}),
        .S({\gmiimode0.r[tx_en]_i_10_n_0 ,\gmiimode0.r[tx_en]_i_11_n_0 ,\gmiimode0.r[tx_en]_i_12_n_0 ,\gmiimode0.r[tx_en]_i_13_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \gmiimode0.r_reg[txd][0]_i_1 
       (.I0(\gmiimode0.r[txd][0]_i_3_n_0 ),
        .I1(\gmiimode0.r[txd][0]_i_4_n_0 ),
        .O(\gmiimode0.r_reg[txd][0]_i_1_n_0 ),
        .S(\gmiimode0.r[txd][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \gmiimode0.r_reg[txd][0]_i_8 
       (.I0(\gmiimode0.r[txd][0]_i_11_n_0 ),
        .I1(\gmiimode0.r[txd][0]_i_12_n_0 ),
        .O(\gmiimode0.r_reg[txd][0]_i_8_n_0 ),
        .S(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \gmiimode0.r_reg[txd][1]_i_1 
       (.I0(\gmiimode0.r[txd][1]_i_2_n_0 ),
        .I1(\gmiimode0.r[txd][1]_i_3_n_0 ),
        .O(\gmiimode0.r_reg[txd][1]_i_1_n_0 ),
        .S(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \gmiimode0.r_reg[txd][3]_i_1 
       (.I0(\gmiimode0.r[txd][3]_i_2_n_0 ),
        .I1(\gmiimode0.r[txd][3]_i_3_n_0 ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/rin[txd_msb] [1]),
        .S(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* PWROPT_WRITE_MODE_CHANGE_A = "WRITE_FIRST:NO_CHANGE_1" *) 
  (* XILINX_LEGACY_PRIM = "RAMB16_S36_S36" *) 
  (* XILINX_TRANSFORM_PINMAP = "ADDRA[0]:ADDRARDADDR[0],ADDRARDADDR[10] ADDRA[1]:ADDRARDADDR[1],ADDRARDADDR[11] ADDRA[2]:ADDRARDADDR[2],ADDRARDADDR[12] ADDRA[3]:ADDRARDADDR[3],ADDRARDADDR[13] ADDRA[4]:ADDRARDADDR[4],ADDRARDADDR[9] ADDRB[0]:ADDRBWRADDR[0],ADDRBWRADDR[10] ADDRB[1]:ADDRBWRADDR[1],ADDRBWRADDR[11] ADDRB[2]:ADDRBWRADDR[2],ADDRBWRADDR[12] ADDRB[3]:ADDRBWRADDR[3],ADDRBWRADDR[13] ADDRB[4]:ADDRBWRADDR[4],ADDRBWRADDR[9] WEA:WEA[3],WEA[2],WEA[1],WEA[0] WEB:WEBWE[3],WEBWE[2],WEBWE[1],WEBWE[0] ADDRA[14]:ADDRARDADDR[14] ADDRA[5]:ADDRARDADDR[5] ADDRA[6]:ADDRARDADDR[6] ADDRA[7]:ADDRARDADDR[7] ADDRA[8]:ADDRARDADDR[8] ADDRB[14]:ADDRBWRADDR[14] ADDRB[5]:ADDRBWRADDR[5] ADDRB[6]:ADDRBWRADDR[6] ADDRB[7]:ADDRBWRADDR[7] ADDRB[8]:ADDRBWRADDR[8] CLKA:CLKARDCLK CLKB:CLKBWRCLK DIA[0]:DIADI[0] DIA[10]:DIADI[10] DIA[11]:DIADI[11] DIA[12]:DIADI[12] DIA[13]:DIADI[13] DIA[14]:DIADI[14] DIA[15]:DIADI[15] DIA[16]:DIADI[16] DIA[17]:DIADI[17] DIA[18]:DIADI[18] DIA[19]:DIADI[19] DIA[1]:DIADI[1] DIA[20]:DIADI[20] DIA[21]:DIADI[21] DIA[22]:DIADI[22] DIA[23]:DIADI[23] DIA[24]:DIADI[24] DIA[25]:DIADI[25] DIA[26]:DIADI[26] DIA[27]:DIADI[27] DIA[28]:DIADI[28] DIA[29]:DIADI[29] DIA[2]:DIADI[2] DIA[30]:DIADI[30] DIA[31]:DIADI[31] DIA[3]:DIADI[3] DIA[4]:DIADI[4] DIA[5]:DIADI[5] DIA[6]:DIADI[6] DIA[7]:DIADI[7] DIA[8]:DIADI[8] DIA[9]:DIADI[9] DIB[0]:DIBDI[0] DIB[10]:DIBDI[10] DIB[11]:DIBDI[11] DIB[12]:DIBDI[12] DIB[13]:DIBDI[13] DIB[14]:DIBDI[14] DIB[15]:DIBDI[15] DIB[16]:DIBDI[16] DIB[17]:DIBDI[17] DIB[18]:DIBDI[18] DIB[19]:DIBDI[19] DIB[1]:DIBDI[1] DIB[20]:DIBDI[20] DIB[21]:DIBDI[21] DIB[22]:DIBDI[22] DIB[23]:DIBDI[23] DIB[24]:DIBDI[24] DIB[25]:DIBDI[25] DIB[26]:DIBDI[26] DIB[27]:DIBDI[27] DIB[28]:DIBDI[28] DIB[29]:DIBDI[29] DIB[2]:DIBDI[2] DIB[30]:DIBDI[30] DIB[31]:DIBDI[31] DIB[3]:DIBDI[3] DIB[4]:DIBDI[4] DIB[5]:DIBDI[5] DIB[6]:DIBDI[6] DIB[7]:DIBDI[7] DIB[8]:DIBDI[8] DIB[9]:DIBDI[9] DIPA[0]:DIPADIP[0] DIPA[1]:DIPADIP[1] DIPA[2]:DIPADIP[2] DIPA[3]:DIPADIP[3] DIPB[0]:DIPBDIP[0] DIPB[1]:DIPBDIP[1] DIPB[2]:DIPBDIP[2] DIPB[3]:DIPBDIP[3] DOA[0]:DOADO[0] DOA[10]:DOADO[10] DOA[11]:DOADO[11] DOA[12]:DOADO[12] DOA[13]:DOADO[13] DOA[14]:DOADO[14] DOA[15]:DOADO[15] DOA[16]:DOADO[16] DOA[17]:DOADO[17] DOA[18]:DOADO[18] DOA[19]:DOADO[19] DOA[1]:DOADO[1] DOA[20]:DOADO[20] DOA[21]:DOADO[21] DOA[22]:DOADO[22] DOA[23]:DOADO[23] DOA[24]:DOADO[24] DOA[25]:DOADO[25] DOA[26]:DOADO[26] DOA[27]:DOADO[27] DOA[28]:DOADO[28] DOA[29]:DOADO[29] DOA[2]:DOADO[2] DOA[30]:DOADO[30] DOA[31]:DOADO[31] DOA[3]:DOADO[3] DOA[4]:DOADO[4] DOA[5]:DOADO[5] DOA[6]:DOADO[6] DOA[7]:DOADO[7] DOA[8]:DOADO[8] DOA[9]:DOADO[9] DOB[0]:DOBDO[0] DOB[10]:DOBDO[10] DOB[11]:DOBDO[11] DOB[12]:DOBDO[12] DOB[13]:DOBDO[13] DOB[14]:DOBDO[14] DOB[15]:DOBDO[15] DOB[16]:DOBDO[16] DOB[17]:DOBDO[17] DOB[18]:DOBDO[18] DOB[19]:DOBDO[19] DOB[1]:DOBDO[1] DOB[20]:DOBDO[20] DOB[21]:DOBDO[21] DOB[22]:DOBDO[22] DOB[23]:DOBDO[23] DOB[24]:DOBDO[24] DOB[25]:DOBDO[25] DOB[26]:DOBDO[26] DOB[27]:DOBDO[27] DOB[28]:DOBDO[28] DOB[29]:DOBDO[29] DOB[2]:DOBDO[2] DOB[30]:DOBDO[30] DOB[31]:DOBDO[31] DOB[3]:DOBDO[3] DOB[4]:DOBDO[4] DOB[5]:DOBDO[5] DOB[6]:DOBDO[6] DOB[7]:DOBDO[7] DOB[8]:DOBDO[8] DOB[9]:DOBDO[9] DOPA[0]:DOPADOP[0] DOPA[1]:DOPADOP[1] DOPA[2]:DOPADOP[2] DOPA[3]:DOPADOP[3] DOPB[0]:DOPBDOP[0] DOPB[1]:DOPBDOP[1] DOPB[2]:DOPBDOP[2] DOPB[3]:DOPBDOP[3] ENA:ENARDEN ENB:ENBWREN REGCEA:REGCEAREGCE SSRA:RSTRAMARSTRAM SSRB:RSTRAMB" *) 
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
    .READ_WIDTH_A(36),
    .READ_WIDTH_B(36),
    .RSTREG_PRIORITY_A("REGCE"),
    .RSTREG_PRIORITY_B("REGCE"),
    .SIM_COLLISION_CHECK("GENERATE_X_ONLY"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("NO_CHANGE"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(36),
    .WRITE_WIDTH_B(36)) 
    \m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0 
       (.ADDRARDADDR({VCC_2,GND_2,\m100.u0/ewaddressm ,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .ADDRBWRADDR({VCC_2,GND_2,\m100.u0/eraddress ,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,\m100.u0/datain [31:16]}),
        .DIBDI({etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho}),
        .DIPADIP({etho,etho,etho,etho}),
        .DIPBDIP({etho,etho,etho,etho}),
        .DOBDO({\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_53 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_54 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_55 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_56 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_57 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_58 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_59 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_60 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_61 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_62 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_63 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_64 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_65 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_66 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_67 ,\m100.u0/edclramnft.r0/xc2v.x0/a6.x0/a9.x[0].r0_n_68 ,\m100.u0/erdata [31:16]}),
        .ENARDEN(\m100.u0/ewritem ),
        .ENBWREN(\m100.u0/erenable ),
        .REGCEAREGCE(GND_2),
        .REGCEB(GND_2),
        .RSTRAMARSTRAM(etho),
        .RSTRAMB(etho),
        .RSTREGARSTREG(GND_2),
        .RSTREGB(GND_2),
        .WEA({\m100.u0/ewritem ,\m100.u0/ewritem ,\m100.u0/ewritem ,\m100.u0/ewritem }),
        .WEBWE({GND_2,GND_2,GND_2,GND_2,etho,etho,etho,etho}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* PWROPT_WRITE_MODE_CHANGE_A = "WRITE_FIRST:NO_CHANGE_1" *) 
  (* XILINX_LEGACY_PRIM = "RAMB16_S36_S36" *) 
  (* XILINX_TRANSFORM_PINMAP = "ADDRA[0]:ADDRARDADDR[0],ADDRARDADDR[10] ADDRA[1]:ADDRARDADDR[1],ADDRARDADDR[11] ADDRA[2]:ADDRARDADDR[2],ADDRARDADDR[12] ADDRA[3]:ADDRARDADDR[3],ADDRARDADDR[13] ADDRA[4]:ADDRARDADDR[4],ADDRARDADDR[9] ADDRB[0]:ADDRBWRADDR[0],ADDRBWRADDR[10] ADDRB[1]:ADDRBWRADDR[1],ADDRBWRADDR[11] ADDRB[2]:ADDRBWRADDR[2],ADDRBWRADDR[12] ADDRB[3]:ADDRBWRADDR[3],ADDRBWRADDR[13] ADDRB[4]:ADDRBWRADDR[4],ADDRBWRADDR[9] WEA:WEA[3],WEA[2],WEA[1],WEA[0] WEB:WEBWE[3],WEBWE[2],WEBWE[1],WEBWE[0] ADDRA[14]:ADDRARDADDR[14] ADDRA[5]:ADDRARDADDR[5] ADDRA[6]:ADDRARDADDR[6] ADDRA[7]:ADDRARDADDR[7] ADDRA[8]:ADDRARDADDR[8] ADDRB[14]:ADDRBWRADDR[14] ADDRB[5]:ADDRBWRADDR[5] ADDRB[6]:ADDRBWRADDR[6] ADDRB[7]:ADDRBWRADDR[7] ADDRB[8]:ADDRBWRADDR[8] CLKA:CLKARDCLK CLKB:CLKBWRCLK DIA[0]:DIADI[0] DIA[10]:DIADI[10] DIA[11]:DIADI[11] DIA[12]:DIADI[12] DIA[13]:DIADI[13] DIA[14]:DIADI[14] DIA[15]:DIADI[15] DIA[16]:DIADI[16] DIA[17]:DIADI[17] DIA[18]:DIADI[18] DIA[19]:DIADI[19] DIA[1]:DIADI[1] DIA[20]:DIADI[20] DIA[21]:DIADI[21] DIA[22]:DIADI[22] DIA[23]:DIADI[23] DIA[24]:DIADI[24] DIA[25]:DIADI[25] DIA[26]:DIADI[26] DIA[27]:DIADI[27] DIA[28]:DIADI[28] DIA[29]:DIADI[29] DIA[2]:DIADI[2] DIA[30]:DIADI[30] DIA[31]:DIADI[31] DIA[3]:DIADI[3] DIA[4]:DIADI[4] DIA[5]:DIADI[5] DIA[6]:DIADI[6] DIA[7]:DIADI[7] DIA[8]:DIADI[8] DIA[9]:DIADI[9] DIB[0]:DIBDI[0] DIB[10]:DIBDI[10] DIB[11]:DIBDI[11] DIB[12]:DIBDI[12] DIB[13]:DIBDI[13] DIB[14]:DIBDI[14] DIB[15]:DIBDI[15] DIB[16]:DIBDI[16] DIB[17]:DIBDI[17] DIB[18]:DIBDI[18] DIB[19]:DIBDI[19] DIB[1]:DIBDI[1] DIB[20]:DIBDI[20] DIB[21]:DIBDI[21] DIB[22]:DIBDI[22] DIB[23]:DIBDI[23] DIB[24]:DIBDI[24] DIB[25]:DIBDI[25] DIB[26]:DIBDI[26] DIB[27]:DIBDI[27] DIB[28]:DIBDI[28] DIB[29]:DIBDI[29] DIB[2]:DIBDI[2] DIB[30]:DIBDI[30] DIB[31]:DIBDI[31] DIB[3]:DIBDI[3] DIB[4]:DIBDI[4] DIB[5]:DIBDI[5] DIB[6]:DIBDI[6] DIB[7]:DIBDI[7] DIB[8]:DIBDI[8] DIB[9]:DIBDI[9] DIPA[0]:DIPADIP[0] DIPA[1]:DIPADIP[1] DIPA[2]:DIPADIP[2] DIPA[3]:DIPADIP[3] DIPB[0]:DIPBDIP[0] DIPB[1]:DIPBDIP[1] DIPB[2]:DIPBDIP[2] DIPB[3]:DIPBDIP[3] DOA[0]:DOADO[0] DOA[10]:DOADO[10] DOA[11]:DOADO[11] DOA[12]:DOADO[12] DOA[13]:DOADO[13] DOA[14]:DOADO[14] DOA[15]:DOADO[15] DOA[16]:DOADO[16] DOA[17]:DOADO[17] DOA[18]:DOADO[18] DOA[19]:DOADO[19] DOA[1]:DOADO[1] DOA[20]:DOADO[20] DOA[21]:DOADO[21] DOA[22]:DOADO[22] DOA[23]:DOADO[23] DOA[24]:DOADO[24] DOA[25]:DOADO[25] DOA[26]:DOADO[26] DOA[27]:DOADO[27] DOA[28]:DOADO[28] DOA[29]:DOADO[29] DOA[2]:DOADO[2] DOA[30]:DOADO[30] DOA[31]:DOADO[31] DOA[3]:DOADO[3] DOA[4]:DOADO[4] DOA[5]:DOADO[5] DOA[6]:DOADO[6] DOA[7]:DOADO[7] DOA[8]:DOADO[8] DOA[9]:DOADO[9] DOB[0]:DOBDO[0] DOB[10]:DOBDO[10] DOB[11]:DOBDO[11] DOB[12]:DOBDO[12] DOB[13]:DOBDO[13] DOB[14]:DOBDO[14] DOB[15]:DOBDO[15] DOB[16]:DOBDO[16] DOB[17]:DOBDO[17] DOB[18]:DOBDO[18] DOB[19]:DOBDO[19] DOB[1]:DOBDO[1] DOB[20]:DOBDO[20] DOB[21]:DOBDO[21] DOB[22]:DOBDO[22] DOB[23]:DOBDO[23] DOB[24]:DOBDO[24] DOB[25]:DOBDO[25] DOB[26]:DOBDO[26] DOB[27]:DOBDO[27] DOB[28]:DOBDO[28] DOB[29]:DOBDO[29] DOB[2]:DOBDO[2] DOB[30]:DOBDO[30] DOB[31]:DOBDO[31] DOB[3]:DOBDO[3] DOB[4]:DOBDO[4] DOB[5]:DOBDO[5] DOB[6]:DOBDO[6] DOB[7]:DOBDO[7] DOB[8]:DOBDO[8] DOB[9]:DOBDO[9] DOPA[0]:DOPADOP[0] DOPA[1]:DOPADOP[1] DOPA[2]:DOPADOP[2] DOPA[3]:DOPADOP[3] DOPB[0]:DOPBDOP[0] DOPB[1]:DOPBDOP[1] DOPB[2]:DOPBDOP[2] DOPB[3]:DOPBDOP[3] ENA:ENARDEN ENB:ENBWREN REGCEA:REGCEAREGCE SSRA:RSTRAMARSTRAM SSRB:RSTRAMB" *) 
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
    .READ_WIDTH_A(36),
    .READ_WIDTH_B(36),
    .RSTREG_PRIORITY_A("REGCE"),
    .RSTREG_PRIORITY_B("REGCE"),
    .SIM_COLLISION_CHECK("GENERATE_X_ONLY"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("NO_CHANGE"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(36),
    .WRITE_WIDTH_B(36)) 
    \m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0 
       (.ADDRARDADDR({VCC_2,GND_2,\m100.u0/ewaddressm [8:7],\m100.u0/ewaddressl ,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .ADDRBWRADDR({VCC_2,GND_2,\m100.u0/eraddress ,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,\m100.u0/datain [15:0]}),
        .DIBDI({etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho}),
        .DIPADIP({etho,etho,etho,etho}),
        .DIPBDIP({etho,etho,etho,etho}),
        .DOBDO({\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_53 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_54 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_55 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_56 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_57 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_58 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_59 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_60 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_61 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_62 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_63 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_64 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_65 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_66 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_67 ,\m100.u0/edclramnft.r1/xc2v.x0/a6.x0/a9.x[0].r0_n_68 ,\m100.u0/erdata [15:0]}),
        .ENARDEN(\m100.u0/ewritel ),
        .ENBWREN(\m100.u0/erenable ),
        .REGCEAREGCE(GND_2),
        .REGCEB(GND_2),
        .RSTRAMARSTRAM(etho),
        .RSTRAMB(etho),
        .RSTREGARSTREG(GND_2),
        .RSTREGB(GND_2),
        .WEA({\m100.u0/ewritel ,\m100.u0/ewritel ,\m100.u0/ewritel ,\m100.u0/ewritel }),
        .WEBWE({GND_2,GND_2,GND_2,GND_2,etho,etho,etho,etho}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[edclrstate][0] 
       (.C(clk),
        .CE(\FSM_sequential_r[edclrstate][3]_i_1_n_0 ),
        .D(FSM_sequential_r),
        .Q(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[edclrstate][1] 
       (.C(clk),
        .CE(\FSM_sequential_r[edclrstate][3]_i_1_n_0 ),
        .D(\FSM_sequential_r[edclrstate][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[edclrstate][2] 
       (.C(clk),
        .CE(\FSM_sequential_r[edclrstate][3]_i_1_n_0 ),
        .D(\FSM_sequential_r[edclrstate][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[edclrstate][3] 
       (.C(clk),
        .CE(\FSM_sequential_r[edclrstate][3]_i_1_n_0 ),
        .D(\FSM_sequential_r[edclrstate][3]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[mdio_state][0] 
       (.C(clk),
        .CE(\FSM_sequential_r_reg[mdio_state][3]_i_1_n_0 ),
        .D(\FSM_sequential_r[mdio_state][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[mdio_state][1] 
       (.C(clk),
        .CE(\FSM_sequential_r_reg[mdio_state][3]_i_1_n_0 ),
        .D(\FSM_sequential_r[mdio_state][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[mdio_state][2] 
       (.C(clk),
        .CE(\FSM_sequential_r_reg[mdio_state][3]_i_1_n_0 ),
        .D(\FSM_sequential_r[mdio_state][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[mdio_state][3] 
       (.C(clk),
        .CE(\FSM_sequential_r_reg[mdio_state][3]_i_1_n_0 ),
        .D(\FSM_sequential_r[mdio_state][3]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[regaddr][0] 
       (.C(clk),
        .CE(apbo),
        .D(\FSM_sequential_r[regaddr][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[regaddr][1] 
       (.C(clk),
        .CE(apbo),
        .D(\FSM_sequential_r[regaddr][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[regaddr][2] 
       (.C(clk),
        .CE(apbo),
        .D(\FSM_sequential_r[regaddr][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[rxdstate][0] 
       (.C(clk),
        .CE(apbo),
        .D(\FSM_sequential_r[rxdstate][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[rxdstate][1] 
       (.C(clk),
        .CE(apbo),
        .D(\FSM_sequential_r[rxdstate][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/v[rmsto][write] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/FSM_sequential_r_reg[rxdstate][2] 
       (.C(clk),
        .CE(apbo),
        .D(\FSM_sequential_r[rxdstate][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/ahb0/r_reg[ba] 
       (.C(clk),
        .CE(apbo),
        .D(\r[ba]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/ahb0/r_reg ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/ahb0/r_reg[bb] 
       (.C(clk),
        .CE(apbo),
        .D(\r[bb]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/ahb0/r_reg[bb]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/ahb0/r_reg[bg] 
       (.C(clk),
        .CE(apbo),
        .D(\r[bg]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/ahb0/r_reg[bg]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/ahb0/r_reg[bo] 
       (.C(clk),
        .CE(apbo),
        .D(\r[bo]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/ahb0/r_reg[error] 
       (.C(clk),
        .CE(apbo),
        .D(\r[error]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/ahb0/r_reg[error]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/ahb0/r_reg[retry] 
       (.C(clk),
        .CE(apbo),
        .D(\r[retry]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[abufs][0] 
       (.C(clk),
        .CE(apbo),
        .D(r),
        .Q(\m100.u0/ethc0/r_reg ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[abufs][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[abufs][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[abufs][2] 
       (.C(clk),
        .CE(apbo),
        .D(\r[abufs][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[abufs_n_0_][2] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[addrdone] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r ),
        .Q(\m100.u0/ethc0/r_reg[addrdone]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[addrok] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[addrok]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[addrok_n_0_] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[applength][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\r[applength][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[applength]__0 [0]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[applength][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\r[applength][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[applength]__0 [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[applength][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\r[applength][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[applength]__0 [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[applength][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\r[applength][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[applength]__0 [3]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[applength][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\r[applength][4]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[applength]__0 [4]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[applength][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\r[applength][5]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[applength]__0 [5]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[applength][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\r[applength][6]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[applength]__0 [6]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[applength][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\r[applength][7]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[applength]__0 [7]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[applength][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\r[applength][8]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[applength]__0 [8]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[applength][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\r[applength][9]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[applength]__0 [9]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[bcast] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[bcast]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[bcast_n_0_] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[capbil][1] 
       (.C(clk),
        .CE(\r[capbil][4]_i_1_n_0 ),
        .D(\r[capbil][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[capbil_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[capbil][2] 
       (.C(clk),
        .CE(\r[capbil][4]_i_1_n_0 ),
        .D(\r[capbil][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[capbil_n_0_][2] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[capbil][3] 
       (.C(clk),
        .CE(\r[capbil][4]_i_1_n_0 ),
        .D(\r[capbil][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/p_116_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[capbil][4] 
       (.C(clk),
        .CE(\r[capbil][4]_i_1_n_0 ),
        .D(\r[capbil][4]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/p_0_in1_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[check] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/v[check] ),
        .Q(\m100.u0/ethc0/r_reg[check]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][0] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [0]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][10] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][10] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [10]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][11] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][11] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [11]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][12] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][12] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [12]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][13] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][13] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [13]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][14] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][14] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [14]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][15] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][15] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [15]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][16] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][16] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [16]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][17] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][17] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [17]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][18] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][18] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [18]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][19] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][19] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [19]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][1] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [1]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][20] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][20] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [20]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][21] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][21] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [21]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][22] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][22] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [22]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][23] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][23] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [23]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][24] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][24] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [24]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][25] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][25] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [25]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][26] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][26] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [26]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][27] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][27] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [27]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][28] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][28] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [28]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][29] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][29] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [29]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][2] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [2]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][30] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][30] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [30]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][31] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][31] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [31]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][3] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [3]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][4] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [4]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][5] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [5]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][6] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [6]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][7] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [7]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][8] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [8]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[checkdata][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[check] ),
        .D(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][9] ),
        .Q(\m100.u0/ethc0/r_reg[checkdata]__0 [9]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[cnt][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[cnt] ),
        .D(\r[cnt][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[cnt][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[cnt] ),
        .D(\r[cnt][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[cnt][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[cnt] ),
        .D(\r[cnt][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[cnt][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[cnt] ),
        .D(\r[cnt][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[cnt][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[cnt] ),
        .D(\r[cnt][4]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ctrl][edcldis] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[ctrl][edcldis]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/p_6_in [14]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ctrl][full_duplex] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[ctrl][full_duplex]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/p_6_in [4]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ctrl][prom] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[ctrl][txen] ),
        .D(\apbi[pwdata] [5]),
        .Q(\m100.u0/ethc0/p_6_in [5]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ctrl][reset] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[ctrl][txen] ),
        .D(\apbi[pwdata] [6]),
        .Q(\m100.u0/ethc0/p_6_in [6]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ctrl][rx_irqen] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[ctrl][txen] ),
        .D(\apbi[pwdata] [3]),
        .Q(\m100.u0/ethc0/p_6_in [3]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ctrl][rxen] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[ctrl][rxen]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/p_6_in [1]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ctrl][speed] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[ctrl][speed]_i_2_n_0 ),
        .Q(\etho[speed] ),
        .S(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ctrl][tx_irqen] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[ctrl][txen] ),
        .D(\apbi[pwdata] [2]),
        .Q(\m100.u0/ethc0/p_6_in [2]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ctrl][txen] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[ctrl][txen]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/p_6_in [0]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ctrlpkt] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[ctrlpkt]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[ctrlpkt]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[disableduplex] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[disableduplex]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/p_6_in [12]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[duplexstate][0] 
       (.C(clk),
        .CE(apbo),
        .D(\r[duplexstate][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[duplexstate][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[duplexstate][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[duplexstate][2] 
       (.C(clk),
        .CE(apbo),
        .D(\r[duplexstate][2]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ecnt][0] 
       (.C(clk),
        .CE(\r[ecnt][3]_i_1_n_0 ),
        .D(\r[ecnt][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ecnt][1] 
       (.C(clk),
        .CE(\r[ecnt][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ecnt] [1]),
        .Q(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ecnt][2] 
       (.C(clk),
        .CE(\r[ecnt][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ecnt] [2]),
        .Q(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ecnt][3] 
       (.C(clk),
        .CE(\r[ecnt][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ecnt] [3]),
        .Q(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclactive] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[edclactive]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[edclactive_n_0_] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclbcast] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[edclbcast]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[edclbcast]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [0]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][0] ),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][10] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [10]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][10] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][11] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [11]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][11] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][12] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [12]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][12] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][13] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [13]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][13] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][14] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [14]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][14] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][15] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [15]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][15] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][16] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [16]),
        .Q(\m100.u0/ethc0/p_0_in0_in [0]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][17] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [17]),
        .Q(\m100.u0/ethc0/p_0_in0_in [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][18] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [18]),
        .Q(\m100.u0/ethc0/p_0_in0_in [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][19] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [19]),
        .Q(\m100.u0/ethc0/p_0_in0_in [3]),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [1]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][1] ),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][20] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [20]),
        .Q(\m100.u0/ethc0/p_0_in0_in [4]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][21] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [21]),
        .Q(\m100.u0/ethc0/p_0_in0_in [5]),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][22] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [22]),
        .Q(\m100.u0/ethc0/p_0_in0_in [6]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][23] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [23]),
        .Q(\m100.u0/ethc0/p_0_in0_in [7]),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][24] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [24]),
        .Q(\m100.u0/ethc0/p_0_in0_in [8]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][25] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [25]),
        .Q(\m100.u0/ethc0/p_0_in0_in [9]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][26] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [26]),
        .Q(\m100.u0/ethc0/p_0_in0_in [10]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][27] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [27]),
        .Q(\m100.u0/ethc0/p_0_in0_in [11]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][28] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [28]),
        .Q(\m100.u0/ethc0/p_0_in0_in [12]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][29] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [29]),
        .Q(\m100.u0/ethc0/p_0_in0_in [13]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [2]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][2] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][30] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [30]),
        .Q(\m100.u0/ethc0/p_0_in0_in [14]),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][31] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [31]),
        .Q(\m100.u0/ethc0/p_0_in0_in [15]),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [3]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][3] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [4]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][4] ),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [5]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][5] ),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [6]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][6] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [7]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][7] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [8]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][8] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[edclip][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[edclip] ),
        .D(\apbi[pwdata] [9]),
        .Q(\m100.u0/ethc0/r_reg[edclip_n_0_][9] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [0]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][0] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][10] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [10]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][10] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][11] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [11]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][11] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][12] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [12]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][12] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][13] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [13]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][13] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][14] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [14]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][14] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][15] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [15]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][15] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][16] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [16]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][16] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][17] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [17]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][17] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][18] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [18]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][18] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][19] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [19]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][19] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [1]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][1] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][20] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [20]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][20] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][21] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [21]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][21] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][22] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [22]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][22] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][23] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [23]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][23] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][24] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [24]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][24] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][25] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [25]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][25] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][26] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [26]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][26] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][27] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [27]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][27] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][28] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [28]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][28] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][29] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [29]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][29] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [2]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][2] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][30] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [30]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][30] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][31] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [31]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][31] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][32] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [0]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][32] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][33] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [1]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][33] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][34] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [2]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][34] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][35] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [3]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][35] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][36] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [4]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][36] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][37] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [5]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][37] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][38] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [6]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][38] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][39] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [7]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][39] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [3]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][3] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][40] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [8]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][40] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][41] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [9]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][41] ),
        .S(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][42] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [10]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][42] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][43] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [11]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][43] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][44] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [12]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][44] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][45] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [13]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][45] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][46] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [14]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][46] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][47] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [47]),
        .D(\apbi[pwdata] [15]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][47] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [4]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][4] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [5]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][5] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [6]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][6] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [7]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][7] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [8]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][8] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[emacaddr][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[emacaddr] [31]),
        .D(\apbi[pwdata] [9]),
        .Q(\m100.u0/ethc0/r_reg[emacaddr_n_0_][9] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[erenable] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[erenable]_i_1_n_0 ),
        .Q(\m100.u0/erenable ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[erxidle] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[erxidle]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[erxidle]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[etxidle] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/rin ),
        .Q(\m100.u0/ethc0/r_reg[etxidle]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ewr] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\m100.u0/rxwdata [17]),
        .Q(\m100.u0/ethc0/r_reg[ewr]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[gotframe] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[gotframe]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[gotframe_n_0_] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[init_busy] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[init_busy]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[init_busy_n_0_] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][0] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [0]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][0] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][10] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [10]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][10] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][11] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [11]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][11] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][12] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [12]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][12] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][13] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [13]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][13] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][14] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [14]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][14] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][15] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [15]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][15] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][16] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [16]),
        .Q(\m100.u0/ethc0/a [0]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][17] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [17]),
        .Q(\m100.u0/ethc0/a [1]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][1] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [1]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][2] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [2]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][2] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][3] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [3]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][3] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][4] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [4]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][4] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][5] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [5]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][5] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][6] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [6]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][6] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][7] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [7]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][7] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][8] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [8]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][8] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[ipcrc][9] 
       (.C(clk),
        .CE(\r[ipcrc][17]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[ipcrc] [9]),
        .Q(\m100.u0/ethc0/r_reg[ipcrc_n_0_][9] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [0]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][0] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][10] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [10]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][10] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][11] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [11]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][11] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][12] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [12]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][12] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][13] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [13]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][13] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][14] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [14]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][14] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][15] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [15]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][15] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][16] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [16]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][16] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][17] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [17]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][17] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][18] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [18]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][18] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][19] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [19]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][19] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [1]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][20] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [20]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][20] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][21] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [21]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][21] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][22] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [22]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][22] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][23] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [23]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][23] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][24] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [24]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][24] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][25] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [25]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][25] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][26] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [26]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][26] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][27] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [27]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][27] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][28] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [28]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][28] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][29] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [29]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][29] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [2]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][2] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][30] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [30]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][30] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][31] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [31]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][31] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][32] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [0]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][32] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][33] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [1]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][33] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][34] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [2]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][34] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][35] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [3]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][35] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][36] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [4]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][36] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][37] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [5]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][37] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][38] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [6]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][38] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][39] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [7]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][39] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [3]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][3] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][40] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [8]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][40] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][41] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [9]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][41] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][42] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [10]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][42] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][43] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [11]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][43] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][44] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [12]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][44] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][45] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [13]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][45] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][46] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [14]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][46] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][47] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [47]),
        .D(\apbi[pwdata] [15]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][47] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [4]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][4] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [5]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][5] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [6]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][6] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [7]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][7] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [8]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][8] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mac_addr][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[mac_addr] [31]),
        .D(\apbi[pwdata] [9]),
        .Q(\m100.u0/ethc0/r_reg[mac_addr_n_0_][9] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdccnt][0] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/v[mdccnt] [0]),
        .Q(\m100.u0/ethc0/d [0]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdccnt][1] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/v[mdccnt] [1]),
        .Q(\m100.u0/ethc0/d [1]),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdccnt][2] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/v[mdccnt] [2]),
        .Q(\m100.u0/ethc0/d [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdccnt][3] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/v[mdccnt] [3]),
        .Q(\m100.u0/ethc0/d [3]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdccnt][4] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/v[mdccnt] [4]),
        .Q(\m100.u0/ethc0/d [4]),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdccnt][5] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdccnt][5]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/d [5]),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][busy] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[mdio_ctrl][busy]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][busy]__0 ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][0] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][10] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][10]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][10] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][11] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][11]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][11] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][12] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][12]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][12] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][13] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][13]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][13] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][14] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][14]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][14] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][15] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][15]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][15] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][1] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][2] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][2] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][3] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][3] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][4] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][4]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][4] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][5] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][5]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][5] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][6] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][6]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][6] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][7] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][7]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][7] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][8] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][8]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/p_1_in128_in ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][data][9] 
       (.C(clk),
        .CE(apbo),
        .D(\r[mdio_ctrl][data][9]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][9] ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][linkfail] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[mdio_ctrl][linkfail]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][linkfail_n_0_] ),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][phyadr][0] 
       (.C(clk),
        .CE(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .D(\apbi[pwdata] [11]),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][phyadr_n_0_][0] ),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][phyadr][1] 
       (.C(clk),
        .CE(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .D(\apbi[pwdata] [12]),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][phyadr_n_0_][1] ),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][phyadr][2] 
       (.C(clk),
        .CE(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .D(\apbi[pwdata] [13]),
        .Q(\m100.u0/ethc0/data2 ),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][phyadr][3] 
       (.C(clk),
        .CE(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .D(\apbi[pwdata] [14]),
        .Q(\m100.u0/ethc0/data1 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][phyadr][4] 
       (.C(clk),
        .CE(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .D(\apbi[pwdata] [15]),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][phyadr_n_0_][4] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][read] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[mdio_ctrl][read]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][regadr][0] 
       (.C(clk),
        .CE(\r[mdio_ctrl][regadr][4]_i_1_n_0 ),
        .D(\r[mdio_ctrl][regadr][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [0]),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][regadr][1] 
       (.C(clk),
        .CE(\r[mdio_ctrl][regadr][4]_i_1_n_0 ),
        .D(\r[mdio_ctrl][regadr][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [1]),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][regadr][2] 
       (.C(clk),
        .CE(\r[mdio_ctrl][regadr][4]_i_1_n_0 ),
        .D(\r[mdio_ctrl][regadr][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [2]),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][regadr][3] 
       (.C(clk),
        .CE(\r[mdio_ctrl][regadr][4]_i_1_n_0 ),
        .D(\r[mdio_ctrl][regadr][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [3]),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][regadr][4] 
       (.C(clk),
        .CE(\r[mdio_ctrl][regadr][4]_i_1_n_0 ),
        .D(\r[mdio_ctrl][regadr][4]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [4]),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdio_ctrl][write] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[mdio_ctrl][write]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[mdio_ctrl][write]__0 ),
        .R(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdioclk] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[mdioclk]_i_2_n_0 ),
        .Q(\etho[mdc] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdioclkold][0] 
       (.C(clk),
        .CE(apbo),
        .D(\etho[mdc] ),
        .Q(\m100.u0/ethc0/p_1_in143_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdioen] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[mdioen]_i_1_n_0 ),
        .Q(\etho[mdio_oe] ),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdioi] 
       (.C(clk),
        .CE(apbo),
        .D(\ethi[mdio_i] ),
        .Q(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[mdioo] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[mdioo]_i_1_n_0 ),
        .Q(\etho[mdio_o] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[msbgood] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[msbgood]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[msbgood_n_0_] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[nak] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\r[nak]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[nak_n_0_] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[oplen][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\m100.u0/rxwdata [7]),
        .Q(\m100.u0/ethc0/r_reg[oplen_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[oplen][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\m100.u0/rxwdata [8]),
        .Q(\m100.u0/ethc0/r_reg[oplen_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[oplen][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\m100.u0/rxwdata [9]),
        .Q(\m100.u0/ethc0/r_reg[oplen_n_0_][2] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[oplen][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\m100.u0/rxwdata [10]),
        .Q(\m100.u0/ethc0/r_reg[oplen_n_0_][3] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[oplen][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\m100.u0/rxwdata [11]),
        .Q(\m100.u0/ethc0/r_reg[oplen_n_0_][4] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[oplen][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\m100.u0/rxwdata [12]),
        .Q(\m100.u0/ethc0/r_reg[oplen_n_0_][5] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[oplen][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\m100.u0/rxwdata [13]),
        .Q(\m100.u0/ethc0/r_reg[oplen_n_0_][6] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[oplen][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\m100.u0/rxwdata [14]),
        .Q(\m100.u0/ethc0/r_reg[oplen_n_0_][7] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[oplen][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\m100.u0/rxwdata [15]),
        .Q(\m100.u0/ethc0/r_reg[oplen_n_0_][8] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[oplen][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[nak] ),
        .D(\m100.u0/rxwdata [16]),
        .Q(\m100.u0/ethc0/r_reg[oplen_n_0_][9] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[phywr] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[phywr]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntl][0] 
       (.C(clk),
        .CE(\r[rcntl][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntl] [0]),
        .Q(\m100.u0/ewaddressl [0]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntl][1] 
       (.C(clk),
        .CE(\r[rcntl][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntl] [1]),
        .Q(\m100.u0/ewaddressl [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntl][2] 
       (.C(clk),
        .CE(\r[rcntl][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntl] [2]),
        .Q(\m100.u0/ewaddressl [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntl][3] 
       (.C(clk),
        .CE(\r[rcntl][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntl] [3]),
        .Q(\m100.u0/ewaddressl [3]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntl][4] 
       (.C(clk),
        .CE(\r[rcntl][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntl] [4]),
        .Q(\m100.u0/ewaddressl [4]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntl][5] 
       (.C(clk),
        .CE(\r[rcntl][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntl] [5]),
        .Q(\m100.u0/ewaddressl [5]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntl][6] 
       (.C(clk),
        .CE(\r[rcntl][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntl] [6]),
        .Q(\m100.u0/ewaddressl [6]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntm][0] 
       (.C(clk),
        .CE(\r[rcntm][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntm] [0]),
        .Q(\m100.u0/ewaddressm [0]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntm][1] 
       (.C(clk),
        .CE(\r[rcntm][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntm] [1]),
        .Q(\m100.u0/ewaddressm [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntm][2] 
       (.C(clk),
        .CE(\r[rcntm][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntm] [2]),
        .Q(\m100.u0/ewaddressm [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntm][3] 
       (.C(clk),
        .CE(\r[rcntm][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntm] [3]),
        .Q(\m100.u0/ewaddressm [3]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntm][4] 
       (.C(clk),
        .CE(\r[rcntm][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntm] [4]),
        .Q(\m100.u0/ewaddressm [4]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntm][5] 
       (.C(clk),
        .CE(\r[rcntm][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntm] [5]),
        .Q(\m100.u0/ewaddressm [5]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rcntm][6] 
       (.C(clk),
        .CE(\r[rcntm][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rcntm] [6]),
        .Q(\m100.u0/ewaddressm [6]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rfcnt][0] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/v[rfcnt]__0 [0]),
        .Q(\m100.u0/ethc0/r_reg[rfcnt_n_0_][0] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rfcnt][1] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/v[rfcnt]__0 [1]),
        .Q(\m100.u0/ethc0/r_reg[rfcnt_n_0_][1] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rfcnt][2] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/v[rfcnt]__0 [2]),
        .Q(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rfrpnt][0] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/rxraddress [0]),
        .Q(\m100.u0/ethc0/r_reg[rfrpnt_n_0_][0] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rfrpnt][1] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/rxraddress [1]),
        .Q(\m100.u0/ethc0/r_reg[rfrpnt_n_0_][1] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rfwpnt][0] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rfwpnt][0]_i_1_n_0 ),
        .Q(\m100.u0/rxwaddress [0]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rfwpnt][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rfwpnt][1]_i_1_n_0 ),
        .Q(\m100.u0/rxwaddress [1]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][10] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][9]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [10]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][11] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][9]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [11]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][12] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][9]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [12]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][13] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][13]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [13]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][14] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][13]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [14]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][15] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][13]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [15]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][16] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][13]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [16]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][17] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][17]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [17]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][18] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][17]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [18]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][19] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][17]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [19]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][1] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][1]_i_2_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][20] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][17]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [20]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][21] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][21]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [21]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][22] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][21]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [22]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][23] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][21]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [23]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][24] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][21]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [24]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][25] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][25]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [25]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][26] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][25]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [26]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][27] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][25]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [27]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][28] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][25]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [28]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][29] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][29]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [29]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][2] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][1]_i_2_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][30] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][29]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [30]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][31] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][29]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [31]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][3] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][1]_i_2_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [3]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][4] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][1]_i_2_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [4]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][5] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][5]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [5]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][6] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][5]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [6]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][7] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][5]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [7]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][8] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][5]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [8]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][addr][9] 
       (.C(clk),
        .CE(\r[rmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[rmsto][addr][9]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][addr] [9]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][0] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [0]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][0] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][10] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [10]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][10] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][11] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [11]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][11] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][12] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [12]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][12] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][13] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [13]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][13] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][14] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [14]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][14] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][15] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [15]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][15] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][16] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [16]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][16] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][17] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [17]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][17] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][18] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [18]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][18] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][19] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [19]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][19] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][1] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [1]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][20] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [20]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][20] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][21] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [21]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][21] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][22] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [22]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][22] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][23] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [23]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][23] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][24] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [24]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][24] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][25] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [25]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][25] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][26] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [26]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][26] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][27] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [27]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][27] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][28] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [28]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][28] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][29] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [29]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][29] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][2] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [2]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][2] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][30] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [30]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][30] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][31] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/rxrdata [31]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][31] ),
        .R(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][3] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [3]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][3] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][4] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [4]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][4] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][5] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [5]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][5] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][6] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [6]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][6] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][7] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [7]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][7] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][8] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [8]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][8] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][data][9] 
       (.C(clk),
        .CE(\r[rmsto][data][18]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rmsto][data] [9]),
        .Q(\m100.u0/ethc0/r_reg[rmsto][data_n_0_][9] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][req] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rmsto][req]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rmsto][write] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[rmsto][write]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rmsto][write_n_0_] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rpnt][0] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rpnt][0]_i_1_n_0 ),
        .Q(\m100.u0/ewaddressm [7]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rpnt][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rpnt][1]_i_1_n_0 ),
        .Q(\m100.u0/ewaddressm [8]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rstaneg] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[rstaneg]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rstaneg_n_0_] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rstphy] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[rstphy]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rstphy]__0 ),
        .S(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][10] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [10]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][10] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][11] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [11]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][11] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][12] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [12]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][12] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][13] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [13]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][13] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][14] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [14]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][14] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][15] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [15]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][15] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][16] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [16]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][16] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][17] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [17]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][17] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][18] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [18]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][18] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][19] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [19]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][19] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][20] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [20]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][20] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][21] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [21]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][21] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][22] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [22]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][22] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][23] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [23]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][23] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][24] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [24]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][24] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][25] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [25]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][25] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][26] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [26]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][26] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][27] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [27]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][27] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][28] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [28]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][28] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][29] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [29]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][29] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [2]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][2] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][30] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [30]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][30] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][31] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [31]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][31] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [3]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][3] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [4]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][4] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [5]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][5] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [6]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][6] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [7]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][7] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [8]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][8] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxaddr][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxaddr] ),
        .D(\ahbmi[hrdata] [9]),
        .Q(\m100.u0/ethc0/r_reg[rxaddr_n_0_][9] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxburstav] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/v[rxburstav] ),
        .Q(\m100.u0/ethc0/r_reg[rxburstav]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxburstcnt][0] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rxburstcnt][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxburstcnt_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxburstcnt][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rxburstcnt][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxburstcnt_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxbytecount][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxbytecount][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxbytecount]__0 [0]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxbytecount][10] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxbytecount][10]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxbytecount]__0 [10]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxbytecount][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxbytecount][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxbytecount]__0 [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxbytecount][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxbytecount][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxbytecount]__0 [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxbytecount][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxbytecount][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxbytecount]__0 [3]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxbytecount][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxbytecount][4]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxbytecount]__0 [4]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxbytecount][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxbytecount][5]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxbytecount]__0 [5]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxbytecount][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxbytecount][6]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxbytecount]__0 [6]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxbytecount][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxbytecount][7]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxbytecount]__0 [7]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxbytecount][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxbytecount][8]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxbytecount]__0 [8]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxbytecount][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxbytecount][9]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxbytecount]__0 [9]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxcnt][0] 
       (.C(clk),
        .CE(\r[rxcnt][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxcnt] [0]),
        .Q(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxcnt][10] 
       (.C(clk),
        .CE(\r[rxcnt][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxcnt] [10]),
        .Q(\m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxcnt][1] 
       (.C(clk),
        .CE(\r[rxcnt][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxcnt] [1]),
        .Q(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxcnt][2] 
       (.C(clk),
        .CE(\r[rxcnt][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxcnt] [2]),
        .Q(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxcnt][3] 
       (.C(clk),
        .CE(\r[rxcnt][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxcnt] [3]),
        .Q(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxcnt][4] 
       (.C(clk),
        .CE(\r[rxcnt][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxcnt] [4]),
        .Q(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxcnt][5] 
       (.C(clk),
        .CE(\r[rxcnt][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxcnt] [5]),
        .Q(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxcnt][6] 
       (.C(clk),
        .CE(\r[rxcnt][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxcnt] [6]),
        .Q(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxcnt][7] 
       (.C(clk),
        .CE(\r[rxcnt][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxcnt] [7]),
        .Q(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxcnt][8] 
       (.C(clk),
        .CE(\r[rxcnt][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxcnt] [8]),
        .Q(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxcnt][9] 
       (.C(clk),
        .CE(\r[rxcnt][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxcnt] [9]),
        .Q(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxden] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[rxden]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxden]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][10] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [10]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][10] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][11] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [11]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][11] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][12] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [12]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][12] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][13] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [13]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][13] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][14] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [14]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][14] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][15] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [15]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][15] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][16] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [16]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][16] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][17] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [17]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][17] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][18] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [18]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][18] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][19] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [19]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][19] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][20] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [20]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][20] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][21] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [21]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][21] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][22] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [22]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][22] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][23] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [23]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][23] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][24] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [24]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][24] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][25] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [25]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][25] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][26] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [26]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][26] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][27] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [27]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][27] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][28] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [28]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][28] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][29] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [29]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][29] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][30] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [30]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][30] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdesc][31] 
       (.C(clk),
        .CE(\r[rxdesc][31]_i_1_n_0 ),
        .D(\apbi[pwdata] [31]),
        .Q(\m100.u0/ethc0/r_reg[rxdesc_n_0_][31] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdone][0] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/rxo ),
        .Q(\m100.u0/ethc0/r_reg[rxdone] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdoneack] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[rxdoneack]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdoneold] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rxdoneold]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdsel][3] 
       (.C(clk),
        .CE(\r[rxdsel][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxdsel] [3]),
        .Q(\m100.u0/ethc0/r_reg[rxdsel_n_0_][3] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdsel][4] 
       (.C(clk),
        .CE(\r[rxdsel][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxdsel] [4]),
        .Q(\m100.u0/ethc0/r_reg[rxdsel_n_0_][4] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdsel][5] 
       (.C(clk),
        .CE(\r[rxdsel][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxdsel] [5]),
        .Q(\m100.u0/ethc0/r_reg[rxdsel_n_0_][5] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdsel][6] 
       (.C(clk),
        .CE(\r[rxdsel][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxdsel] [6]),
        .Q(\m100.u0/ethc0/r_reg[rxdsel_n_0_][6] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdsel][7] 
       (.C(clk),
        .CE(\r[rxdsel][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxdsel] [7]),
        .Q(\m100.u0/ethc0/r_reg[rxdsel_n_0_][7] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdsel][8] 
       (.C(clk),
        .CE(\r[rxdsel][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxdsel] [8]),
        .Q(\m100.u0/ethc0/r_reg[rxdsel_n_0_][8] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxdsel][9] 
       (.C(clk),
        .CE(\r[rxdsel][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[rxdsel] [9]),
        .Q(\m100.u0/ethc0/r_reg[rxdsel_n_0_][9] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxirq] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[rxirq]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxirq]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxlength][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxlength][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxlength_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxlength][10] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxlength][10]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxlength_n_0_][10] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxlength][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxlength][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxlength_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxlength][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxlength][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxlength][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxlength][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxlength][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxlength][4]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxlength_n_0_][4] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxlength][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxlength][5]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxlength_n_0_][5] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxlength][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxlength][6]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxlength_n_0_][6] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxlength][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxlength][7]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxlength_n_0_][7] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxlength][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxlength][8]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxlength_n_0_][8] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxlength][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[rxbytecount] ),
        .D(\r[rxlength][9]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxlength_n_0_][9] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxstart][0] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/rxo[start] ),
        .Q(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxstart][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rxstart][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxstatus][0] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rxstatus][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxstatus_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxstatus][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rxstatus][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxstatus_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxstatus][2] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rxstatus][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxstatus_n_0_][2] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxstatus][3] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rxstatus][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/p_0_in153_in ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxstatus][4] 
       (.C(clk),
        .CE(apbo),
        .D(\r[rxstatus][4]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/p_1_in4_in ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxwrap] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[rxwrap]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[rxwrap_n_0_] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxwrite][0] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/rxo[write] ),
        .Q(\m100.u0/ethc0/r_reg[rxwrite] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[rxwriteack] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/r_reg[rxwrite] ),
        .Q(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][0]_i_2_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [0]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][10] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][8]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [10]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][11] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][8]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [11]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][12] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][12]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [12]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][13] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][12]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [13]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][0]_i_2_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][0]_i_2_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][0]_i_2_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [3]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][4]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [4]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][4]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [5]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][4]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [6]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][4]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [7]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][8]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [8]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[seq][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[seq] ),
        .D(\r_reg[seq][8]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[seq] [9]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[status][invaddr] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[status][invaddr]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[status][invaddr_n_0_] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[status][rx_err] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[status][rx_err]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[status][rx_err_n_0_] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[status][rx_int] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[status][rx_int]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[status][rx_int_n_0_] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[status][rxahberr] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[status][rxahberr]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[status][rxahberr_n_0_] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[status][toosmall] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[status][toosmall]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[status][toosmall_n_0_] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[status][tx_err] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[status][tx_err]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[status][tx_err_n_0_] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[status][tx_int] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[status][tx_int]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[status][tx_int_n_0_] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[status][txahberr] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[status][txahberr]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[status][txahberr_n_0_] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tarp] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[tarp]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tarp]__0 ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tcnt][0] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/eraddress [0]),
        .Q(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tcnt][1] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/eraddress [1]),
        .Q(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tcnt][2] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/eraddress [2]),
        .Q(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tcnt][3] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/eraddress [3]),
        .Q(\m100.u0/ethc0/r_reg[tcnt_n_0_][3] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tcnt][4] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/eraddress [4]),
        .Q(\m100.u0/ethc0/r_reg[tcnt_n_0_][4] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tcnt][5] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/eraddress [5]),
        .Q(\m100.u0/ethc0/r_reg[tcnt_n_0_][5] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tcnt][6] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/eraddress [6]),
        .Q(\m100.u0/ethc0/r_reg[tcnt_n_0_][6] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tedcl] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[tedcl]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfcnt][0] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tfcnt][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tfcnt_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfcnt][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tfcnt][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tfcnt_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfcnt][2] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tfcnt][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tfcnt_n_0_][2] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfcnt][3] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tfcnt][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tfcnt_n_0_][3] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfcnt][4] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tfcnt][4]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tfcnt_n_0_][4] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfcnt][5] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tfcnt][5]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tfcnt_n_0_][5] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfcnt][6] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tfcnt][6]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tfcnt_n_0_][6] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfcnt][7] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tfcnt][7]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tfcnt_n_0_][7] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfrpnt][0] 
       (.C(clk),
        .CE(\r[tfrpnt][6]_i_1_n_0 ),
        .D(\r[tfrpnt][0]_i_1_n_0 ),
        .Q(\m100.u0/txraddress [0]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfrpnt][1] 
       (.C(clk),
        .CE(\r[tfrpnt][6]_i_1_n_0 ),
        .D(\r[tfrpnt][1]_i_1_n_0 ),
        .Q(\m100.u0/txraddress [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfrpnt][2] 
       (.C(clk),
        .CE(\r[tfrpnt][6]_i_1_n_0 ),
        .D(\r[tfrpnt][2]_i_1_n_0 ),
        .Q(\m100.u0/txraddress [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfrpnt][3] 
       (.C(clk),
        .CE(\r[tfrpnt][6]_i_1_n_0 ),
        .D(\r[tfrpnt][3]_i_1_n_0 ),
        .Q(\m100.u0/txraddress [3]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfrpnt][4] 
       (.C(clk),
        .CE(\r[tfrpnt][6]_i_1_n_0 ),
        .D(\r[tfrpnt][4]_i_1_n_0 ),
        .Q(\m100.u0/txraddress [4]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfrpnt][5] 
       (.C(clk),
        .CE(\r[tfrpnt][6]_i_1_n_0 ),
        .D(\r[tfrpnt][5]_i_1_n_0 ),
        .Q(\m100.u0/txraddress [5]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfrpnt][6] 
       (.C(clk),
        .CE(\r[tfrpnt][6]_i_1_n_0 ),
        .D(\r[tfrpnt][6]_i_2_n_0 ),
        .Q(\m100.u0/txraddress [6]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfwpnt][0] 
       (.C(clk),
        .CE(\r[tfwpnt][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[tfwpnt] [0]),
        .Q(\m100.u0/txwaddress [0]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfwpnt][1] 
       (.C(clk),
        .CE(\r[tfwpnt][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[tfwpnt] [1]),
        .Q(\m100.u0/txwaddress [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfwpnt][2] 
       (.C(clk),
        .CE(\r[tfwpnt][6]_i_1_n_0 ),
        .D(\r[tfwpnt][2]_i_1_n_0 ),
        .Q(\m100.u0/txwaddress [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfwpnt][3] 
       (.C(clk),
        .CE(\r[tfwpnt][6]_i_1_n_0 ),
        .D(\r[tfwpnt][3]_i_1_n_0 ),
        .Q(\m100.u0/txwaddress [3]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfwpnt][4] 
       (.C(clk),
        .CE(\r[tfwpnt][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[tfwpnt] [4]),
        .Q(\m100.u0/txwaddress [4]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfwpnt][5] 
       (.C(clk),
        .CE(\r[tfwpnt][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/v[tfwpnt] [5]),
        .Q(\m100.u0/txwaddress [5]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tfwpnt][6] 
       (.C(clk),
        .CE(\r[tfwpnt][6]_i_1_n_0 ),
        .D(\r[tfwpnt][6]_i_2_n_0 ),
        .Q(\m100.u0/txwaddress [6]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][10] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][9]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [10]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][11] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][9]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [11]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][12] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][9]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [12]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][13] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][13]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [13]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][14] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][13]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [14]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][15] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][13]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [15]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][16] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][13]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [16]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][17] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][17]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [17]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][18] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][17]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [18]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][19] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][17]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [19]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][1] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][1]_i_2_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][20] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][17]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [20]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][21] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][21]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [21]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][22] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][21]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [22]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][23] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][21]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [23]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][24] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][21]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [24]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][25] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][25]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [25]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][26] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][25]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [26]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][27] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][25]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [27]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][28] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][25]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [28]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][29] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][29]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [29]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][2] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][1]_i_2_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][30] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][29]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [30]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][31] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][29]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [31]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][3] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][1]_i_2_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [3]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][4] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][1]_i_2_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [4]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][5] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][5]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [5]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][6] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][5]_i_1_n_6 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [6]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][7] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][5]_i_1_n_5 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [7]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][8] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][5]_i_1_n_4 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [8]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][addr][9] 
       (.C(clk),
        .CE(\r[tmsto][addr][1]_i_1_n_0 ),
        .D(\r_reg[tmsto][addr][9]_i_1_n_7 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][addr] [9]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [0]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][0] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][10] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [10]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][10] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][11] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [11]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][11] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][12] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [12]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][12] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][13] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [13]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][13] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][14] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tmsto][data][14]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][14] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][15] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tmsto][data][15]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][15] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][16] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [16]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][16] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][17] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [17]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][17] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][18] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [18]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][18] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][19] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [19]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][19] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [1]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][1] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][20] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [20]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][20] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][21] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [21]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][21] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][22] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [22]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][22] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][23] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [23]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][23] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][24] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [24]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][24] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][25] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [25]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][25] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][26] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [26]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][26] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][27] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [27]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][27] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][28] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [28]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][28] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][29] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [29]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][29] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [2]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][2] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][30] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [30]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][30] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][31] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [31]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][31] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [3]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][3] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [4]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][4] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [5]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][5] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [6]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][6] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [7]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][7] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [8]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][8] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][data][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tmsto][data] ),
        .D(\m100.u0/erdata [9]),
        .Q(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][9] ),
        .R(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][req] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tmsto][req]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tmsto][write] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[tmsto][write]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tmsto][write_n_0_] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tnak] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[tnak]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[tnak]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tpnt][0] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tpnt][0]_i_1_n_0 ),
        .Q(\m100.u0/eraddress [7]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[tpnt][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[tpnt][1]_i_1_n_0 ),
        .Q(\m100.u0/eraddress [8]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][10] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][10]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [8]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][11] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][11]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [9]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][12] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][12]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [10]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][13] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][13]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [11]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][14] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][14]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [12]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][15] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][15]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [13]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][16] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][16]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [14]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][17] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][17]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [15]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][18] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][18]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [16]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][19] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][19]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [17]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][20] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][20]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [18]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][21] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][21]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [19]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][22] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][22]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [20]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][23] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][23]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [21]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][24] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][24]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [22]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][25] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][25]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [23]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][26] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][26]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [24]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][27] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][27]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [25]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][28] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][28]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [26]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][29] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][29]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [27]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][2] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [0]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][30] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][30]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [28]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][31] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][31]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [29]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][3] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [1]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][4] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][4]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [2]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][5] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][5]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [3]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][6] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][6]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [4]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][7] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][7]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [5]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][8] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][8]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [6]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txaddr][9] 
       (.C(clk),
        .CE(\r[txaddr][31]_i_1_n_0 ),
        .D(\r[txaddr][9]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txaddr]__0 [7]),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txburstav] 
       (.C(clk),
        .CE(apbo),
        .D(\r[txburstav]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txburstav]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txburstcnt][0] 
       (.C(clk),
        .CE(apbo),
        .D(\r[txburstcnt][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txburstcnt_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txburstcnt][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[txburstcnt][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txburstcnt_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txcnt][0] 
       (.C(clk),
        .CE(\r[txcnt][10]_i_1_n_0 ),
        .D(\r[txcnt][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txcnt][10] 
       (.C(clk),
        .CE(\r[txcnt][10]_i_1_n_0 ),
        .D(\r[txcnt][10]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txcnt_n_0_][10] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txcnt][1] 
       (.C(clk),
        .CE(\r[txcnt][10]_i_1_n_0 ),
        .D(\r[txcnt][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txcnt][2] 
       (.C(clk),
        .CE(\r[txcnt][10]_i_1_n_0 ),
        .D(\r[txcnt][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txcnt][3] 
       (.C(clk),
        .CE(\r[txcnt][10]_i_1_n_0 ),
        .D(\r[txcnt][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txcnt][4] 
       (.C(clk),
        .CE(\r[txcnt][10]_i_1_n_0 ),
        .D(\r[txcnt][4]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txcnt][5] 
       (.C(clk),
        .CE(\r[txcnt][10]_i_1_n_0 ),
        .D(\r[txcnt][5]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txcnt][6] 
       (.C(clk),
        .CE(\r[txcnt][10]_i_1_n_0 ),
        .D(\r[txcnt][6]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txcnt_n_0_][6] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txcnt][7] 
       (.C(clk),
        .CE(\r[txcnt][10]_i_1_n_0 ),
        .D(\r[txcnt][7]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txcnt_n_0_][7] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txcnt][8] 
       (.C(clk),
        .CE(\r[txcnt][10]_i_1_n_0 ),
        .D(\r[txcnt][8]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txcnt_n_0_][8] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txcnt][9] 
       (.C(clk),
        .CE(\r[txcnt][10]_i_1_n_0 ),
        .D(\r[txcnt][9]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txcnt_n_0_][9] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [0]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][0] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][10] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [10]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][10] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][11] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [11]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][11] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][12] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [12]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][12] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][13] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [13]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][13] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][14] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [14]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][14] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][15] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [15]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][15] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][16] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [16]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][16] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][17] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [17]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][17] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][18] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [18]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][18] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][19] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [19]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][19] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [1]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][20] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [20]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][20] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][21] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [21]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][21] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][22] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [22]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][22] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][23] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [23]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][23] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][24] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [24]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][24] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][25] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [25]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][25] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][26] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [26]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][26] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][27] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [27]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][27] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][28] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [28]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][28] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][29] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [29]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][29] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [2]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][2] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][30] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [30]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][30] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][31] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [31]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][31] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [3]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][3] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [4]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][4] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [5]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][5] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [6]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][6] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [7]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][7] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [8]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][8] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdata][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/txrdata [9]),
        .Q(\m100.u0/ethc0/r_reg[txdata_n_0_][9] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdataav] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/txrenable ),
        .Q(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txden] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[txden]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txden]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][10] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [10]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [0]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][11] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [11]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [1]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][12] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [12]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [2]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][13] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [13]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [3]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][14] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [14]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [4]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][15] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [15]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [5]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][16] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [16]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [6]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][17] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [17]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [7]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][18] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [18]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [8]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][19] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [19]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [9]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][20] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [20]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [10]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][21] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [21]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [11]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][22] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [22]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [12]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][23] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [23]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [13]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][24] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [24]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [14]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][25] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [25]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [15]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][26] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [26]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [16]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][27] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [27]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [17]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][28] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [28]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [18]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][29] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [29]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [19]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][30] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [30]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [20]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdesc][31] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[txdsel] ),
        .D(\apbi[pwdata] [31]),
        .Q(\m100.u0/ethc0/r_reg[txdesc]__0 [21]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdone][0] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/txo ),
        .Q(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdone][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[txdone][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdsel][3] 
       (.C(clk),
        .CE(\r[txdsel][9]_i_1_n_0 ),
        .D(\r[txdsel][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txdsel_n_0_][3] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdsel][4] 
       (.C(clk),
        .CE(\r[txdsel][9]_i_1_n_0 ),
        .D(\r[txdsel][4]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txdsel_n_0_][4] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdsel][5] 
       (.C(clk),
        .CE(\r[txdsel][9]_i_1_n_0 ),
        .D(\r[txdsel][5]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txdsel_n_0_][5] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdsel][6] 
       (.C(clk),
        .CE(\r[txdsel][9]_i_1_n_0 ),
        .D(\r[txdsel][6]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txdsel_n_0_][6] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdsel][7] 
       (.C(clk),
        .CE(\r[txdsel][9]_i_1_n_0 ),
        .D(\r[txdsel][7]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txdsel_n_0_][7] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdsel][8] 
       (.C(clk),
        .CE(\r[txdsel][9]_i_1_n_0 ),
        .D(\r[txdsel][8]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txdsel_n_0_][8] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdsel][9] 
       (.C(clk),
        .CE(\r[txdsel][9]_i_1_n_0 ),
        .D(\r[txdsel][9]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txdsel_n_0_][9] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdstate][0] 
       (.C(clk),
        .CE(apbo),
        .D(\r[txdstate][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdstate][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[txdstate][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdstate][2] 
       (.C(clk),
        .CE(apbo),
        .D(\r[txdstate][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txdstate][3] 
       (.C(clk),
        .CE(apbo),
        .D(\r[txdstate][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txirq] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[txirq]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txirq]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txirqgen] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[txirqgen]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txirqgen_n_0_] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txlength][0] 
       (.C(clk),
        .CE(\r[txlength][10]_i_1_n_0 ),
        .D(\r[txlength][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txlength_n_0_][0] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txlength][10] 
       (.C(clk),
        .CE(\r[txlength][10]_i_1_n_0 ),
        .D(\r[txlength][10]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txlength_n_0_][10] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txlength][1] 
       (.C(clk),
        .CE(\r[txlength][10]_i_1_n_0 ),
        .D(\r[txlength][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txlength_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txlength][2] 
       (.C(clk),
        .CE(\r[txlength][10]_i_1_n_0 ),
        .D(\r[txlength][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txlength_n_0_][2] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txlength][3] 
       (.C(clk),
        .CE(\r[txlength][10]_i_1_n_0 ),
        .D(\r[txlength][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txlength_n_0_][3] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txlength][4] 
       (.C(clk),
        .CE(\r[txlength][10]_i_1_n_0 ),
        .D(\r[txlength][4]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txlength_n_0_][4] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txlength][5] 
       (.C(clk),
        .CE(\r[txlength][10]_i_1_n_0 ),
        .D(\r[txlength][5]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txlength_n_0_][5] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txlength][6] 
       (.C(clk),
        .CE(\r[txlength][10]_i_1_n_0 ),
        .D(\r[txlength][6]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txlength_n_0_][6] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txlength][7] 
       (.C(clk),
        .CE(\r[txlength][10]_i_1_n_0 ),
        .D(\r_reg[txlength][7]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txlength_n_0_][7] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txlength][8] 
       (.C(clk),
        .CE(\r[txlength][10]_i_1_n_0 ),
        .D(\r[txlength][8]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txlength_n_0_][8] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txlength][9] 
       (.C(clk),
        .CE(\r[txlength][10]_i_1_n_0 ),
        .D(\r_reg[txlength][9]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txlength_n_0_][9] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txread][0] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/txo[read] ),
        .Q(\m100.u0/ethc0/r_reg[txread] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txreadack] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/r_reg[txread] ),
        .Q(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txrestart][0] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/ethc0/txo[restart] ),
        .Q(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txrestart][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[txrestart][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txstart] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[txstart]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txstart]__0 ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txstart_sync] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[txstart_sync]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txstart_sync_n_0_] ),
        .R(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txstatus][0] 
       (.C(clk),
        .CE(apbo),
        .D(\r[txstatus][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txstatus_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txstatus][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[txstatus][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txstatus_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txvalid] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[tfrpnt]1 ),
        .D(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .Q(\m100.u0/ethc0/r_reg[txvalid_n_0_] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[txwrap] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[txwrap]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[txwrap_n_0_] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][0] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [0]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][10] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [10]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][10] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][11] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [11]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][11] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][12] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [12]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][12] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][13] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [13]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][13] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][14] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [14]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][14] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][15] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [15]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][15] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][1] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [1]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][2] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [2]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][2] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][3] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [3]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][3] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][4] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [4]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][4] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][5] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [5]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][5] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][6] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [6]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][6] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][7] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [7]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][7] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][8] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [8]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][8] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[udpsrc][9] 
       (.C(clk),
        .CE(\m100.u0/ethc0/v[udpsrc] ),
        .D(\m100.u0/rxwdata [9]),
        .Q(\m100.u0/ethc0/r_reg[udpsrc_n_0_][9] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[write][0] 
       (.C(clk),
        .CE(apbo),
        .D(\r[write][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[write_n_0_][0] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[write][1] 
       (.C(clk),
        .CE(apbo),
        .D(\r[write][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[write_n_0_][1] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[write][2] 
       (.C(clk),
        .CE(apbo),
        .D(\r[write][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[write_n_0_][2] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[write][3] 
       (.C(clk),
        .CE(apbo),
        .D(\r[write][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[write_n_0_][3] ),
        .R(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/r_reg[writeok] 
       (.C(clk),
        .CE(apbo),
        .D(\m100.u0/r[writeok]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/r_reg[writeok_n_0_] ),
        .S(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/FSM_sequential_gmiimode0.r_reg[rx_state][0] 
       (.C(ethi),
        .CE(\FSM_sequential_gmiimode0.r[rx_state][3]_i_2_n_0 ),
        .D(\FSM_sequential_gmiimode0.r[rx_state][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [0]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/FSM_sequential_gmiimode0.r_reg[rx_state][1] 
       (.C(ethi),
        .CE(\FSM_sequential_gmiimode0.r[rx_state][3]_i_2_n_0 ),
        .D(\FSM_sequential_gmiimode0.r_reg ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [1]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/FSM_sequential_gmiimode0.r_reg[rx_state][2] 
       (.C(ethi),
        .CE(\FSM_sequential_gmiimode0.r[rx_state][3]_i_2_n_0 ),
        .D(\FSM_sequential_gmiimode0.r[rx_state][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [2]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/FSM_sequential_gmiimode0.r_reg[rx_state][3] 
       (.C(ethi),
        .CE(\FSM_sequential_gmiimode0.r[rx_state][3]_i_2_n_0 ),
        .D(\FSM_sequential_gmiimode0.r[rx_state][3]_i_3_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rx_state] [3]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r[lentype][3]_i_2 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/d [19]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r[lentype][3]_i_3 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/d [18]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r[lentype][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r[lentype][3]_i_4 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/d [17]),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r[lentype][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[act] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[byte_count][0] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [0]),
        .Q(\m100.u0/ethc0/rxo[byte_count] [0]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[byte_count][10] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [10]),
        .Q(\m100.u0/ethc0/rxo[byte_count] [10]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[byte_count][1] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [1]),
        .Q(\m100.u0/ethc0/rxo[byte_count] [1]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[byte_count][2] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [2]),
        .Q(\m100.u0/ethc0/rxo[byte_count] [2]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[byte_count][3] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [3]),
        .Q(\m100.u0/ethc0/rxo[byte_count] [3]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[byte_count][4] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [4]),
        .Q(\m100.u0/ethc0/rxo[byte_count] [4]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[byte_count][5] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [5]),
        .Q(\m100.u0/ethc0/rxo[byte_count] [5]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[byte_count][6] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [6]),
        .Q(\m100.u0/ethc0/rxo[byte_count] [6]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[byte_count][7] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [7]),
        .Q(\m100.u0/ethc0/rxo[byte_count] [7]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[byte_count][8] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [8]),
        .Q(\m100.u0/ethc0/rxo[byte_count] [8]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[byte_count][9] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[byte_count] [9]),
        .Q(\m100.u0/ethc0/rxo[byte_count] [9]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[cnt] [0]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[cnt] [1]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt][2] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[cnt] [2]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt][3] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/v[cnt] [3]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[cnt_n_0_][3] ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][0] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [0]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][0] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][10] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [10]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_16_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][11] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [11]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_17_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][12] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [12]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_18_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][13] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [13]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_19_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][14] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [14]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_20_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][15] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [15]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_22_in55_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][16] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [16]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_31_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][17] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [17]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_32_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][18] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [18]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_23_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][19] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [19]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_24_in59_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][1] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [1]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][20] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [20]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_25_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][21] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [21]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_26_in64_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][22] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [22]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_27_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][23] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [23]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_28_in69_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][24] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [24]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_29_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][25] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [25]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_30_in72_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][26] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [26]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_33_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][27] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [27]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][27] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][28] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [28]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in18_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][29] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [29]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in15_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][2] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [2]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][2] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][30] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [30]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in12_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][31] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [31]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_0_in10_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][3] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [3]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_9_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][4] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [4]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_10_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][5] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [5]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_11_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][6] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [6]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc_n_0_][6] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][7] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [7]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_13_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][8] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [8]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_14_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[crc][9] 
       (.C(ethi),
        .CE(\gmiimode0.r[crc][31]_i_1__0_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rin[crc] [9]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_15_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][0] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [3]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][0] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][10] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [11]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][10] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][11] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [11]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][11] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][12] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [15]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][12] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][13] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [15]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][13] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][14] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [15]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][14] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][15] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [15]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][15] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][16] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [19]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [16]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][17] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [19]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [17]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][18] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [19]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [18]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][19] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [19]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [19]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][1] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [3]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][20] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [23]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [20]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][21] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [23]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [21]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][22] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [23]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [22]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][23] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [23]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [23]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][24] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [27]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [24]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][25] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [27]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [25]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][26] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [27]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [26]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][27] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [27]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [27]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][28] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [31]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [28]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][29] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [31]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [29]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][2] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [3]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][2] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][30] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [31]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [30]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][31] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [31]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/d [31]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][3] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [3]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][3] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][4] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [7]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][4] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][5] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [7]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][5] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][6] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [7]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][6] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][7] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [7]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][7] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][8] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [11]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][8] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data][9] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[data] [11]),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][9] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][0] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][0] ),
        .Q(\m100.u0/rxwdata [0]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][10] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][10] ),
        .Q(\m100.u0/rxwdata [10]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][11] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][11] ),
        .Q(\m100.u0/rxwdata [11]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][12] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][12] ),
        .Q(\m100.u0/rxwdata [12]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][13] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][13] ),
        .Q(\m100.u0/rxwdata [13]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][14] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][14] ),
        .Q(\m100.u0/rxwdata [14]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][15] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][15] ),
        .Q(\m100.u0/rxwdata [15]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][16] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [16]),
        .Q(\m100.u0/rxwdata [16]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][17] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [17]),
        .Q(\m100.u0/rxwdata [17]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][18] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [18]),
        .Q(\m100.u0/rxwdata [18]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][19] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [19]),
        .Q(\m100.u0/rxwdata [19]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][1] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][1] ),
        .Q(\m100.u0/rxwdata [1]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][20] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [20]),
        .Q(\m100.u0/rxwdata [20]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][21] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [21]),
        .Q(\m100.u0/rxwdata [21]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][22] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [22]),
        .Q(\m100.u0/rxwdata [22]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][23] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [23]),
        .Q(\m100.u0/rxwdata [23]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][24] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [24]),
        .Q(\m100.u0/rxwdata [24]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][25] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [25]),
        .Q(\m100.u0/rxwdata [25]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][26] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [26]),
        .Q(\m100.u0/rxwdata [26]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][27] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [27]),
        .Q(\m100.u0/rxwdata [27]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][28] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [28]),
        .Q(\m100.u0/rxwdata [28]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][29] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [29]),
        .Q(\m100.u0/rxwdata [29]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][2] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][2] ),
        .Q(\m100.u0/rxwdata [2]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][30] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [30]),
        .Q(\m100.u0/rxwdata [30]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][31] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/d [31]),
        .Q(\m100.u0/rxwdata [31]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][3] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][3] ),
        .Q(\m100.u0/rxwdata [3]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][4] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][4] ),
        .Q(\m100.u0/rxwdata [4]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][5] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][5] ),
        .Q(\m100.u0/rxwdata [5]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][6] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][6] ),
        .Q(\m100.u0/rxwdata [6]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][7] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][7] ),
        .Q(\m100.u0/rxwdata [7]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][8] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][8] ),
        .Q(\m100.u0/rxwdata [8]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dataout][9] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[dataout] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[data_n_0_][9] ),
        .Q(\m100.u0/rxwdata [9]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[done] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[done]_i_1__0_n_0 ),
        .Q(\m100.u0/ethc0/rxo ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[done_ack][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[done_ack_n_0_][0] ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dv] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[dv]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[dv]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[en] 
       (.C(ethi),
        .CE(apbo),
        .D(\ethi[rx_crs] ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[en]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[enold] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[enold]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[enold]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[got4b]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[got4b]__0 ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[gotframe] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[gotframe]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rxo[gotframe] ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][0] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [0]),
        .Q(\m100.u0/ethc0/rxo[lentype] [0]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][10] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [10]),
        .Q(\m100.u0/ethc0/rxo[lentype] [10]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][11] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [11]),
        .Q(\m100.u0/ethc0/rxo[lentype] [11]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][11]_i_1 
       (.CI(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][7]_i_1_n_0 ),
        .CO({\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][11]_i_1_n_0 ,\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][11]_i_1_n_1 ,\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][11]_i_1_n_2 ,\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][11]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [11:8]),
        .S(\m100.u0/ethc0/rx_rmii1.rx0/d [27:24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][12] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [12]),
        .Q(\m100.u0/ethc0/rxo[lentype] [12]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][13] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [13]),
        .Q(\m100.u0/ethc0/rxo[lentype] [13]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][14] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [14]),
        .Q(\m100.u0/ethc0/rxo[lentype] [14]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][15] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [15]),
        .Q(\m100.u0/ethc0/rxo[lentype] [15]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][15]_i_2 
       (.CI(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][11]_i_1_n_0 ),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [15:12]),
        .S(\m100.u0/ethc0/rx_rmii1.rx0/d [31:28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][1] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [1]),
        .Q(\m100.u0/ethc0/rxo[lentype] [1]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][2] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [2]),
        .Q(\m100.u0/ethc0/rxo[lentype] [2]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][3] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [3]),
        .Q(\m100.u0/ethc0/rxo[lentype] [3]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][3]_i_1 
       (.CI(etho),
        .CO({\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][3]_i_1_n_0 ,\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][3]_i_1_n_1 ,\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][3]_i_1_n_2 ,\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][3]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/rx_rmii1.rx0/d [19:17],etho}),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [3:0]),
        .S({\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r ,\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r[lentype][3]_i_3_n_0 ,\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r[lentype][3]_i_4_n_0 ,\m100.u0/ethc0/rx_rmii1.rx0/d [16]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][4] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [4]),
        .Q(\m100.u0/ethc0/rxo[lentype] [4]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][5] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [5]),
        .Q(\m100.u0/ethc0/rxo[lentype] [5]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][6] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [6]),
        .Q(\m100.u0/ethc0/rxo[lentype] [6]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][7] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [7]),
        .Q(\m100.u0/ethc0/rxo[lentype] [7]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][7]_i_1 
       (.CI(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][3]_i_1_n_0 ),
        .CO({\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][7]_i_1_n_0 ,\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][7]_i_1_n_1 ,\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][7]_i_1_n_2 ,\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][7]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [7:4]),
        .S(\m100.u0/ethc0/rx_rmii1.rx0/d [23:20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][8] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [8]),
        .Q(\m100.u0/ethc0/rxo[lentype] [8]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[lentype][9] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/rx_rmii1.rx0/v[lentype] ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/plusOp [9]),
        .Q(\m100.u0/ethc0/rxo[lentype] [9]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[ltfound] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[ltfound]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[ltfound_n_0_] ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[odd_nibble] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[odd_nibble]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[odd_nibble_n_0_] ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxd2][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[rxd2][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxd2][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[rxd2][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxd][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\ethi[rxd] [0]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxd][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\ethi[rxd] [1]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp][0] 
       (.C(ethi),
        .CE(\gmiimode0.r[rxdp][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [24]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp_n_0_][0] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp][1] 
       (.C(ethi),
        .CE(\gmiimode0.r[rxdp][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [25]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp][2] 
       (.C(ethi),
        .CE(\gmiimode0.r[rxdp][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [26]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp_n_0_][2] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp][3] 
       (.C(ethi),
        .CE(\gmiimode0.r[rxdp][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/p_4_in [27]),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[rxdp_n_0_][3] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[start] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[start]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[start]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[status][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[status][0]_i_1__0_n_0 ),
        .Q(\m100.u0/ethc0/rxo[status] [0]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[status][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[status][1]_i_1__0_n_0 ),
        .Q(\m100.u0/ethc0/rxo[status] [1]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[status][2] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[status][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rxo[status] [2]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[status][3] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[status][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rxo[status] [3]),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[sync_start] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[sync_start]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rxo[start] ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[write] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[write]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/rxo[write] ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[write_ack][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[write_ack] ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[zero]_i_1__0_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[zero]__0 ),
        .R(\FSM_sequential_gmiimode0.r[rx_state][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg[0] 
       (.C(ethi),
        .CE(apbo),
        .CLR(\r[ctrl][speed]_i_1_n_0 ),
        .D(apbo),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg_n_0_ ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg[1] 
       (.C(ethi),
        .CE(apbo),
        .CLR(\r[ctrl][speed]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg_n_0_ ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg_n_0_[1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg[2] 
       (.C(ethi),
        .CE(apbo),
        .CLR(\r[ctrl][speed]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg_n_0_[1] ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/p_1_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg[3] 
       (.C(ethi),
        .CE(apbo),
        .CLR(\r[ctrl][speed]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/p_1_in ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg[4] 
       (.C(ethi),
        .CE(apbo),
        .CLR(\r[ctrl][speed]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/p_0_in ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/rstout0 
       (.I0(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/p_1_in ),
        .I1(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/r_reg_n_0_[4] ),
        .I2(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/p_0_in ),
        .O(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/rstout0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \m100.u0/ethc0/rx_rmii1.rx0/rx_rst/rstout_reg 
       (.C(ethi),
        .CE(apbo),
        .CLR(\r[ctrl][speed]_i_1_n_0 ),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/rx_rst/rstout0_n_0 ),
        .Q(\m100.u0/ethc0/rx_rmii1.rx0/rxrst ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/FSM_sequential_gmiimode0.r_reg[def_state][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\FSM_sequential_gmiimode0.r ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [0]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/FSM_sequential_gmiimode0.r_reg[def_state][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\FSM_sequential_gmiimode0.r[def_state][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [1]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/FSM_sequential_gmiimode0.r_reg[def_state][2] 
       (.C(ethi),
        .CE(apbo),
        .D(\FSM_sequential_gmiimode0.r[def_state][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[def_state] [2]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/FSM_sequential_gmiimode0.r_reg[main_state][0] 
       (.C(ethi),
        .CE(\FSM_sequential_gmiimode0.r[main_state][3]_i_1_n_0 ),
        .D(\FSM_sequential_gmiimode0.r[main_state][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [0]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/FSM_sequential_gmiimode0.r_reg[main_state][1] 
       (.C(ethi),
        .CE(\FSM_sequential_gmiimode0.r[main_state][3]_i_1_n_0 ),
        .D(\FSM_sequential_gmiimode0.r[main_state][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [1]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/FSM_sequential_gmiimode0.r_reg[main_state][2] 
       (.C(ethi),
        .CE(\FSM_sequential_gmiimode0.r[main_state][3]_i_1_n_0 ),
        .D(\FSM_sequential_gmiimode0.r[main_state][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [2]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/FSM_sequential_gmiimode0.r_reg[main_state][3] 
       (.C(ethi),
        .CE(\FSM_sequential_gmiimode0.r[main_state][3]_i_1_n_0 ),
        .D(\FSM_sequential_gmiimode0.r[main_state][3]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[main_state] [3]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count][0] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_2_n_0 ),
        .D(\gmiimode0.r[byte_count][0]_i_1__0_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg ),
        .S(\gmiimode0.r[byte_count][10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count][10] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_2_n_0 ),
        .D(\gmiimode0.r[byte_count][10]_i_3_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][10] ),
        .S(\gmiimode0.r[byte_count][10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count][1] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_2_n_0 ),
        .D(\gmiimode0.r[byte_count][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][1] ),
        .S(\gmiimode0.r[byte_count][10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count][2] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_2_n_0 ),
        .D(\gmiimode0.r[byte_count][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][2] ),
        .S(\gmiimode0.r[byte_count][10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count][3] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_2_n_0 ),
        .D(\gmiimode0.r[byte_count][3]_i_1__0_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][3] ),
        .S(\gmiimode0.r[byte_count][10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count][4] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_2_n_0 ),
        .D(\gmiimode0.r[byte_count][4]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][4] ),
        .S(\gmiimode0.r[byte_count][10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count][5] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_2_n_0 ),
        .D(\gmiimode0.r[byte_count][5]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][5] ),
        .S(\gmiimode0.r[byte_count][10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count][6] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_2_n_0 ),
        .D(\gmiimode0.r[byte_count][6]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][6] ),
        .S(\gmiimode0.r[byte_count][10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count][7] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_2_n_0 ),
        .D(\gmiimode0.r[byte_count][7]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][7] ),
        .S(\gmiimode0.r[byte_count][10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count][8] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_2_n_0 ),
        .D(\gmiimode0.r[byte_count][8]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][8] ),
        .S(\gmiimode0.r[byte_count][10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count][9] 
       (.C(ethi),
        .CE(\gmiimode0.r[byte_count][10]_i_2_n_0 ),
        .D(\gmiimode0.r[byte_count][9]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[byte_count_n_0_][9] ),
        .S(\gmiimode0.r[byte_count][10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt][0] 
       (.C(ethi),
        .CE(\gmiimode0.r[cnt][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[cnt] [0]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][0] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt][1] 
       (.C(ethi),
        .CE(\gmiimode0.r[cnt][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[cnt] [1]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][1] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt][2] 
       (.C(ethi),
        .CE(\gmiimode0.r[cnt][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[cnt] [2]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][2] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt][3] 
       (.C(ethi),
        .CE(\gmiimode0.r[cnt][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[cnt] [3]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[cnt_n_0_][3] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [0]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][0] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][10] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [10]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][10] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][11] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [11]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_17_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][12] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [12]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][12] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][13] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [13]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][13] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][14] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [14]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][14] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][15] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [15]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_22_in55_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][16] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [16]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_31_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][17] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [17]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_32_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][18] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [18]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_23_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][19] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [19]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_24_in59_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [1]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][20] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [20]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_25_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][21] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [21]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_26_in64_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][22] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [22]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_27_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][23] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [23]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_28_in69_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][24] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [24]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][24] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][25] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [25]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_30_in72_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][26] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [26]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_33_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][27] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [27]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][27] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][28] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [28]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in18_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][29] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [29]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in15_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][2] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [2]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_8_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][30] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [30]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in12_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][31] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [31]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in10_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][3] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [3]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_9_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][4] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [4]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_10_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][5] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [5]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_11_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][6] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [6]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_12_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][7] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [7]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_13_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][8] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [8]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_14_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc][9] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[crc] [9]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_n_0_][9] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[crc_en]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crc_en]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/rx_rmii1.rx0/gmiimode0.r_reg[en]__0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/rin ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_act] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[crs_act]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_act]__1 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_prev] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/rin ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[crs_prev_n_0_] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][0] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][0] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][0] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][10] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][10] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_15_in [2]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][11] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][11] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_15_in [3]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][12] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][12] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_19_in [0]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][13] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][13] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_19_in [1]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][14] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][14] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_19_in [2]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][15] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][15] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_19_in [3]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][16] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][16] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_16_in [0]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][17] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][17] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_16_in [1]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][18] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][18] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_16_in [2]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][19] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][19] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_16_in [3]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][1] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][1] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][20] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][20] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_20_in [0]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][21] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][21] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_20_in [1]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][22] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][22] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_20_in [2]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][23] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][23] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_20_in [3]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][24] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][24] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][24] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][25] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][25] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][25] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][26] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][26] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][26] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][27] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][27] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][27] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][28] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][28] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][28] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][29] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][29] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][29] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][2] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][2] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][2] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][30] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][30] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][30] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][31] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][31] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][31] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][3] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][3] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data_n_0_][3] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][4] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][4] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_18_in [0]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][5] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][5] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_18_in [1]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][6] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][6] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_18_in [2]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][7] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][7] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_18_in [3]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][8] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][8] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_15_in [0]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[data][9] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[data] ),
        .D(\m100.u0/ethc0/r_reg[txdata_n_0_][9] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_15_in [1]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[deferring] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[deferring]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[deferring_n_0_] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[delay_val][0] 
       (.C(ethi),
        .CE(\gmiimode0.r[delay_val][9]_i_1_n_0 ),
        .D(\gmiimode0.r[delay_val][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/v [0]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[delay_val][1] 
       (.C(ethi),
        .CE(\gmiimode0.r[delay_val][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [1]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/v [1]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[delay_val][2] 
       (.C(ethi),
        .CE(\gmiimode0.r[delay_val][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [2]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/v [2]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[delay_val][3] 
       (.C(ethi),
        .CE(\gmiimode0.r[delay_val][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [3]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/v [3]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[delay_val][4] 
       (.C(ethi),
        .CE(\gmiimode0.r[delay_val][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [4]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/v [4]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[delay_val][5] 
       (.C(ethi),
        .CE(\gmiimode0.r[delay_val][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [5]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/v [5]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[delay_val][6] 
       (.C(ethi),
        .CE(\gmiimode0.r[delay_val][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [6]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/v [6]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[delay_val][7] 
       (.C(ethi),
        .CE(\gmiimode0.r[delay_val][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [7]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/v [7]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[delay_val][8] 
       (.C(ethi),
        .CE(\gmiimode0.r[delay_val][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [8]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/v [8]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[delay_val][9] 
       (.C(ethi),
        .CE(\gmiimode0.r[delay_val][9]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[delay_val] [9]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/v [9]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[done] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[done]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/txo ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[fullduplex][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/p_6_in [4]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/rin[fullduplex] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[fullduplex][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/rin[fullduplex] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in38_in ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[icnt][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][0] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[icnt][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[icnt_n_0_][1] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[ifg_cycls][0] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[ifg_cycls] ),
        .D(\gmiimode0.r[ifg_cycls][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/d [0]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[ifg_cycls][1] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[ifg_cycls] ),
        .D(\gmiimode0.r[ifg_cycls][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/d [1]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[ifg_cycls][2] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[ifg_cycls] ),
        .D(\gmiimode0.r[ifg_cycls][2]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/d [2]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[ifg_cycls][3] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[ifg_cycls] ),
        .D(\gmiimode0.r[ifg_cycls][3]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/d [3]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[ifg_cycls][4] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[ifg_cycls] ),
        .D(\gmiimode0.r[ifg_cycls][4]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/d [4]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[ifg_cycls][5] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[ifg_cycls] ),
        .D(\gmiimode0.r[ifg_cycls][5]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/d [5]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[ifg_cycls][6] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[ifg_cycls] ),
        .D(\gmiimode0.r[ifg_cycls][6]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/d [6]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[ifg_cycls][7] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[ifg_cycls] ),
        .D(\gmiimode0.r[ifg_cycls][7]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/d [7]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[ifg_cycls][8] 
       (.C(ethi),
        .CE(\m100.u0/ethc0/tx_rmii1.tx0/v[ifg_cycls] ),
        .D(\gmiimode0.r[ifg_cycls][8]_i_2_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/d [8]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[random][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][0] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][0] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][1] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random][2] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][1] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_1_in75_in ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random][3] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/p_1_in75_in ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_5_in ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random][4] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/p_5_in ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_7_in ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random][5] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/p_7_in ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][5] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random][6] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][5] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][6] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random][7] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][6] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][7] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random][8] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][7] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][8] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random][9] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[random_n_0_][8] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/p_0_in74_in ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt][0] 
       (.C(ethi),
        .CE(\gmiimode0.r[rcnt][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[rcnt] [0]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][0] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt][1] 
       (.C(ethi),
        .CE(\gmiimode0.r[rcnt][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[rcnt] [1]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][1] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt][2] 
       (.C(ethi),
        .CE(\gmiimode0.r[rcnt][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[rcnt] [2]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][2] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt][3] 
       (.C(ethi),
        .CE(\gmiimode0.r[rcnt][3]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[rcnt] [3]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rcnt_n_0_][3] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[read] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[read]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/txo[read] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[read_ack][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[read_ack] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[restart] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[restart]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/txo[restart] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt][0] 
       (.C(ethi),
        .CE(\gmiimode0.r[retry_cnt][4]_i_1_n_0 ),
        .D(\gmiimode0.r[retry_cnt][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][0] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt][1] 
       (.C(ethi),
        .CE(\gmiimode0.r[retry_cnt][4]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[retry_cnt] [1]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][1] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt][2] 
       (.C(ethi),
        .CE(\gmiimode0.r[retry_cnt][4]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[retry_cnt] [2]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][2] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt][3] 
       (.C(ethi),
        .CE(\gmiimode0.r[retry_cnt][4]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[retry_cnt] [3]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][3] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt][4] 
       (.C(ethi),
        .CE(\gmiimode0.r[retry_cnt][4]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[retry_cnt] [4]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[retry_cnt_n_0_][4] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[rmii_crc_en]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[rmii_crc_en]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count][0] 
       (.C(ethi),
        .CE(\gmiimode0.r[slot_count][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [0]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][0] ),
        .S(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count][1] 
       (.C(ethi),
        .CE(\gmiimode0.r[slot_count][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [1]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][1] ),
        .S(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count][2] 
       (.C(ethi),
        .CE(\gmiimode0.r[slot_count][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [2]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][2] ),
        .S(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count][3] 
       (.C(ethi),
        .CE(\gmiimode0.r[slot_count][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [3]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][3] ),
        .S(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count][4] 
       (.C(ethi),
        .CE(\gmiimode0.r[slot_count][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [4]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][4] ),
        .S(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count][5] 
       (.C(ethi),
        .CE(\gmiimode0.r[slot_count][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [5]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][5] ),
        .S(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count][6] 
       (.C(ethi),
        .CE(\gmiimode0.r[slot_count][6]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/v[slot_count] [6]),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[slot_count_n_0_][6] ),
        .S(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[speed][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\etho[speed] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/rin[speed] ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[speed][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/rin[speed] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/speed ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/r_reg[txstart_sync_n_0_] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [0]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[start][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[start]__0 [1]),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[status][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[status][0]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/txo[status] [0]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[status][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[status][1]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/txo[status] [1]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[switch]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[switch]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[transmitting] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[transmitting]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[transmitting]__0 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[tx_en] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[tx_en]_i_2_n_0 ),
        .Q(\etho[tx_en] ),
        .R(\gmiimode0.r[tx_en]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[txd][0] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r_reg[txd][0]_i_1_n_0 ),
        .Q(\^etho[txd] [0]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[txd][1] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r_reg[txd][1]_i_1_n_0 ),
        .Q(\^etho[txd] [1]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[txd][2] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/rin[txd_msb] [0]),
        .Q(\^etho[txd] [2]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[txd][3] 
       (.C(ethi),
        .CE(apbo),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/rin[txd_msb] [1]),
        .Q(\^etho[txd] [3]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero] 
       (.C(ethi),
        .CE(apbo),
        .D(\gmiimode0.r[zero]_i_1_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/gmiimode0.r_reg[zero]__1 ),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg[0] 
       (.C(ethi),
        .CE(apbo),
        .CLR(\r[ctrl][speed]_i_1_n_0 ),
        .D(apbo),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg_n_0_ ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg[1] 
       (.C(ethi),
        .CE(apbo),
        .CLR(\r[ctrl][speed]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg_n_0_ ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg_n_0_[1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg[2] 
       (.C(ethi),
        .CE(apbo),
        .CLR(\r[ctrl][speed]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg_n_0_[1] ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/p_1_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg[3] 
       (.C(ethi),
        .CE(apbo),
        .CLR(\r[ctrl][speed]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/p_1_in ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  (* equivalent_register_removal = "no" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg[4] 
       (.C(ethi),
        .CE(apbo),
        .CLR(\r[ctrl][speed]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/p_0_in ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/rstout0 
       (.I0(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/p_1_in ),
        .I1(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/r_reg_n_0_[4] ),
        .I2(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/p_0_in ),
        .O(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/rstout0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \m100.u0/ethc0/tx_rmii1.tx0/tx_rst/rstout_reg 
       (.C(ethi),
        .CE(apbo),
        .CLR(\r[ctrl][speed]_i_1_n_0 ),
        .D(\m100.u0/ethc0/tx_rmii1.tx0/tx_rst/rstout0_n_0 ),
        .Q(\m100.u0/ethc0/tx_rmii1.tx0/txrst ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[0] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[0]),
        .Q(\m100.u0/rxrdata [0]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[10] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[10]),
        .Q(\m100.u0/rxrdata [10]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[11] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[11]),
        .Q(\m100.u0/rxrdata [11]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[12] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[12]),
        .Q(\m100.u0/rxrdata [12]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[13] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[13]),
        .Q(\m100.u0/rxrdata [13]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[14] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[14]),
        .Q(\m100.u0/rxrdata [14]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[15] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[15]),
        .Q(\m100.u0/rxrdata [15]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[16] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[16]),
        .Q(\m100.u0/rxrdata [16]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[17] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[17]),
        .Q(\m100.u0/rxrdata [17]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[18] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[18]),
        .Q(\m100.u0/rxrdata [18]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[19] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[19]),
        .Q(\m100.u0/rxrdata [19]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[1] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[1]),
        .Q(\m100.u0/rxrdata [1]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[20] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[20]),
        .Q(\m100.u0/rxrdata [20]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[21] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[21]),
        .Q(\m100.u0/rxrdata [21]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[22] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[22]),
        .Q(\m100.u0/rxrdata [22]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[23] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[23]),
        .Q(\m100.u0/rxrdata [23]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[24] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[24]),
        .Q(\m100.u0/rxrdata [24]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[25] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[25]),
        .Q(\m100.u0/rxrdata [25]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[26] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[26]),
        .Q(\m100.u0/rxrdata [26]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[27] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[27]),
        .Q(\m100.u0/rxrdata [27]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[28] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[28]),
        .Q(\m100.u0/rxrdata [28]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[29] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[29]),
        .Q(\m100.u0/rxrdata [29]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[2] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[2]),
        .Q(\m100.u0/rxrdata [2]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[30] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[30]),
        .Q(\m100.u0/rxrdata [30]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[31] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[31]),
        .Q(\m100.u0/rxrdata [31]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[3] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[3]),
        .Q(\m100.u0/rxrdata [3]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[4] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[4]),
        .Q(\m100.u0/rxrdata [4]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[5] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[5]),
        .Q(\m100.u0/rxrdata [5]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[6] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[6]),
        .Q(\m100.u0/rxrdata [6]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[7] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[7]),
        .Q(\m100.u0/rxrdata [7]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[8] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[8]),
        .Q(\m100.u0/rxrdata [8]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/oneclk.q_reg[9] 
       (.C(clk),
        .CE(apbo),
        .D(p_0_out[9]),
        .Q(\m100.u0/rxrdata [9]),
        .R(etho));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/rfd_reg_0_3_0_5 
       (.ADDRA({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRB({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRC({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRD({etho,etho,etho,\m100.u0/rxwaddress }),
        .DIA(\m100.u0/rxwdata [1:0]),
        .DIB(\m100.u0/rxwdata [3:2]),
        .DIC(\m100.u0/rxwdata [5:4]),
        .DID({etho,etho}),
        .DOA(p_0_out[1:0]),
        .DOB(p_0_out[3:2]),
        .DOC(p_0_out[5:4]),
        .WCLK(clk),
        .WE(\m100.u0/rxwrite ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/rfd_reg_0_3_12_17 
       (.ADDRA({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRB({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRC({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRD({etho,etho,etho,\m100.u0/rxwaddress }),
        .DIA(\m100.u0/rxwdata [13:12]),
        .DIB(\m100.u0/rxwdata [15:14]),
        .DIC(\m100.u0/rxwdata [17:16]),
        .DID({etho,etho}),
        .DOA(p_0_out[13:12]),
        .DOB(p_0_out[15:14]),
        .DOC(p_0_out[17:16]),
        .WCLK(clk),
        .WE(\m100.u0/rxwrite ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/rfd_reg_0_3_18_23 
       (.ADDRA({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRB({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRC({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRD({etho,etho,etho,\m100.u0/rxwaddress }),
        .DIA(\m100.u0/rxwdata [19:18]),
        .DIB(\m100.u0/rxwdata [21:20]),
        .DIC(\m100.u0/rxwdata [23:22]),
        .DID({etho,etho}),
        .DOA(p_0_out[19:18]),
        .DOB(p_0_out[21:20]),
        .DOC(p_0_out[23:22]),
        .WCLK(clk),
        .WE(\m100.u0/rxwrite ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/rfd_reg_0_3_24_29 
       (.ADDRA({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRB({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRC({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRD({etho,etho,etho,\m100.u0/rxwaddress }),
        .DIA(\m100.u0/rxwdata [25:24]),
        .DIB(\m100.u0/rxwdata [27:26]),
        .DIC(\m100.u0/rxwdata [29:28]),
        .DID({etho,etho}),
        .DOA(p_0_out[25:24]),
        .DOB(p_0_out[27:26]),
        .DOC(p_0_out[29:28]),
        .WCLK(clk),
        .WE(\m100.u0/rxwrite ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/rfd_reg_0_3_30_31 
       (.ADDRA({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRB({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRC({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRD({etho,etho,etho,\m100.u0/rxwaddress }),
        .DIA(\m100.u0/rxwdata [31:30]),
        .DIB({etho,etho}),
        .DIC({etho,etho}),
        .DID({etho,etho}),
        .DOA(p_0_out[31:30]),
        .WCLK(clk),
        .WE(\m100.u0/rxwrite ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "" *) 
  RAM32M #(
    .INIT_A(64'h0000000000000000),
    .INIT_B(64'h0000000000000000),
    .INIT_C(64'h0000000000000000),
    .INIT_D(64'h0000000000000000),
    .IS_WCLK_INVERTED(1'b0)) 
    \m100.u0/nft.rx_fifo0/xc2v.x0/a0.x0/rfd_reg_0_3_6_11 
       (.ADDRA({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRB({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRC({etho,etho,etho,\m100.u0/rxraddress }),
        .ADDRD({etho,etho,etho,\m100.u0/rxwaddress }),
        .DIA(\m100.u0/rxwdata [7:6]),
        .DIB(\m100.u0/rxwdata [9:8]),
        .DIC(\m100.u0/rxwdata [11:10]),
        .DID({etho,etho}),
        .DOA(p_0_out[7:6]),
        .DOB(p_0_out[9:8]),
        .DOC(p_0_out[11:10]),
        .WCLK(clk),
        .WE(\m100.u0/rxwrite ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* PWROPT_WRITE_MODE_CHANGE_A = "WRITE_FIRST:NO_CHANGE_1" *) 
  (* XILINX_LEGACY_PRIM = "RAMB16_S36_S36" *) 
  (* XILINX_TRANSFORM_PINMAP = "ADDRA[0]:ADDRARDADDR[0],ADDRARDADDR[10] ADDRA[1]:ADDRARDADDR[1],ADDRARDADDR[11] ADDRA[2]:ADDRARDADDR[2],ADDRARDADDR[12] ADDRA[3]:ADDRARDADDR[3],ADDRARDADDR[13] ADDRA[4]:ADDRARDADDR[4],ADDRARDADDR[9] ADDRB[0]:ADDRBWRADDR[0],ADDRBWRADDR[10] ADDRB[1]:ADDRBWRADDR[1],ADDRBWRADDR[11] ADDRB[2]:ADDRBWRADDR[2],ADDRBWRADDR[12] ADDRB[3]:ADDRBWRADDR[3],ADDRBWRADDR[13] ADDRB[4]:ADDRBWRADDR[4],ADDRBWRADDR[9] WEA:WEA[3],WEA[2],WEA[1],WEA[0] WEB:WEBWE[3],WEBWE[2],WEBWE[1],WEBWE[0] ADDRA[14]:ADDRARDADDR[14] ADDRA[5]:ADDRARDADDR[5] ADDRA[6]:ADDRARDADDR[6] ADDRA[7]:ADDRARDADDR[7] ADDRA[8]:ADDRARDADDR[8] ADDRB[14]:ADDRBWRADDR[14] ADDRB[5]:ADDRBWRADDR[5] ADDRB[6]:ADDRBWRADDR[6] ADDRB[7]:ADDRBWRADDR[7] ADDRB[8]:ADDRBWRADDR[8] CLKA:CLKARDCLK CLKB:CLKBWRCLK DIA[0]:DIADI[0] DIA[10]:DIADI[10] DIA[11]:DIADI[11] DIA[12]:DIADI[12] DIA[13]:DIADI[13] DIA[14]:DIADI[14] DIA[15]:DIADI[15] DIA[16]:DIADI[16] DIA[17]:DIADI[17] DIA[18]:DIADI[18] DIA[19]:DIADI[19] DIA[1]:DIADI[1] DIA[20]:DIADI[20] DIA[21]:DIADI[21] DIA[22]:DIADI[22] DIA[23]:DIADI[23] DIA[24]:DIADI[24] DIA[25]:DIADI[25] DIA[26]:DIADI[26] DIA[27]:DIADI[27] DIA[28]:DIADI[28] DIA[29]:DIADI[29] DIA[2]:DIADI[2] DIA[30]:DIADI[30] DIA[31]:DIADI[31] DIA[3]:DIADI[3] DIA[4]:DIADI[4] DIA[5]:DIADI[5] DIA[6]:DIADI[6] DIA[7]:DIADI[7] DIA[8]:DIADI[8] DIA[9]:DIADI[9] DIB[0]:DIBDI[0] DIB[10]:DIBDI[10] DIB[11]:DIBDI[11] DIB[12]:DIBDI[12] DIB[13]:DIBDI[13] DIB[14]:DIBDI[14] DIB[15]:DIBDI[15] DIB[16]:DIBDI[16] DIB[17]:DIBDI[17] DIB[18]:DIBDI[18] DIB[19]:DIBDI[19] DIB[1]:DIBDI[1] DIB[20]:DIBDI[20] DIB[21]:DIBDI[21] DIB[22]:DIBDI[22] DIB[23]:DIBDI[23] DIB[24]:DIBDI[24] DIB[25]:DIBDI[25] DIB[26]:DIBDI[26] DIB[27]:DIBDI[27] DIB[28]:DIBDI[28] DIB[29]:DIBDI[29] DIB[2]:DIBDI[2] DIB[30]:DIBDI[30] DIB[31]:DIBDI[31] DIB[3]:DIBDI[3] DIB[4]:DIBDI[4] DIB[5]:DIBDI[5] DIB[6]:DIBDI[6] DIB[7]:DIBDI[7] DIB[8]:DIBDI[8] DIB[9]:DIBDI[9] DIPA[0]:DIPADIP[0] DIPA[1]:DIPADIP[1] DIPA[2]:DIPADIP[2] DIPA[3]:DIPADIP[3] DIPB[0]:DIPBDIP[0] DIPB[1]:DIPBDIP[1] DIPB[2]:DIPBDIP[2] DIPB[3]:DIPBDIP[3] DOA[0]:DOADO[0] DOA[10]:DOADO[10] DOA[11]:DOADO[11] DOA[12]:DOADO[12] DOA[13]:DOADO[13] DOA[14]:DOADO[14] DOA[15]:DOADO[15] DOA[16]:DOADO[16] DOA[17]:DOADO[17] DOA[18]:DOADO[18] DOA[19]:DOADO[19] DOA[1]:DOADO[1] DOA[20]:DOADO[20] DOA[21]:DOADO[21] DOA[22]:DOADO[22] DOA[23]:DOADO[23] DOA[24]:DOADO[24] DOA[25]:DOADO[25] DOA[26]:DOADO[26] DOA[27]:DOADO[27] DOA[28]:DOADO[28] DOA[29]:DOADO[29] DOA[2]:DOADO[2] DOA[30]:DOADO[30] DOA[31]:DOADO[31] DOA[3]:DOADO[3] DOA[4]:DOADO[4] DOA[5]:DOADO[5] DOA[6]:DOADO[6] DOA[7]:DOADO[7] DOA[8]:DOADO[8] DOA[9]:DOADO[9] DOB[0]:DOBDO[0] DOB[10]:DOBDO[10] DOB[11]:DOBDO[11] DOB[12]:DOBDO[12] DOB[13]:DOBDO[13] DOB[14]:DOBDO[14] DOB[15]:DOBDO[15] DOB[16]:DOBDO[16] DOB[17]:DOBDO[17] DOB[18]:DOBDO[18] DOB[19]:DOBDO[19] DOB[1]:DOBDO[1] DOB[20]:DOBDO[20] DOB[21]:DOBDO[21] DOB[22]:DOBDO[22] DOB[23]:DOBDO[23] DOB[24]:DOBDO[24] DOB[25]:DOBDO[25] DOB[26]:DOBDO[26] DOB[27]:DOBDO[27] DOB[28]:DOBDO[28] DOB[29]:DOBDO[29] DOB[2]:DOBDO[2] DOB[30]:DOBDO[30] DOB[31]:DOBDO[31] DOB[3]:DOBDO[3] DOB[4]:DOBDO[4] DOB[5]:DOBDO[5] DOB[6]:DOBDO[6] DOB[7]:DOBDO[7] DOB[8]:DOBDO[8] DOB[9]:DOBDO[9] DOPA[0]:DOPADOP[0] DOPA[1]:DOPADOP[1] DOPA[2]:DOPADOP[2] DOPA[3]:DOPADOP[3] DOPB[0]:DOPBDOP[0] DOPB[1]:DOPBDOP[1] DOPB[2]:DOPBDOP[2] DOPB[3]:DOPBDOP[3] ENA:ENARDEN ENB:ENBWREN REGCEA:REGCEAREGCE SSRA:RSTRAMARSTRAM SSRB:RSTRAMB" *) 
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
    .READ_WIDTH_A(36),
    .READ_WIDTH_B(36),
    .RSTREG_PRIORITY_A("REGCE"),
    .RSTREG_PRIORITY_B("REGCE"),
    .SIM_COLLISION_CHECK("GENERATE_X_ONLY"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("NO_CHANGE"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(36),
    .WRITE_WIDTH_B(36)) 
    \m100.u0/nft.tx_fifo0/xc2v.x0/a6.x0/a9.x[0].r0 
       (.ADDRARDADDR({VCC_2,GND_2,etho,etho,\m100.u0/txwaddress ,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .ADDRBWRADDR({VCC_2,GND_2,etho,etho,\m100.u0/txraddress ,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI(\m100.u0/txwdata ),
        .DIBDI({etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho,etho}),
        .DIPADIP({etho,etho,etho,etho}),
        .DIPBDIP({etho,etho,etho,etho}),
        .DOBDO(\m100.u0/txrdata ),
        .ENARDEN(\m100.u0/txwrite ),
        .ENBWREN(\m100.u0/txrenable ),
        .REGCEAREGCE(GND_2),
        .REGCEB(GND_2),
        .RSTRAMARSTRAM(etho),
        .RSTRAMB(etho),
        .RSTREGARSTREG(GND_2),
        .RSTREGB(GND_2),
        .WEA({\m100.u0/txwrite ,\m100.u0/txwrite ,\m100.u0/txwrite ,\m100.u0/txwrite }),
        .WEBWE({GND_2,GND_2,GND_2,GND_2,etho,etho,etho,etho}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFF00)) 
    \m100.u0/r[addrdone]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\m100.u0/ethc0/v ),
        .I4(\m100.u0/ethc0/r_reg[addrdone]__0 ),
        .O(\m100.u0/r ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFF00)) 
    \m100.u0/r[addrok]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\m100.u0/ethc0/v[addrok]62_out ),
        .I4(\m100.u0/ethc0/r_reg[addrok_n_0_] ),
        .O(\m100.u0/r[addrok]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7533753045004500)) 
    \m100.u0/r[bcast]_i_1 
       (.I0(\r[msbgood]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/v[addrok] ),
        .I2(\r[bcast]_i_3_n_0 ),
        .I3(\r[bcast]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[bcast_n_0_] ),
        .O(\m100.u0/r[bcast]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \m100.u0/r[ctrl][edcldis]_i_1 
       (.I0(\apbi[pwdata] [14]),
        .I1(\m100.u0/ethc0/v[ctrl][txen] ),
        .I2(\m100.u0/ethc0/p_6_in [14]),
        .O(\m100.u0/r[ctrl][edcldis]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111F0FF1111F000)) 
    \m100.u0/r[ctrl][full_duplex]_i_1 
       (.I0(\r[ctrl][full_duplex]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I2(\apbi[pwdata] [4]),
        .I3(\m100.u0/ethc0/v[ctrl][txen] ),
        .I4(\r[ctrl][full_duplex]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/p_6_in [4]),
        .O(\m100.u0/r[ctrl][full_duplex]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \m100.u0/r[ctrl][rxen]_i_1 
       (.I0(\m100.u0/ethc0/v[ctrl][rxen] ),
        .I1(\r[ctrl][rxen]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/p_6_in [1]),
        .O(\m100.u0/r[ctrl][rxen]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAEFEFEFAAE0E0E0)) 
    \m100.u0/r[ctrl][speed]_i_2 
       (.I0(\r[ctrl][speed]_i_3_n_0 ),
        .I1(\apbi[pwdata] [7]),
        .I2(\m100.u0/ethc0/v[ctrl][txen] ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\etho[speed] ),
        .O(\m100.u0/r[ctrl][speed]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8888F0FF8888F000)) 
    \m100.u0/r[ctrl][txen]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\ahbmi[hrdata] [11]),
        .I2(\apbi[pwdata] [0]),
        .I3(\m100.u0/ethc0/v[ctrl][txen] ),
        .I4(\r[ctrl][txen]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/p_6_in [0]),
        .O(\m100.u0/r[ctrl][txen]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF7EFEFFFF0000)) 
    \m100.u0/r[ctrlpkt]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I3(\m100.u0/ethc0/v[ctrlpkt]69_out ),
        .I4(\m100.u0/ethc0/v[ctrlpkt]68_out ),
        .I5(\m100.u0/ethc0/r_reg[ctrlpkt]__0 ),
        .O(\m100.u0/r[ctrlpkt]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \m100.u0/r[disableduplex]_i_1 
       (.I0(\apbi[pwdata] [12]),
        .I1(\m100.u0/ethc0/v[ctrl][txen] ),
        .I2(\m100.u0/ethc0/p_6_in [12]),
        .O(\m100.u0/r[disableduplex]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h808080FF80808000)) 
    \m100.u0/r[edclactive]_i_1 
       (.I0(\m100.u0/ethc0/v[edclactive]58_out ),
        .I1(\r[rcntm][2]_i_2_n_0 ),
        .I2(\r[edclactive]_i_3_n_0 ),
        .I3(\r[edclactive]_i_4_n_0 ),
        .I4(\r[edclactive]_i_5_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[edclactive_n_0_] ),
        .O(\m100.u0/r[edclactive]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0440FFFF04400000)) 
    \m100.u0/r[edclbcast]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I4(\r[edclbcast]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[edclbcast]__0 ),
        .O(\m100.u0/r[edclbcast]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFE00000002)) 
    \m100.u0/r[erenable]_i_1 
       (.I0(\m100.u0/ethc0/v[tmsto][req]1149_out ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\m100.u0/erenable ),
        .O(\m100.u0/r[erenable]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFB0000000B)) 
    \m100.u0/r[erxidle]_i_1 
       (.I0(\m100.u0/ethc0/p_6_in [14]),
        .I1(\r[erxidle]_i_2_n_0 ),
        .I2(\r[erxidle]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I5(\m100.u0/ethc0/r_reg[erxidle]__0 ),
        .O(\m100.u0/r[erxidle]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFFFEB28000028)) 
    \m100.u0/r[gotframe]_i_1 
       (.I0(\m100.u0/ethc0/rxo[gotframe] ),
        .I1(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rxdone] ),
        .I3(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I4(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I5(\m100.u0/ethc0/r_reg[gotframe_n_0_] ),
        .O(\m100.u0/r[gotframe]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000CEEE)) 
    \m100.u0/r[init_busy]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[init_busy_n_0_] ),
        .I1(\r[mdio_ctrl][data][15]_i_2_n_0 ),
        .I2(\r[init_busy]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I4(\m100.u0/ethc0/v[mdio_ctrl][write]113_out ),
        .O(\m100.u0/r[init_busy]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEFFCECECECC)) 
    \m100.u0/r[mdio_ctrl][busy]_i_1 
       (.I0(\r[mdio_ctrl][busy]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][15]_i_2_n_0 ),
        .I2(\r[mdio_ctrl][busy]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/v[mdio_ctrl][busy] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][busy]__0 ),
        .O(\m100.u0/r[mdio_ctrl][busy]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F004FFF40004000)) 
    \m100.u0/r[mdio_ctrl][linkfail]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I1(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I2(\r[mdio_ctrl][linkfail]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I4(\r[mdio_ctrl][linkfail]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][linkfail_n_0_] ),
        .O(\m100.u0/r[mdio_ctrl][linkfail]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFABFBFFFFA808)) 
    \m100.u0/r[mdio_ctrl][read]_i_1 
       (.I0(\r[mdio_ctrl][read]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I3(\r[mdio_ctrl][write]_i_4_n_0 ),
        .I4(\r[mdio_ctrl][read]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .O(\m100.u0/r[mdio_ctrl][read]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFABFBFFFFA808)) 
    \m100.u0/r[mdio_ctrl][write]_i_1 
       (.I0(\r_reg[mdio_ctrl][write]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][write]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I3(\r[mdio_ctrl][write]_i_4_n_0 ),
        .I4(\r[mdio_ctrl][write]_i_5_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][write]__0 ),
        .O(\m100.u0/r[mdio_ctrl][write]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE01)) 
    \m100.u0/r[mdioclk]_i_2 
       (.I0(\r[mdioclk]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/d [4]),
        .I2(\m100.u0/ethc0/d [5]),
        .I3(\etho[mdc] ),
        .O(\m100.u0/r[mdioclk]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \m100.u0/r[mdioen]_i_1 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][write]1 ),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/v[mdioen] ),
        .I5(\etho[mdio_oe] ),
        .O(\m100.u0/r[mdioen]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \m100.u0/r[mdioo]_i_1 
       (.I0(\r[mdioo]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/v[mdioo] ),
        .I2(\etho[mdio_o] ),
        .O(\m100.u0/r[mdioo]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFEFE00FF0000)) 
    \m100.u0/r[msbgood]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\r[msbgood]_i_2_n_0 ),
        .I4(\r_reg[msbgood]_i_3_n_1 ),
        .I5(\m100.u0/ethc0/r_reg[msbgood_n_0_] ),
        .O(\m100.u0/r[msbgood]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFBFF0800)) 
    \m100.u0/r[phywr]_i_1 
       (.I0(\r[phywr]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/v[phywr] ),
        .I2(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .O(\m100.u0/r[phywr]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \m100.u0/r[rmsto][write]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[rmsto][write_n_0_] ),
        .O(\m100.u0/r[rmsto][write]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF02000000)) 
    \m100.u0/r[rstaneg]_i_1 
       (.I0(\r[rstaneg]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I4(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I5(\m100.u0/ethc0/r_reg[rstaneg_n_0_] ),
        .O(\m100.u0/r[rstaneg]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAA8AAAA)) 
    \m100.u0/r[rstphy]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rstphy]__0 ),
        .I1(\m100.u0/ethc0/r_reg[init_busy_n_0_] ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][linkfail_n_0_] ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .O(\m100.u0/r[rstphy]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \m100.u0/r[rxden]_i_1 
       (.I0(\ahbmi[hrdata] [11]),
        .I1(\m100.u0/ethc0/v[rxwrap] ),
        .I2(\m100.u0/ethc0/r_reg[rxden]__0 ),
        .O(\m100.u0/r[rxden]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF690)) 
    \m100.u0/r[rxdoneack]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I2(\m100.u0/ethc0/r_reg[rxdone] ),
        .I3(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\m100.u0/r[rxdoneack]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \m100.u0/r[rxirq]_i_1 
       (.I0(\ahbmi[hrdata] [13]),
        .I1(\m100.u0/ethc0/v[rxwrap] ),
        .I2(\m100.u0/ethc0/r_reg[rxirq]__0 ),
        .O(\m100.u0/r[rxirq]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \m100.u0/r[rxwrap]_i_1 
       (.I0(\ahbmi[hrdata] [12]),
        .I1(\m100.u0/ethc0/v[rxwrap] ),
        .I2(\m100.u0/ethc0/r_reg[rxwrap_n_0_] ),
        .O(\m100.u0/r[rxwrap]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4000FFFF40004000)) 
    \m100.u0/r[status][invaddr]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\r[status][invaddr]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\m100.u0/ethc0/v[status][invaddr]45_out ),
        .I5(\m100.u0/ethc0/r_reg[status][invaddr_n_0_] ),
        .O(\m100.u0/r[status][invaddr]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4000FFFF40004000)) 
    \m100.u0/r[status][rx_err]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\m100.u0/ethc0/v[status][rx_err]15_out ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\m100.u0/ethc0/v[status][rx_err]18_out ),
        .I5(\m100.u0/ethc0/r_reg[status][rx_err_n_0_] ),
        .O(\m100.u0/r[status][rx_err]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4000FFFF40004000)) 
    \m100.u0/r[status][rx_int]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\r[status][rx_int]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\m100.u0/ethc0/v[status][rx_int]26_out ),
        .I5(\m100.u0/ethc0/r_reg[status][rx_int_n_0_] ),
        .O(\m100.u0/r[status][rx_int]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4088FFFF40884088)) 
    \m100.u0/r[status][rxahberr]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/rmsti ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/v[status][rxahberr]32_out ),
        .I5(\m100.u0/ethc0/r_reg[status][rxahberr_n_0_] ),
        .O(\m100.u0/r[status][rxahberr]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4000FFFF40004000)) 
    \m100.u0/r[status][toosmall]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/v[status][toosmall]39_out ),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\m100.u0/ethc0/v[status][toosmall]42_out ),
        .I5(\m100.u0/ethc0/r_reg[status][toosmall_n_0_] ),
        .O(\m100.u0/r[status][toosmall]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFE0FFFFE0E0E0E0)) 
    \m100.u0/r[status][tx_err]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txstatus_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txstatus_n_0_][0] ),
        .I2(\r[txdsel][9]_i_3_n_0 ),
        .I3(\r[status][tx_int]_i_2_n_0 ),
        .I4(\apbi[pwdata] [1]),
        .I5(\m100.u0/ethc0/r_reg[status][tx_err_n_0_] ),
        .O(\m100.u0/r[status][tx_err]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF10FFFF10101010)) 
    \m100.u0/r[status][tx_int]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txstatus_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txstatus_n_0_][0] ),
        .I2(\r[txdsel][9]_i_3_n_0 ),
        .I3(\r[status][tx_int]_i_2_n_0 ),
        .I4(\apbi[pwdata] [3]),
        .I5(\m100.u0/ethc0/r_reg[status][tx_int_n_0_] ),
        .O(\m100.u0/r[status][tx_int]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFFAAAAAAAA)) 
    \m100.u0/r[status][txahberr]_i_1 
       (.I0(\m100.u0/ethc0/rin[status][txahberr] ),
        .I1(\apbi[paddr] [5]),
        .I2(\apbi[paddr] [3]),
        .I3(\r[status][txahberr]_i_2_n_0 ),
        .I4(\apbi[pwdata] [5]),
        .I5(\m100.u0/ethc0/r_reg[status][txahberr_n_0_] ),
        .O(\m100.u0/r[status][txahberr]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F20)) 
    \m100.u0/r[tarp]_i_1 
       (.I0(\r[tarp]_i_2_n_0 ),
        .I1(\r[tarp]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[tarp]0 ),
        .I3(\m100.u0/ethc0/r_reg[tarp]__0 ),
        .O(\m100.u0/r[tarp]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEFE01000000)) 
    \m100.u0/r[tedcl]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\r[tedcl]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I5(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .O(\m100.u0/r[tedcl]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F8F8FFF8F8F8F00)) 
    \m100.u0/r[tmsto][write]_i_1 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\r[tmsto][write]_i_3_n_0 ),
        .I3(\r[tmsto][write]_i_4_n_0 ),
        .I4(\r[tmsto][write]_i_5_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[tmsto][write_n_0_] ),
        .O(\m100.u0/r[tmsto][write]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \m100.u0/r[tnak]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[tnak]__0 ),
        .I1(\r[txlength][10]_i_5_n_0 ),
        .I2(\m100.u0/erdata [10]),
        .O(\m100.u0/r[tnak]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \m100.u0/r[txden]_i_1 
       (.I0(\ahbmi[hrdata] [11]),
        .I1(\m100.u0/ethc0/v[txirq] ),
        .I2(\m100.u0/ethc0/r_reg[txden]__0 ),
        .O(\m100.u0/r[txden]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \m100.u0/r[txirq]_i_1 
       (.I0(\ahbmi[hrdata] [13]),
        .I1(\m100.u0/ethc0/v[txirq] ),
        .I2(\m100.u0/ethc0/r_reg[txirq]__0 ),
        .O(\m100.u0/r[txirq]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h808080FF80808000)) 
    \m100.u0/r[txirqgen]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/p_6_in [2]),
        .I2(\m100.u0/ethc0/r_reg[txirq]__0 ),
        .I3(\r[txdsel][9]_i_3_n_0 ),
        .I4(\apbo[pirq][12]_INST_0_i_2_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txirqgen_n_0_] ),
        .O(\m100.u0/r[txirqgen]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFF0000000004)) 
    \m100.u0/r[txstart]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r[txstart]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txstart]__0 ),
        .O(\m100.u0/r[txstart]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDDDDDD02222222F)) 
    \m100.u0/r[txstart_sync]_i_1 
       (.I0(\r[txstart_sync]_i_2_n_0 ),
        .I1(\r[txstart_sync]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\r[txstart_sync]_i_4_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txstart_sync_n_0_] ),
        .O(\m100.u0/r[txstart_sync]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \m100.u0/r[txwrap]_i_1 
       (.I0(\ahbmi[hrdata] [12]),
        .I1(\m100.u0/ethc0/v[txirq] ),
        .I2(\m100.u0/ethc0/r_reg[txwrap_n_0_] ),
        .O(\m100.u0/r[txwrap]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBAAB8AA8)) 
    \m100.u0/r[writeok]_i_1 
       (.I0(\r[writeok]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/v[rxlength] ),
        .I2(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I4(\m100.u0/ethc0/r_reg[writeok_n_0_] ),
        .O(\m100.u0/r[writeok]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD5D755FF2A28AA00)) 
    \r[abufs][0]_i_1 
       (.I0(\r[abufs][0]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\r[abufs][0]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\r[abufs][2]_i_6_n_0 ),
        .O(r));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEEEEFEFFFE)) 
    \r[abufs][0]_i_2 
       (.I0(\r[abufs][2]_i_15_n_0 ),
        .I1(\r[abufs][0]_i_4_n_0 ),
        .I2(\r[abufs][0]_i_3_n_0 ),
        .I3(\r[rpnt][1]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/r_reg ),
        .I5(\r[erxidle]_i_3_n_0 ),
        .O(\r[abufs][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAA6AAAAAA)) 
    \r[abufs][0]_i_3 
       (.I0(\m100.u0/ethc0/r_reg ),
        .I1(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[abufs][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[abufs][0]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\r[abufs][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h9A)) 
    \r[abufs][1]_i_1 
       (.I0(\m100.u0/ethc0/v[abufs] [1]),
        .I1(\m100.u0/ethc0/v[abufs] [0]),
        .I2(\r[abufs][2]_i_6_n_0 ),
        .O(\r[abufs][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE0E0E0E0E01FE0E0)) 
    \r[abufs][2]_i_1 
       (.I0(\r[abufs][2]_i_2_n_0 ),
        .I1(\r[abufs][2]_i_3_n_0 ),
        .I2(\r[abufs][2]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/v[abufs] [1]),
        .I4(\r[abufs][2]_i_6_n_0 ),
        .I5(\m100.u0/ethc0/v[abufs] [0]),
        .O(\r[abufs][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r[abufs][2]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[abufs][2]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF708)) 
    \r[abufs][2]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I1(\m100.u0/ethc0/rin[status][txahberr] ),
        .I2(\m100.u0/ethc0/r_reg ),
        .I3(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .O(\r[abufs][2]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000A8ABABA8)) 
    \r[abufs][2]_i_12 
       (.I0(\r[abufs][2]_i_11_n_0 ),
        .I1(\r[abufs][2]_i_16_n_0 ),
        .I2(\r[rxstatus][4]_i_1_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg ),
        .I5(\r[erxidle]_i_3_n_0 ),
        .O(\r[abufs][2]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA8BB80000)) 
    \r[abufs][2]_i_13 
       (.I0(\r[abufs][2]_i_11_n_0 ),
        .I1(\r[erxidle]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg ),
        .I3(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\r[abufs][2]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000A8AB)) 
    \r[abufs][2]_i_14 
       (.I0(\r[abufs][0]_i_3_n_0 ),
        .I1(\r[abufs][2]_i_16_n_0 ),
        .I2(\r[rxstatus][4]_i_1_n_0 ),
        .I3(\m100.u0/ethc0/r_reg ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\r[abufs][2]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA28EB0000)) 
    \r[abufs][2]_i_15 
       (.I0(\r[abufs][0]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\r[abufs][2]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    \r[abufs][2]_i_16 
       (.I0(\r[rxstatus][1]_i_1_n_0 ),
        .I1(\r[rxstatus][3]_i_1_n_0 ),
        .I2(\r[rxstatus][2]_i_1_n_0 ),
        .I3(\m100.u0/ethc0/rxo[gotframe] ),
        .I4(\m100.u0/ethc0/rxo[status] [0]),
        .I5(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[abufs][2]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAEB280000)) 
    \r[abufs][2]_i_2 
       (.I0(\r[abufs][2]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\r[abufs][2]_i_9_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\r[abufs][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4540FFFFFFFFFFFF)) 
    \r[abufs][2]_i_3 
       (.I0(\r[erxidle]_i_3_n_0 ),
        .I1(\r[abufs][2]_i_9_n_0 ),
        .I2(\r[rpnt][1]_i_3_n_0 ),
        .I3(\r[abufs][2]_i_8_n_0 ),
        .I4(\r[abufs][2]_i_10_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\r[abufs][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h76F0)) 
    \r[abufs][2]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\r[abufs][2]_i_8_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\r[abufs][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0FFAAAAA0CCAAAAA)) 
    \r[abufs][2]_i_5 
       (.I0(\r[abufs][2]_i_11_n_0 ),
        .I1(\r[abufs][2]_i_12_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\r[abufs][2]_i_13_n_0 ),
        .O(\m100.u0/ethc0/v[abufs] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000002800000000)) 
    \r[abufs][2]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[abufs][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0FFAAAAA0CCAAAAA)) 
    \r[abufs][2]_i_7 
       (.I0(\r[abufs][0]_i_3_n_0 ),
        .I1(\r[abufs][2]_i_14_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\r[abufs][2]_i_15_n_0 ),
        .O(\m100.u0/ethc0/v[abufs] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA9AAAAAA)) 
    \r[abufs][2]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[abufs_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg ),
        .I2(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .I3(\m100.u0/ethc0/rin[status][txahberr] ),
        .I4(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .O(\r[abufs][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    \r[abufs][2]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[abufs_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg ),
        .O(\r[abufs][2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \r[addrdone]_i_2 
       (.I0(\r[addrdone]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .O(\m100.u0/ethc0/v ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \r[addrdone]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .I3(\r[msbgood]_i_9_n_0 ),
        .O(\r[addrdone]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[addrok]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [21]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [19]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][4] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [20]),
        .O(\r[addrok]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[addrok]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [17]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [18]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[checkdata]__0 [16]),
        .I5(\m100.u0/ethc0/r_reg[mac_addr_n_0_][0] ),
        .O(\r[addrok]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02300200)) 
    \r[addrok]_i_2 
       (.I0(\m100.u0/ethc0/p_6_in [5]),
        .I1(\r[msbgood]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I4(\r[addrok]_i_3_n_0 ),
        .O(\m100.u0/ethc0/v[addrok]62_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \r[addrok]_i_3 
       (.I0(r_reg[1]),
        .I1(\m100.u0/ethc0/r_reg[msbgood_n_0_] ),
        .I2(\r[bcast]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[bcast_n_0_] ),
        .O(\r[addrok]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r[addrok]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][15] ),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [31]),
        .O(\r[addrok]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[addrok]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [29]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][13] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [28]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][12] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][14] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [30]),
        .O(\r[addrok]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[addrok]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [25]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][9] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [26]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][10] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][11] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [27]),
        .O(\r[addrok]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[addrok]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [22]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][6] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [23]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][7] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][8] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [24]),
        .O(\r[addrok]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \r[applength][0]_i_1 
       (.I0(\m100.u0/rxwdata [7]),
        .I1(\m100.u0/ethc0/v[nak]1 ),
        .I2(\m100.u0/rxwdata [17]),
        .O(\r[applength][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \r[applength][1]_i_1 
       (.I0(\m100.u0/rxwdata [8]),
        .I1(\m100.u0/ethc0/v[nak]1 ),
        .I2(\m100.u0/rxwdata [17]),
        .O(\r[applength][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \r[applength][2]_i_1 
       (.I0(\m100.u0/rxwdata [9]),
        .I1(\m100.u0/rxwdata [17]),
        .I2(\m100.u0/ethc0/v[nak]1 ),
        .O(\r[applength][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \r[applength][3]_i_1 
       (.I0(\m100.u0/rxwdata [10]),
        .I1(\m100.u0/rxwdata [17]),
        .I2(\m100.u0/ethc0/v[nak]1 ),
        .O(\r[applength][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \r[applength][4]_i_1 
       (.I0(\m100.u0/rxwdata [11]),
        .I1(\m100.u0/ethc0/v[nak]1 ),
        .I2(\m100.u0/rxwdata [17]),
        .O(\r[applength][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \r[applength][5]_i_1 
       (.I0(\m100.u0/rxwdata [12]),
        .I1(\m100.u0/ethc0/v[nak]1 ),
        .I2(\m100.u0/rxwdata [17]),
        .O(\r[applength][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \r[applength][6]_i_1 
       (.I0(\m100.u0/rxwdata [13]),
        .I1(\m100.u0/ethc0/v[nak]1 ),
        .I2(\m100.u0/rxwdata [17]),
        .O(\r[applength][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \r[applength][7]_i_1 
       (.I0(\m100.u0/rxwdata [14]),
        .I1(\m100.u0/ethc0/v[nak]1 ),
        .I2(\m100.u0/rxwdata [17]),
        .O(\r[applength][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \r[applength][8]_i_1 
       (.I0(\m100.u0/rxwdata [15]),
        .I1(\m100.u0/ethc0/v[nak]1 ),
        .I2(\m100.u0/rxwdata [17]),
        .O(\r[applength][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \r[applength][9]_i_1 
       (.I0(\m100.u0/rxwdata [16]),
        .I1(\m100.u0/ethc0/v[nak]1 ),
        .I2(\m100.u0/rxwdata [17]),
        .O(\r[applength][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00C0A0A0)) 
    \r[ba]_i_1 
       (.I0(\m100.u0/ethc0/ahb0/r_reg ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bg]__0 ),
        .I2(rst),
        .I3(\r[ba]_i_2_n_0 ),
        .I4(\ahbmi[hready] ),
        .O(\r[ba]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEEEF)) 
    \r[ba]_i_2 
       (.I0(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[error]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .O(\r[ba]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[bb]_i_1 
       (.I0(\m100.u0/ethc0/ahb0/v ),
        .I1(\ahbmi[hready] ),
        .I2(\m100.u0/ethc0/ahb0/r_reg[bb]__0 ),
        .O(\r[bb]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF800080008000)) 
    \r[bb]_i_2 
       (.I0(\m100.u0/ethc0/ahb0/nbo ),
        .I1(\m100.u0/ethc0/r_reg[tmsto][addr] [3]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][addr] [2]),
        .I3(\r[bb]_i_4_n_0 ),
        .I4(\r[bb]_i_5_n_0 ),
        .I5(\r[bb]_i_6_n_0 ),
        .O(\m100.u0/ethc0/ahb0/v ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCD88)) 
    \r[bb]_i_3 
       (.I0(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .O(\m100.u0/ethc0/ahb0/nbo ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \r[bb]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [6]),
        .I1(\m100.u0/ethc0/r_reg[tmsto][addr] [7]),
        .I2(\m100.u0/ethc0/r_reg[tmsto][addr] [4]),
        .I3(\m100.u0/ethc0/r_reg[tmsto][addr] [5]),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [9]),
        .I5(\m100.u0/ethc0/r_reg[tmsto][addr] [8]),
        .O(\r[bb]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \r[bb]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[rmsto][addr] [6]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [7]),
        .I2(\m100.u0/ethc0/r_reg[rmsto][addr] [4]),
        .I3(\m100.u0/ethc0/r_reg[rmsto][addr] [5]),
        .I4(\m100.u0/ethc0/r_reg[rmsto][addr] [9]),
        .I5(\m100.u0/ethc0/r_reg[rmsto][addr] [8]),
        .O(\r[bb]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0808080008088888)) 
    \r[bb]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rmsto][addr] [3]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [2]),
        .I2(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I3(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I4(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I5(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .O(\r[bb]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    \r[bcast]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [5]),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [7]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [8]),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [13]),
        .I4(\r[bcast]_i_12_n_0 ),
        .O(\r[bcast]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \r[bcast]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [27]),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [16]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [29]),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [28]),
        .O(\r[bcast]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \r[bcast]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [4]),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [2]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [11]),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [1]),
        .O(\r[bcast]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \r[bcast]_i_2 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .O(\m100.u0/ethc0/v[addrok] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFABF)) 
    \r[bcast]_i_3 
       (.I0(\r[msbgood]_i_4_n_0 ),
        .I1(\r[bcast]_i_5_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .O(\r[bcast]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[bcast]_i_4 
       (.I0(\r[bcast]_i_5_n_0 ),
        .I1(\r[bcast]_i_6_n_0 ),
        .O(\r[bcast]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    \r[bcast]_i_5 
       (.I0(\r[bcast]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [18]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [17]),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [20]),
        .I4(\m100.u0/ethc0/r_reg[checkdata]__0 [19]),
        .I5(\r[bcast]_i_8_n_0 ),
        .O(\r[bcast]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    \r[bcast]_i_6 
       (.I0(\r[bcast]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [6]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [3]),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [14]),
        .I4(\m100.u0/ethc0/r_reg[checkdata]__0 [12]),
        .I5(\r[bcast]_i_10_n_0 ),
        .O(\r[bcast]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \r[bcast]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [22]),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [21]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [24]),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [23]),
        .O(\r[bcast]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    \r[bcast]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [30]),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [31]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [25]),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [26]),
        .I4(\r[bcast]_i_11_n_0 ),
        .O(\r[bcast]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \r[bcast]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [10]),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [9]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [15]),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [0]),
        .O(\r[bcast]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[bg]_i_1 
       (.I0(ahbmi[6]),
        .I1(\ahbmi[hready] ),
        .I2(\m100.u0/ethc0/ahb0/r_reg[bg]__0 ),
        .O(\r[bg]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFAFF1000)) 
    \r[bo]_i_1 
       (.I0(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I1(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I3(\ahbmi[hready] ),
        .I4(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[bo]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h57005500)) 
    \r[capbil][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][6] ),
        .I4(\m100.u0/ethc0/r_reg[capbil_n_0_][1] ),
        .O(\r[capbil][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h57005500)) 
    \r[capbil][2]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][7] ),
        .I4(\m100.u0/ethc0/r_reg[capbil_n_0_][2] ),
        .O(\r[capbil][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h57005500)) 
    \r[capbil][3]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I3(\m100.u0/ethc0/p_1_in128_in ),
        .I4(\m100.u0/ethc0/p_116_in ),
        .O(\r[capbil][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00240000)) 
    \r[capbil][4]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .O(\r[capbil][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h57005500)) 
    \r[capbil][4]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][9] ),
        .I4(\m100.u0/ethc0/p_0_in1_in ),
        .O(\r[capbil][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0080)) 
    \r[checkdata][31]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\m100.u0/ethc0/rmsti[ready] ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .O(\m100.u0/ethc0/v[check] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0022002205FF04AA)) 
    \r[cnt][0]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I2(\r[cnt][0]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I5(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .O(\r[cnt][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \r[cnt][0]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .O(\r[cnt][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2442277224422222)) 
    \r[cnt][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I5(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .O(\r[cnt][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F4A40404A4A4040)) 
    \r[cnt][2]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I1(\r[cnt][2]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I3(\r[cnt][2]_i_3_n_0 ),
        .I4(\r[cnt][2]_i_4_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .O(\r[cnt][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00EEEE0EEE000000)) 
    \r[cnt][2]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I2(\r[cnt][2]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .O(\r[cnt][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    \r[cnt][2]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .O(\r[cnt][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE1FF)) 
    \r[cnt][2]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .O(\r[cnt][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \r[cnt][2]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .O(\r[cnt][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5F0A50004A0A4000)) 
    \r[cnt][3]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I3(\r[cnt][3]_i_2_n_0 ),
        .I4(\r[cnt][3]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .O(\r[cnt][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \r[cnt][3]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .O(\r[cnt][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFE01FFFF)) 
    \r[cnt][3]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .O(\r[cnt][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000003770000)) 
    \r[cnt][4]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I4(\etho[mdc] ),
        .I5(\m100.u0/ethc0/p_1_in143_in ),
        .O(\m100.u0/ethc0/v[cnt] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h33BB008830800080)) 
    \r[cnt][4]_i_2 
       (.I0(\r[cnt][4]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\r[cnt][4]_i_4_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .O(\r[cnt][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAAAA9)) 
    \r[cnt][4]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .O(\r[cnt][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \r[cnt][4]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .O(\r[cnt][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5455)) 
    \r[ctrl][full_duplex]_i_2 
       (.I0(\m100.u0/ethc0/p_116_in ),
        .I1(\m100.u0/ethc0/r_reg[capbil_n_0_][2] ),
        .I2(\m100.u0/ethc0/p_0_in1_in ),
        .I3(\m100.u0/ethc0/r_reg[capbil_n_0_][1] ),
        .O(\r[ctrl][full_duplex]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[ctrl][full_duplex]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .O(\r[ctrl][full_duplex]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFFF3F3B00000008)) 
    \r[ctrl][rxen]_i_2 
       (.I0(\r[ctrl][rxen]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I2(\m100.u0/ethc0/rmsti ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\apbi[pwdata] [1]),
        .O(\m100.u0/ethc0/v[ctrl][rxen] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF3000C0C8)) 
    \r[ctrl][rxen]_i_3 
       (.I0(\r[ctrl][rxen]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I2(\m100.u0/ethc0/rmsti ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/v[ctrl][txen] ),
        .O(\r[ctrl][rxen]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0020)) 
    \r[ctrl][rxen]_i_4 
       (.I0(\ahbmi[hrdata] [11]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/rmsti[ready] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I4(\apbi[pwdata] [1]),
        .O(\r[ctrl][rxen]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \r[ctrl][rxen]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/rmsti[ready] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .O(\r[ctrl][rxen]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r[ctrl][speed]_i_1 
       (.I0(\m100.u0/ethc0/p_6_in [6]),
        .I1(rst),
        .O(\r[ctrl][speed]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4040404040404000)) 
    \r[ctrl][speed]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[capbil_n_0_][2] ),
        .I4(\m100.u0/ethc0/p_0_in1_in ),
        .I5(\m100.u0/ethc0/p_116_in ),
        .O(\r[ctrl][speed]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \r[ctrl][tx_irqen]_i_1 
       (.I0(\apbi[penable] ),
        .I1(apbi[15]),
        .I2(\apbi[pwrite] ),
        .I3(\apbo[prdata][14]_INST_0_i_2_n_0 ),
        .O(\m100.u0/ethc0/v[ctrl][txen] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0404040400000200)) 
    \r[ctrl][txen]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/tmsti[ready] ),
        .I4(\r[ctrl][txen]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[ctrl][txen]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r[ctrl][txen]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .O(\r[ctrl][txen]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \r[ctrlpkt]_i_2 
       (.I0(\r_reg[rxcnt][10]_i_8_n_2 ),
        .I1(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I2(\m100.u0/ethc0/p_0_in153_in ),
        .O(\m100.u0/ethc0/v[ctrlpkt]69_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[ctrlpkt]_i_3 
       (.I0(\m100.u0/ethc0/v ),
        .I1(\r[ctrlpkt]_i_4_n_0 ),
        .O(\m100.u0/ethc0/v[ctrlpkt]68_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFB)) 
    \r[ctrlpkt]_i_4 
       (.I0(\r[ctrlpkt]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [31]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [30]),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [20]),
        .I4(\m100.u0/ethc0/r_reg[checkdata]__0 [17]),
        .I5(\r[ctrlpkt]_i_6_n_0 ),
        .O(\r[ctrlpkt]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r[ctrlpkt]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [24]),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [21]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [22]),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [18]),
        .O(\r[ctrlpkt]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    \r[ctrlpkt]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [28]),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [29]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [25]),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [19]),
        .I4(\r[ctrlpkt]_i_7_n_0 ),
        .O(\r[ctrlpkt]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFD)) 
    \r[ctrlpkt]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [27]),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [26]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [23]),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [16]),
        .O(\r[ctrlpkt]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF550F04FF550004)) 
    \r[duplexstate][0]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I1(\r[duplexstate][0]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I4(\r[duplexstate][1]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[init_busy_n_0_] ),
        .O(\r[duplexstate][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[duplexstate][0]_i_2 
       (.I0(\m100.u0/ethc0/p_6_in [12]),
        .I1(\m100.u0/ethc0/p_6_in [14]),
        .O(\r[duplexstate][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF100F1F1)) 
    \r[duplexstate][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rstphy]__0 ),
        .I1(\r[duplexstate][1]_i_2_n_0 ),
        .I2(\r[duplexstate][1]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .O(\r[duplexstate][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFD)) 
    \r[duplexstate][1]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][linkfail_n_0_] ),
        .I3(\m100.u0/ethc0/r_reg[init_busy_n_0_] ),
        .O(\r[duplexstate][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAEAA)) 
    \r[duplexstate][1]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I3(\r[duplexstate][1]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I5(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .O(\r[duplexstate][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAABAA)) 
    \r[duplexstate][1]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I1(\m100.u0/ethc0/p_6_in [12]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][15] ),
        .I3(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rstaneg_n_0_] ),
        .O(\r[duplexstate][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r[duplexstate][2]_i_1 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][write]113_out ),
        .I1(rst),
        .O(\r[duplexstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFAAAAFFFF0200)) 
    \r[duplexstate][2]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I3(\m100.u0/ethc0/p_6_in [12]),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .O(\r[duplexstate][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFEFEFE00)) 
    \r[duplexstate][2]_i_3 
       (.I0(\r[duplexstate][1]_i_1_n_0 ),
        .I1(\r[duplexstate][2]_i_2_n_0 ),
        .I2(\r[duplexstate][0]_i_1_n_0 ),
        .I3(\m100.u0/ethc0/p_6_in [14]),
        .I4(\m100.u0/ethc0/p_6_in [12]),
        .O(\m100.u0/ethc0/v[mdio_ctrl][write]113_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h002A)) 
    \r[ecnt][0]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\r[ecnt][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h002A2A00)) 
    \r[ecnt][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\m100.u0/ethc0/v[ecnt] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h002A2A2A2A000000)) 
    \r[ecnt][2]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .O(\m100.u0/ethc0/v[ecnt] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0028000000007D00)) 
    \r[ecnt][3]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I2(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\r[ecnt][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h002A2A2A2A000000)) 
    \r[ecnt][3]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\r[ecnt][3]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\m100.u0/ethc0/v[ecnt] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[ecnt][3]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\r[ecnt][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[edclactive]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][11] ),
        .I1(\m100.u0/rxwdata [27]),
        .I2(\m100.u0/rxwdata [25]),
        .I3(\m100.u0/ethc0/r_reg[edclip_n_0_][9] ),
        .I4(\m100.u0/rxwdata [26]),
        .I5(\m100.u0/ethc0/r_reg[edclip_n_0_][10] ),
        .O(\r[edclactive]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[edclactive]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][7] ),
        .I1(\m100.u0/rxwdata [23]),
        .I2(\m100.u0/rxwdata [24]),
        .I3(\m100.u0/ethc0/r_reg[edclip_n_0_][8] ),
        .I4(\m100.u0/rxwdata [22]),
        .I5(\m100.u0/ethc0/r_reg[edclip_n_0_][6] ),
        .O(\r[edclactive]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[edclactive]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][4] ),
        .I1(\m100.u0/rxwdata [20]),
        .I2(\m100.u0/rxwdata [21]),
        .I3(\m100.u0/ethc0/r_reg[edclip_n_0_][5] ),
        .I4(\m100.u0/rxwdata [19]),
        .I5(\m100.u0/ethc0/r_reg[edclip_n_0_][3] ),
        .O(\r[edclactive]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[edclactive]_i_13 
       (.I0(\m100.u0/rxwdata [18]),
        .I1(\m100.u0/ethc0/r_reg[edclip_n_0_][2] ),
        .I2(\m100.u0/rxwdata [16]),
        .I3(\m100.u0/ethc0/r_reg[edclip_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[edclip_n_0_][1] ),
        .I5(\m100.u0/rxwdata [17]),
        .O(\r[edclactive]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \r[edclactive]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I4(\m100.u0/ethc0/v[writeok]1 ),
        .I5(\r_reg[edclactive]_i_6_n_2 ),
        .O(\m100.u0/ethc0/v[edclactive]58_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[edclactive]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\r[edclactive]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F00030008000000)) 
    \r[edclactive]_i_4 
       (.I0(\m100.u0/ethc0/v[edclactive]58_out ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\m100.u0/ethc0/v[addrok] ),
        .O(\r[edclactive]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0FEF0FEF00010000)) 
    \r[edclactive]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/v[edclrstate]0 ),
        .I5(\m100.u0/ethc0/v[addrok] ),
        .O(\r[edclactive]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r[edclactive]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][15] ),
        .I1(\m100.u0/rxwdata [31]),
        .O(\r[edclactive]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[edclactive]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[edclip_n_0_][14] ),
        .I1(\m100.u0/rxwdata [30]),
        .I2(\m100.u0/rxwdata [28]),
        .I3(\m100.u0/ethc0/r_reg[edclip_n_0_][12] ),
        .I4(\m100.u0/rxwdata [29]),
        .I5(\m100.u0/ethc0/r_reg[edclip_n_0_][13] ),
        .O(\r[edclactive]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0101000100010001)) 
    \r[edclbcast]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/v[writeok]1 ),
        .I5(\FSM_sequential_r[edclrstate][3]_i_15_n_0 ),
        .O(\r[edclbcast]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4000000000000000)) 
    \r[edclip][31]_i_1 
       (.I0(\apbo[prdata][14]_INST_0_i_5_n_0 ),
        .I1(\apbi[pwrite] ),
        .I2(apbi[15]),
        .I3(\apbi[penable] ),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [2]),
        .O(\m100.u0/ethc0/v[edclip] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0080)) 
    \r[emacaddr][31]_i_1 
       (.I0(\apbi[penable] ),
        .I1(apbi[15]),
        .I2(\apbi[pwrite] ),
        .I3(\r[emacaddr][31]_i_2_n_0 ),
        .O(\m100.u0/ethc0/v[emacaddr] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hDFFF)) 
    \r[emacaddr][31]_i_2 
       (.I0(\apbi[paddr] [5]),
        .I1(\apbi[paddr] [4]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [2]),
        .O(\r[emacaddr][31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00004000)) 
    \r[emacaddr][47]_i_1 
       (.I0(\apbi[paddr] [2]),
        .I1(\apbi[paddr] [3]),
        .I2(\r[mdio_ctrl][phyadr][4]_i_2_n_0 ),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [4]),
        .O(\m100.u0/ethc0/v[emacaddr] [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5554)) 
    \r[erenable]_i_2 
       (.I0(\m100.u0/ethc0/p_6_in [14]),
        .I1(\m100.u0/ethc0/r_reg ),
        .I2(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[abufs_n_0_][2] ),
        .O(\m100.u0/ethc0/v[tmsto][req]1149_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0020)) 
    \r[error]_i_1 
       (.I0(\ahbmi[hresp] [0]),
        .I1(\ahbmi[hresp] [1]),
        .I2(\m100.u0/ethc0/ahb0/r_reg ),
        .I3(\ahbmi[hready] ),
        .O(\r[error]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[erxidle]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .O(\r[erxidle]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r[erxidle]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\r[erxidle]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \r[etxidle]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[abufs_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg ),
        .O(\m100.u0/ethc0/rin ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00080000)) 
    \r[ewr]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\r[ewr]_i_2_n_0 ),
        .O(\m100.u0/ethc0/v[nak] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1400000000000000)) 
    \r[ewr]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I2(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\r[ewr]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \r[init_busy]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .I2(\etho[mdc] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .O(\r[init_busy]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][0]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [0]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][10]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [10]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [10]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][11]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [11]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [11]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6696AAAA66965555)) 
    \r[ipcrc][11]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][9] ),
        .I1(\r[ipcrc][11]_i_12_n_0 ),
        .I2(\m100.u0/rxwdata [16]),
        .I3(\r[ipcrc][11]_i_13_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I5(\m100.u0/rxwdata [25]),
        .O(\r[ipcrc][11]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h59A959A9A95959A9)) 
    \r[ipcrc][11]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][8] ),
        .I1(\m100.u0/rxwdata [24]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\r[ipcrc][11]_i_14_n_0 ),
        .I4(\m100.u0/rxwdata [15]),
        .I5(\r[ipcrc][11]_i_13_n_0 ),
        .O(\r[ipcrc][11]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00A8000000000000)) 
    \r[ipcrc][11]_i_12 
       (.I0(\m100.u0/rxwdata [15]),
        .I1(\r[ipcrc][7]_i_14_n_0 ),
        .I2(\m100.u0/rxwdata [12]),
        .I3(\r[ipcrc][11]_i_13_n_0 ),
        .I4(\m100.u0/rxwdata [13]),
        .I5(\m100.u0/rxwdata [14]),
        .O(\r[ipcrc][11]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r[ipcrc][11]_i_13 
       (.I0(\m100.u0/rxwdata [17]),
        .I1(\m100.u0/ethc0/v[nak]1 ),
        .O(\r[ipcrc][11]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0080008000800000)) 
    \r[ipcrc][11]_i_14 
       (.I0(\m100.u0/rxwdata [14]),
        .I1(\m100.u0/rxwdata [13]),
        .I2(\m100.u0/ethc0/v[nak]1 ),
        .I3(\m100.u0/rxwdata [17]),
        .I4(\m100.u0/rxwdata [12]),
        .I5(\r[ipcrc][7]_i_14_n_0 ),
        .O(\r[ipcrc][11]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \r[ipcrc][11]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][11] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I2(\m100.u0/rxwdata [27]),
        .O(\r[ipcrc][11]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h59A9A9A9)) 
    \r[ipcrc][11]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][10] ),
        .I1(\m100.u0/rxwdata [26]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/rxwdata [16]),
        .I4(\r[ipcrc][11]_i_12_n_0 ),
        .O(\r[ipcrc][11]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][12]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [12]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [12]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][13]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [13]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [13]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][14]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [14]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [14]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][15]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [15]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [15]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \r[ipcrc][15]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][13] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I2(\m100.u0/rxwdata [29]),
        .O(\r[ipcrc][15]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \r[ipcrc][15]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][12] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I2(\m100.u0/rxwdata [28]),
        .O(\r[ipcrc][15]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \r[ipcrc][15]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][15] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I2(\m100.u0/rxwdata [31]),
        .O(\r[ipcrc][15]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \r[ipcrc][15]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][14] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I2(\m100.u0/rxwdata [30]),
        .O(\r[ipcrc][15]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][16]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [16]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [16]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040004044440044)) 
    \r[ipcrc][17]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/v[rxstatus]2 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\r[ipcrc][17]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\r[ipcrc][17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0400)) 
    \r[ipcrc][17]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [17]),
        .O(\m100.u0/ethc0/v[ipcrc] [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000660000606)) 
    \r[ipcrc][17]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I1(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\r[ipcrc][17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [1]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [1]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][2]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [2]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [2]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][3]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [3]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69656565)) 
    \r[ipcrc][3]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\m100.u0/rxwdata [17]),
        .I3(\m100.u0/ethc0/v[nak]1 ),
        .I4(\m100.u0/rxwdata [8]),
        .O(\r[ipcrc][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA959A9A9A9A9A9A9)) 
    \r[ipcrc][3]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][0] ),
        .I1(\m100.u0/rxwdata [16]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/rxwdata [17]),
        .I4(\m100.u0/ethc0/v[nak]1 ),
        .I5(\m100.u0/rxwdata [7]),
        .O(\r[ipcrc][3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCFDF)) 
    \r[ipcrc][3]_i_12 
       (.I0(\m100.u0/rxwdata [9]),
        .I1(\m100.u0/rxwdata [17]),
        .I2(\m100.u0/ethc0/v[nak]1 ),
        .I3(\m100.u0/rxwdata [8]),
        .O(\r[ipcrc][3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[ipcrc][3]_i_6 
       (.I0(\m100.u0/ethc0/a [1]),
        .I1(\m100.u0/ethc0/r_reg[ipcrc_n_0_][1] ),
        .O(\r[ipcrc][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[ipcrc][3]_i_7 
       (.I0(\m100.u0/ethc0/a [0]),
        .I1(\m100.u0/ethc0/r_reg[ipcrc_n_0_][0] ),
        .O(\r[ipcrc][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9699AAAA96995555)) 
    \r[ipcrc][3]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][3] ),
        .I1(\r[ipcrc][3]_i_12_n_0 ),
        .I2(\r[ipcrc][11]_i_13_n_0 ),
        .I3(\m100.u0/rxwdata [10]),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I5(\m100.u0/rxwdata [19]),
        .O(\r[ipcrc][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h595959A95959A959)) 
    \r[ipcrc][3]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][2] ),
        .I1(\m100.u0/rxwdata [18]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/rxwdata [8]),
        .I4(\r[ipcrc][11]_i_13_n_0 ),
        .I5(\m100.u0/rxwdata [9]),
        .O(\r[ipcrc][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][4]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [4]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [4]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][5]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [5]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [5]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][6]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [6]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [6]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][7]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [7]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [7]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA959A95959A9A959)) 
    \r[ipcrc][7]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][5] ),
        .I1(\m100.u0/rxwdata [21]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\r[ipcrc][7]_i_14_n_0 ),
        .I4(\m100.u0/rxwdata [12]),
        .I5(\r[ipcrc][11]_i_13_n_0 ),
        .O(\r[ipcrc][7]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA959A9A959A95959)) 
    \r[ipcrc][7]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][4] ),
        .I1(\m100.u0/rxwdata [20]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\r[ipcrc][11]_i_13_n_0 ),
        .I4(\m100.u0/rxwdata [11]),
        .I5(\r[ipcrc][7]_i_15_n_0 ),
        .O(\r[ipcrc][7]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF1FFFFFF)) 
    \r[ipcrc][7]_i_12 
       (.I0(\r[ipcrc][7]_i_14_n_0 ),
        .I1(\m100.u0/rxwdata [12]),
        .I2(\m100.u0/rxwdata [17]),
        .I3(\m100.u0/ethc0/v[nak]1 ),
        .I4(\m100.u0/rxwdata [13]),
        .O(\r[ipcrc][7]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF11FF15FF55FF55)) 
    \r[ipcrc][7]_i_13 
       (.I0(\m100.u0/rxwdata [12]),
        .I1(\m100.u0/rxwdata [10]),
        .I2(\m100.u0/rxwdata [8]),
        .I3(\r[ipcrc][11]_i_13_n_0 ),
        .I4(\m100.u0/rxwdata [9]),
        .I5(\m100.u0/rxwdata [11]),
        .O(\r[ipcrc][7]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0A00080000000000)) 
    \r[ipcrc][7]_i_14 
       (.I0(\m100.u0/rxwdata [11]),
        .I1(\m100.u0/rxwdata [9]),
        .I2(\m100.u0/rxwdata [17]),
        .I3(\m100.u0/ethc0/v[nak]1 ),
        .I4(\m100.u0/rxwdata [8]),
        .I5(\m100.u0/rxwdata [10]),
        .O(\r[ipcrc][7]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF5FFF7F)) 
    \r[ipcrc][7]_i_15 
       (.I0(\m100.u0/rxwdata [10]),
        .I1(\m100.u0/rxwdata [8]),
        .I2(\m100.u0/ethc0/v[nak]1 ),
        .I3(\m100.u0/rxwdata [17]),
        .I4(\m100.u0/rxwdata [9]),
        .O(\r[ipcrc][7]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA959A95959A9A959)) 
    \r[ipcrc][7]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][7] ),
        .I1(\m100.u0/rxwdata [23]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\r[ipcrc][7]_i_12_n_0 ),
        .I4(\m100.u0/rxwdata [14]),
        .I5(\r[ipcrc][11]_i_13_n_0 ),
        .O(\r[ipcrc][7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9969AAAA99695555)) 
    \r[ipcrc][7]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[ipcrc_n_0_][6] ),
        .I1(\r[ipcrc][7]_i_13_n_0 ),
        .I2(\m100.u0/rxwdata [13]),
        .I3(\r[ipcrc][11]_i_13_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I5(\m100.u0/rxwdata [22]),
        .O(\r[ipcrc][7]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][8]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [8]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [8]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44444444CFC00000)) 
    \r[ipcrc][9]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/crcadder [9]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/p_1_in [9]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[ipcrc] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02000000)) 
    \r[mac_addr][31]_i_1 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[paddr] [5]),
        .I2(\apbi[paddr] [4]),
        .I3(\r[mdio_ctrl][phyadr][4]_i_2_n_0 ),
        .I4(\apbi[paddr] [2]),
        .O(\m100.u0/ethc0/v[mac_addr] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h01000000)) 
    \r[mac_addr][47]_i_1 
       (.I0(\apbi[paddr] [4]),
        .I1(\apbi[paddr] [5]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\r[mdio_ctrl][phyadr][4]_i_2_n_0 ),
        .O(\m100.u0/ethc0/v[mac_addr] [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FFFF0000FFFE)) 
    \r[mdccnt][0]_i_1 
       (.I0(\m100.u0/ethc0/d [3]),
        .I1(\m100.u0/ethc0/d [4]),
        .I2(\m100.u0/ethc0/d [5]),
        .I3(\m100.u0/ethc0/d [2]),
        .I4(\m100.u0/ethc0/d [0]),
        .I5(\m100.u0/ethc0/d [1]),
        .O(\m100.u0/ethc0/v[mdccnt] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r[mdccnt][1]_i_1 
       (.I0(\m100.u0/ethc0/d [1]),
        .I1(\m100.u0/ethc0/d [0]),
        .O(\m100.u0/ethc0/v[mdccnt] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE1E1E1E1E1E1E1E0)) 
    \r[mdccnt][2]_i_1 
       (.I0(\m100.u0/ethc0/d [1]),
        .I1(\m100.u0/ethc0/d [0]),
        .I2(\m100.u0/ethc0/d [2]),
        .I3(\m100.u0/ethc0/d [5]),
        .I4(\m100.u0/ethc0/d [4]),
        .I5(\m100.u0/ethc0/d [3]),
        .O(\m100.u0/ethc0/v[mdccnt] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFE01FE01FE01FE00)) 
    \r[mdccnt][3]_i_1 
       (.I0(\m100.u0/ethc0/d [2]),
        .I1(\m100.u0/ethc0/d [0]),
        .I2(\m100.u0/ethc0/d [1]),
        .I3(\m100.u0/ethc0/d [3]),
        .I4(\m100.u0/ethc0/d [4]),
        .I5(\m100.u0/ethc0/d [5]),
        .O(\m100.u0/ethc0/v[mdccnt] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAAAA9)) 
    \r[mdccnt][4]_i_1 
       (.I0(\m100.u0/ethc0/d [4]),
        .I1(\m100.u0/ethc0/d [2]),
        .I2(\m100.u0/ethc0/d [0]),
        .I3(\m100.u0/ethc0/d [1]),
        .I4(\m100.u0/ethc0/d [3]),
        .O(\m100.u0/ethc0/v[mdccnt] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFE00000001)) 
    \r[mdccnt][5]_i_1 
       (.I0(\m100.u0/ethc0/d [2]),
        .I1(\m100.u0/ethc0/d [0]),
        .I2(\m100.u0/ethc0/d [1]),
        .I3(\m100.u0/ethc0/d [3]),
        .I4(\m100.u0/ethc0/d [4]),
        .I5(\m100.u0/ethc0/d [5]),
        .O(\r[mdccnt][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h03AA00AA)) 
    \r[mdio_ctrl][busy]_i_2 
       (.I0(\r[mdio_ctrl][busy]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\r[mdio_ctrl][busy]_i_6_n_0 ),
        .O(\r[mdio_ctrl][busy]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA22AA22AA022202)) 
    \r[mdio_ctrl][busy]_i_3 
       (.I0(\r[rstaneg]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/v[mdio_ctrl][busy] ),
        .I2(\m100.u0/ethc0/p_6_in [12]),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I5(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .O(\r[mdio_ctrl][busy]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00800000)) 
    \r[mdio_ctrl][busy]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I2(\r[mdio_ctrl][busy]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\m100.u0/ethc0/v[mdio_ctrl][busy] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h007FFFFF00000000)) 
    \r[mdio_ctrl][busy]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I2(\r[mdio_ctrl][busy]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\m100.u0/ethc0/v[mdio_ctrl][busy]0 ),
        .O(\r[mdio_ctrl][busy]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h1A001F00)) 
    \r[mdio_ctrl][busy]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I3(\r[mdio_ctrl][busy]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/p_6_in [12]),
        .O(\r[mdio_ctrl][busy]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAA0008)) 
    \r[mdio_ctrl][busy]_i_7 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][write]1 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/p_6_in [12]),
        .I5(\m100.u0/ethc0/p_6_in [14]),
        .O(\r[mdio_ctrl][busy]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r[mdio_ctrl][busy]_i_8 
       (.I0(\apbi[pwdata] [1]),
        .I1(\apbi[pwdata] [0]),
        .O(\m100.u0/ethc0/v[mdio_ctrl][busy]0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][0]_i_1 
       (.I0(\r[mdio_ctrl][data][0]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][0]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .O(\r[mdio_ctrl][data][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][0]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][0]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][0]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][0]_i_3 
       (.I0(\r[mdio_ctrl][data][0]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][0]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][0]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][0]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [16]),
        .O(\r[mdio_ctrl][data][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC440000FC770000)) 
    \r[mdio_ctrl][data][0]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][0]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][0]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][0]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][0]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][0]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFE00000002)) 
    \r[mdio_ctrl][data][0]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][12]_i_10_n_0 ),
        .I5(\apbi[pwdata] [16]),
        .O(\r[mdio_ctrl][data][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \r[mdio_ctrl][data][0]_i_9 
       (.I0(\r[mdio_ctrl][data][3]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/p_1_in143_in ),
        .I4(\etho[mdc] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .O(\r[mdio_ctrl][data][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][10]_i_1 
       (.I0(\r[mdio_ctrl][data][10]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][10]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][10] ),
        .O(\r[mdio_ctrl][data][10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][10]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][10]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][10]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][10]_i_3 
       (.I0(\r[mdio_ctrl][data][10]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][10]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][10]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][10]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [26]),
        .O(\r[mdio_ctrl][data][10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC440000FC770000)) 
    \r[mdio_ctrl][data][10]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][10]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][10]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][10]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][10]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][10]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][10]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][10]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][10]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEF00000020)) 
    \r[mdio_ctrl][data][10]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][14]_i_10_n_0 ),
        .I5(\apbi[pwdata] [26]),
        .O(\r[mdio_ctrl][data][10]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \r[mdio_ctrl][data][10]_i_9 
       (.I0(\r[mdio_ctrl][data][11]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .I2(\etho[mdc] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .O(\r[mdio_ctrl][data][10]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][11]_i_1 
       (.I0(\r[mdio_ctrl][data][11]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][11]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][11] ),
        .O(\r[mdio_ctrl][data][11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \r[mdio_ctrl][data][11]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .O(\r[mdio_ctrl][data][11]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][11]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][11]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][11]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][11]_i_3 
       (.I0(\r[mdio_ctrl][data][11]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][11]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][11]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][11]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [27]),
        .O(\r[mdio_ctrl][data][11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC440000FC770000)) 
    \r[mdio_ctrl][data][11]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][11]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][11]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][11]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][11]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][11]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][11]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEF00000020)) 
    \r[mdio_ctrl][data][11]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][15]_i_12_n_0 ),
        .I5(\apbi[pwdata] [27]),
        .O(\r[mdio_ctrl][data][11]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \r[mdio_ctrl][data][11]_i_9 
       (.I0(\r[mdio_ctrl][data][11]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/p_1_in143_in ),
        .I4(\etho[mdc] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .O(\r[mdio_ctrl][data][11]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF8FFF800)) 
    \r[mdio_ctrl][data][12]_i_1 
       (.I0(\r[mdio_ctrl][data][15]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rstphy]__0 ),
        .I2(\r[mdio_ctrl][data][12]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][12]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][12] ),
        .O(\r[mdio_ctrl][data][12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFDF)) 
    \r[mdio_ctrl][data][12]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I1(\etho[mdc] ),
        .I2(\m100.u0/ethc0/p_1_in143_in ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .O(\r[mdio_ctrl][data][12]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF10FF00EF00)) 
    \r[mdio_ctrl][data][12]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I3(\r[mdio_ctrl][data][12]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][12]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][12]_i_3 
       (.I0(\r[mdio_ctrl][data][12]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][12]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][12]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][12]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [28]),
        .O(\r[mdio_ctrl][data][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCCC0088FCFF0088)) 
    \r[mdio_ctrl][data][12]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][12]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][12]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][12]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][12]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][12]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][12]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][12]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFEFFF00002000)) 
    \r[mdio_ctrl][data][12]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][12]_i_10_n_0 ),
        .I5(\apbi[pwdata] [28]),
        .O(\r[mdio_ctrl][data][12]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \r[mdio_ctrl][data][12]_i_9 
       (.I0(\r[mdio_ctrl][data][15]_i_13_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/p_1_in143_in ),
        .I4(\etho[mdc] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .O(\r[mdio_ctrl][data][12]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][13]_i_1 
       (.I0(\r[mdio_ctrl][data][13]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][13]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][13] ),
        .O(\r[mdio_ctrl][data][13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFDFFFFF)) 
    \r[mdio_ctrl][data][13]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I3(\etho[mdc] ),
        .I4(\m100.u0/ethc0/p_1_in143_in ),
        .O(\r[mdio_ctrl][data][13]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][13]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][13]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][13]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][13]_i_3 
       (.I0(\r[mdio_ctrl][data][13]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][13]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][13]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][13]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [29]),
        .O(\r[mdio_ctrl][data][13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCCC0088FCFF0088)) 
    \r[mdio_ctrl][data][13]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][13]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][13]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][13]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][13]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][13]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][13]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][13]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][13]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFEFFF00002000)) 
    \r[mdio_ctrl][data][13]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][13]_i_10_n_0 ),
        .I5(\apbi[pwdata] [29]),
        .O(\r[mdio_ctrl][data][13]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \r[mdio_ctrl][data][13]_i_9 
       (.I0(\r[mdio_ctrl][data][15]_i_13_n_0 ),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .I2(\etho[mdc] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .O(\r[mdio_ctrl][data][13]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][14]_i_1 
       (.I0(\r[mdio_ctrl][data][14]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][14]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][14] ),
        .O(\r[mdio_ctrl][data][14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFDFFFFF)) 
    \r[mdio_ctrl][data][14]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I3(\etho[mdc] ),
        .I4(\m100.u0/ethc0/p_1_in143_in ),
        .O(\r[mdio_ctrl][data][14]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][14]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][14]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][14]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][14]_i_3 
       (.I0(\r[mdio_ctrl][data][14]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][14]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][14]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][14]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [30]),
        .O(\r[mdio_ctrl][data][14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC440000FC770000)) 
    \r[mdio_ctrl][data][14]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][14]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][14]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][14]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][14]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][14]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][14]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][14]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][14]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFEFFF00002000)) 
    \r[mdio_ctrl][data][14]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][14]_i_10_n_0 ),
        .I5(\apbi[pwdata] [30]),
        .O(\r[mdio_ctrl][data][14]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \r[mdio_ctrl][data][14]_i_9 
       (.I0(\r[mdio_ctrl][data][15]_i_13_n_0 ),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .I2(\etho[mdc] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .O(\r[mdio_ctrl][data][14]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF8FFF800)) 
    \r[mdio_ctrl][data][15]_i_1 
       (.I0(\r[mdio_ctrl][data][15]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rstphy]__0 ),
        .I2(\r[mdio_ctrl][data][15]_i_3_n_0 ),
        .I3(\r[mdio_ctrl][data][15]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][15] ),
        .O(\r[mdio_ctrl][data][15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFEFFF00002000)) 
    \r[mdio_ctrl][data][15]_i_10 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][15]_i_12_n_0 ),
        .I5(\apbi[pwdata] [31]),
        .O(\r[mdio_ctrl][data][15]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \r[mdio_ctrl][data][15]_i_11 
       (.I0(\r[mdio_ctrl][data][15]_i_13_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/p_1_in143_in ),
        .I4(\etho[mdc] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .O(\r[mdio_ctrl][data][15]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDFFFFFFF)) 
    \r[mdio_ctrl][data][15]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I1(\etho[mdc] ),
        .I2(\m100.u0/ethc0/p_1_in143_in ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .O(\r[mdio_ctrl][data][15]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \r[mdio_ctrl][data][15]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .O(\r[mdio_ctrl][data][15]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \r[mdio_ctrl][data][15]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/p_6_in [12]),
        .I3(\m100.u0/ethc0/p_6_in [14]),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .O(\r[mdio_ctrl][data][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF10FF00EF00)) 
    \r[mdio_ctrl][data][15]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I3(\r[mdio_ctrl][data][15]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][15]_i_6_n_0 ),
        .O(\r[mdio_ctrl][data][15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFA8FF08AA08AA)) 
    \r[mdio_ctrl][data][15]_i_4 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\r[mdio_ctrl][data][15]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][15]_i_9_n_0 ),
        .O(\r[mdio_ctrl][data][15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][15]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][15]_i_10_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [31]),
        .O(\r[mdio_ctrl][data][15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC440000FC770000)) 
    \r[mdio_ctrl][data][15]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][15]_i_5_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1010101010101110)) 
    \r[mdio_ctrl][data][15]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[rstphy]__0 ),
        .I4(\m100.u0/ethc0/p_6_in [14]),
        .I5(\m100.u0/ethc0/p_6_in [12]),
        .O(\r[mdio_ctrl][data][15]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][15]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][15]_i_9_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][15]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][15]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][15]_i_11_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][15]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][1]_i_1 
       (.I0(\r[mdio_ctrl][data][1]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][1]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][1] ),
        .O(\r[mdio_ctrl][data][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][1]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][1]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][1]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][1]_i_3 
       (.I0(\r[mdio_ctrl][data][1]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][1]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][1]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][1]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [17]),
        .O(\r[mdio_ctrl][data][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC440000FC770000)) 
    \r[mdio_ctrl][data][1]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][1]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][1]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][1]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][1]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][1]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFE00000002)) 
    \r[mdio_ctrl][data][1]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][13]_i_10_n_0 ),
        .I5(\apbi[pwdata] [17]),
        .O(\r[mdio_ctrl][data][1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \r[mdio_ctrl][data][1]_i_9 
       (.I0(\r[mdio_ctrl][data][3]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .I2(\etho[mdc] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .O(\r[mdio_ctrl][data][1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][2]_i_1 
       (.I0(\r[mdio_ctrl][data][2]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][2]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][2] ),
        .O(\r[mdio_ctrl][data][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][2]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][2]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][2]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][2]_i_3 
       (.I0(\r[mdio_ctrl][data][2]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][2]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][2]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][2]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [18]),
        .O(\r[mdio_ctrl][data][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC440000FC770000)) 
    \r[mdio_ctrl][data][2]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][2]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][2]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][2]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][2]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][2]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFE00000002)) 
    \r[mdio_ctrl][data][2]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][14]_i_10_n_0 ),
        .I5(\apbi[pwdata] [18]),
        .O(\r[mdio_ctrl][data][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \r[mdio_ctrl][data][2]_i_9 
       (.I0(\r[mdio_ctrl][data][3]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .I2(\etho[mdc] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .O(\r[mdio_ctrl][data][2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][3]_i_1 
       (.I0(\r[mdio_ctrl][data][3]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][3]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][3] ),
        .O(\r[mdio_ctrl][data][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \r[mdio_ctrl][data][3]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .O(\r[mdio_ctrl][data][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][3]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][3]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][3]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][3]_i_3 
       (.I0(\r[mdio_ctrl][data][3]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][3]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][3]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][3]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [19]),
        .O(\r[mdio_ctrl][data][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC440000FC770000)) 
    \r[mdio_ctrl][data][3]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][3]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][3]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][3]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][3]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][3]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFE00000002)) 
    \r[mdio_ctrl][data][3]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][15]_i_12_n_0 ),
        .I5(\apbi[pwdata] [19]),
        .O(\r[mdio_ctrl][data][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \r[mdio_ctrl][data][3]_i_9 
       (.I0(\r[mdio_ctrl][data][3]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/p_1_in143_in ),
        .I4(\etho[mdc] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .O(\r[mdio_ctrl][data][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][4]_i_1 
       (.I0(\r[mdio_ctrl][data][4]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][4]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][4] ),
        .O(\r[mdio_ctrl][data][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][4]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][4]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][4]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][4]_i_3 
       (.I0(\r[mdio_ctrl][data][4]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][4]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][4]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][4]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [20]),
        .O(\r[mdio_ctrl][data][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC440000FC770000)) 
    \r[mdio_ctrl][data][4]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][4]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][4]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][4]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][4]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][4]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEFF00000200)) 
    \r[mdio_ctrl][data][4]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][12]_i_10_n_0 ),
        .I5(\apbi[pwdata] [20]),
        .O(\r[mdio_ctrl][data][4]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \r[mdio_ctrl][data][4]_i_9 
       (.I0(\r[cnt][2]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/p_1_in143_in ),
        .I4(\etho[mdc] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .O(\r[mdio_ctrl][data][4]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][5]_i_1 
       (.I0(\r[mdio_ctrl][data][5]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][5]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][5] ),
        .O(\r[mdio_ctrl][data][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][5]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][5]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][5]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][5]_i_3 
       (.I0(\r[mdio_ctrl][data][5]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][5]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][5]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][5]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [21]),
        .O(\r[mdio_ctrl][data][5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC440000FC770000)) 
    \r[mdio_ctrl][data][5]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][5]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][5]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][5]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][5]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][5]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][5]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEFF00000200)) 
    \r[mdio_ctrl][data][5]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][13]_i_10_n_0 ),
        .I5(\apbi[pwdata] [21]),
        .O(\r[mdio_ctrl][data][5]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \r[mdio_ctrl][data][5]_i_9 
       (.I0(\r[cnt][2]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .I2(\etho[mdc] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .O(\r[mdio_ctrl][data][5]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][6]_i_1 
       (.I0(\r[mdio_ctrl][data][6]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][6]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][6] ),
        .O(\r[mdio_ctrl][data][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][6]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][6]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][6]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][6]_i_3 
       (.I0(\r[mdio_ctrl][data][6]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][6]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][6]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][6]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [22]),
        .O(\r[mdio_ctrl][data][6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC440000FC770000)) 
    \r[mdio_ctrl][data][6]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][6]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][6]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][6]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][6]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][6]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][6]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEFF00000200)) 
    \r[mdio_ctrl][data][6]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][14]_i_10_n_0 ),
        .I5(\apbi[pwdata] [22]),
        .O(\r[mdio_ctrl][data][6]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \r[mdio_ctrl][data][6]_i_9 
       (.I0(\r[cnt][2]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .I2(\etho[mdc] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .O(\r[mdio_ctrl][data][6]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][7]_i_1 
       (.I0(\r[mdio_ctrl][data][7]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][7]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][7] ),
        .O(\r[mdio_ctrl][data][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][7]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][7]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][7]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE0FF20F020F0)) 
    \r[mdio_ctrl][data][7]_i_3 
       (.I0(\r[mdio_ctrl][data][7]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I5(\r[mdio_ctrl][data][7]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][7]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][7]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [23]),
        .O(\r[mdio_ctrl][data][7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC440000FC770000)) 
    \r[mdio_ctrl][data][7]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][7]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF03BBFFFF0388)) 
    \r[mdio_ctrl][data][7]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][7]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][7]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][7]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEFF00000200)) 
    \r[mdio_ctrl][data][7]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][15]_i_12_n_0 ),
        .I5(\apbi[pwdata] [23]),
        .O(\r[mdio_ctrl][data][7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \r[mdio_ctrl][data][7]_i_9 
       (.I0(\r[cnt][2]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/p_1_in143_in ),
        .I4(\etho[mdc] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .O(\r[mdio_ctrl][data][7]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][8]_i_1 
       (.I0(\r[mdio_ctrl][data][8]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][8]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/p_1_in128_in ),
        .O(\r[mdio_ctrl][data][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][8]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][8]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][8]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF8F8C8C)) 
    \r[mdio_ctrl][data][8]_i_3 
       (.I0(\r[mdio_ctrl][data][8]_i_6_n_0 ),
        .I1(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I4(\r[mdio_ctrl][data][8]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][8]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][8]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [24]),
        .O(\r[mdio_ctrl][data][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC880088FCBB0088)) 
    \r[mdio_ctrl][data][8]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][8]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF0155FFFF0144)) 
    \r[mdio_ctrl][data][8]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][8]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][8]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][8]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][8]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEF00000020)) 
    \r[mdio_ctrl][data][8]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][12]_i_10_n_0 ),
        .I5(\apbi[pwdata] [24]),
        .O(\r[mdio_ctrl][data][8]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \r[mdio_ctrl][data][8]_i_9 
       (.I0(\r[mdio_ctrl][data][11]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/p_1_in143_in ),
        .I4(\etho[mdc] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .O(\r[mdio_ctrl][data][8]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[mdio_ctrl][data][9]_i_1 
       (.I0(\r[mdio_ctrl][data][9]_i_2_n_0 ),
        .I1(\r[mdio_ctrl][data][9]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][9] ),
        .O(\r[mdio_ctrl][data][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7500753075005500)) 
    \r[mdio_ctrl][data][9]_i_2 
       (.I0(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\r[rstaneg]_i_2_n_0 ),
        .I3(\r[mdio_ctrl][data][9]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I5(\r[mdio_ctrl][data][9]_i_5_n_0 ),
        .O(\r[mdio_ctrl][data][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF8F8C8C)) 
    \r[mdio_ctrl][data][9]_i_3 
       (.I0(\r[mdio_ctrl][data][9]_i_6_n_0 ),
        .I1(\r[mdio_ctrl][data][15]_i_7_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .I4(\r[mdio_ctrl][data][9]_i_7_n_0 ),
        .O(\r[mdio_ctrl][data][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFF00080000)) 
    \r[mdio_ctrl][data][9]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][9]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [25]),
        .O(\r[mdio_ctrl][data][9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC880088FCBB0088)) 
    \r[mdio_ctrl][data][9]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][9]_i_4_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF0155FFFF0144)) 
    \r[mdio_ctrl][data][9]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I4(\r[mdio_ctrl][data][9]_i_7_n_0 ),
        .I5(\r[phywr]_i_4_n_0 ),
        .O(\r[mdio_ctrl][data][9]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFFFFF00080000)) 
    \r[mdio_ctrl][data][9]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdio_ctrl][data][9]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .O(\r[mdio_ctrl][data][9]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEF00000020)) 
    \r[mdio_ctrl][data][9]_i_8 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I4(\r[mdio_ctrl][data][13]_i_10_n_0 ),
        .I5(\apbi[pwdata] [25]),
        .O(\r[mdio_ctrl][data][9]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \r[mdio_ctrl][data][9]_i_9 
       (.I0(\r[mdio_ctrl][data][11]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .I2(\etho[mdc] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .O(\r[mdio_ctrl][data][9]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \r[mdio_ctrl][linkfail]_i_2 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][linkfail]0 ),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .I2(\etho[mdc] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I5(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .O(\r[mdio_ctrl][linkfail]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \r[mdio_ctrl][linkfail]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I1(\etho[mdc] ),
        .I2(\m100.u0/ethc0/p_1_in143_in ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][busy]__0 ),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I5(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .O(\r[mdio_ctrl][linkfail]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \r[mdio_ctrl][phyadr][4]_i_1 
       (.I0(\apbi[paddr] [5]),
        .I1(\apbi[paddr] [4]),
        .I2(\r[mdio_ctrl][phyadr][4]_i_2_n_0 ),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][busy]__0 ),
        .O(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \r[mdio_ctrl][phyadr][4]_i_2 
       (.I0(\apbi[pwrite] ),
        .I1(apbi[15]),
        .I2(\apbi[penable] ),
        .O(\r[mdio_ctrl][phyadr][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h007FFFFF00000000)) 
    \r[mdio_ctrl][read]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I2(\m100.u0/ethc0/v[mdio_ctrl][write]1 ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\apbi[pwdata] [1]),
        .O(\r[mdio_ctrl][read]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \r[mdio_ctrl][read]_i_3 
       (.I0(\r[mdio_ctrl][data][15]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rstphy]__0 ),
        .I2(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .O(\r[mdio_ctrl][read]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h16FF1600)) 
    \r[mdio_ctrl][regadr][0]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I3(\r[mdio_ctrl][data][15]_i_2_n_0 ),
        .I4(\apbi[pwdata] [6]),
        .O(\r[mdio_ctrl][regadr][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    \r[mdio_ctrl][regadr][1]_i_1 
       (.I0(\apbi[pwdata] [7]),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/p_6_in [14]),
        .I3(\m100.u0/ethc0/p_6_in [12]),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .O(\r[mdio_ctrl][regadr][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h24FF2400)) 
    \r[mdio_ctrl][regadr][2]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I3(\r[mdio_ctrl][data][15]_i_2_n_0 ),
        .I4(\apbi[pwdata] [8]),
        .O(\r[mdio_ctrl][regadr][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \r[mdio_ctrl][regadr][3]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I2(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I3(\r[mdio_ctrl][data][15]_i_2_n_0 ),
        .I4(\apbi[pwdata] [9]),
        .O(\r[mdio_ctrl][regadr][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAAB)) 
    \r[mdio_ctrl][regadr][4]_i_1 
       (.I0(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/p_6_in [14]),
        .I3(\m100.u0/ethc0/p_6_in [12]),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .O(\r[mdio_ctrl][regadr][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    \r[mdio_ctrl][regadr][4]_i_2 
       (.I0(\apbi[pwdata] [10]),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/p_6_in [14]),
        .I3(\m100.u0/ethc0/p_6_in [12]),
        .I4(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .O(\r[mdio_ctrl][regadr][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF01FF00)) 
    \r[mdio_ctrl][write]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I3(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .I4(\r[mdio_ctrl][write]_i_8_n_0 ),
        .O(\r[mdio_ctrl][write]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000AAAAEAAA)) 
    \r[mdio_ctrl][write]_i_4 
       (.I0(\r[mdio_ctrl][phyadr][4]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I3(\etho[mdc] ),
        .I4(\m100.u0/ethc0/p_1_in143_in ),
        .I5(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .O(\r[mdio_ctrl][write]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA8)) 
    \r[mdio_ctrl][write]_i_5 
       (.I0(\r[mdio_ctrl][data][15]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rstphy]__0 ),
        .I2(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .O(\r[mdio_ctrl][write]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFE00FF00)) 
    \r[mdio_ctrl][write]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I3(\apbi[pwdata] [0]),
        .I4(\r[mdio_ctrl][write]_i_8_n_0 ),
        .O(\r[mdio_ctrl][write]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000AAAA2AAA)) 
    \r[mdio_ctrl][write]_i_7 
       (.I0(\apbi[pwdata] [0]),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I3(\etho[mdc] ),
        .I4(\m100.u0/ethc0/p_1_in143_in ),
        .I5(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .O(\r[mdio_ctrl][write]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0080)) 
    \r[mdio_ctrl][write]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][busy]__0 ),
        .I1(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I2(\etho[mdc] ),
        .I3(\m100.u0/ethc0/p_1_in143_in ),
        .O(\r[mdio_ctrl][write]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \r[mdioclk]_i_1 
       (.I0(rst),
        .O(\m100.u0/ethc0/ahb0/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r[mdioclk]_i_3 
       (.I0(\m100.u0/ethc0/d [2]),
        .I1(\m100.u0/ethc0/d [0]),
        .I2(\m100.u0/ethc0/d [1]),
        .I3(\m100.u0/ethc0/d [3]),
        .O(\r[mdioclk]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[mdioen]_i_2 
       (.I0(\etho[mdc] ),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .O(\m100.u0/ethc0/v[mdio_ctrl][write]1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0080FFFF00800000)) 
    \r[mdioen]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I1(\m100.u0/ethc0/v[mdio_ctrl][write]1 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I5(\r[mdioen]_i_4_n_0 ),
        .O(\m100.u0/ethc0/v[mdioen] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8080000000000A00)) 
    \r[mdioen]_i_4 
       (.I0(\m100.u0/ethc0/v[mdio_ctrl][write]1 ),
        .I1(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][busy]__0 ),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I5(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .O(\r[mdioen]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r[mdioo]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .O(\r[mdioo]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r[mdioo]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][6] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][5] ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][4] ),
        .O(\r[mdioo]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000CA00)) 
    \r[mdioo]_i_12 
       (.I0(\r[mdioo]_i_17_n_0 ),
        .I1(\r[mdioo]_i_18_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .O(\r[mdioo]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB800B8FF)) 
    \r[mdioo]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [0]),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I2(\r[mdioo]_i_19_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I4(\etho[mdio_o] ),
        .O(\r[mdioo]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F202F2F2F202020)) 
    \r[mdioo]_i_14 
       (.I0(\etho[mdc] ),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][phyadr_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I5(\r[mdioo]_i_20_n_0 ),
        .O(\r[mdioo]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000005700)) 
    \r[mdioo]_i_15 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/v[mdio_ctrl][write]1 ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I5(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .O(\m100.u0/ethc0/v[mdioo]5_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \r[mdioo]_i_16 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .O(\r[mdioo]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r[mdioo]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][11] ),
        .I1(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][10] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][9] ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/p_1_in128_in ),
        .O(\r[mdioo]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r[mdioo]_i_18 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][15] ),
        .I1(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][14] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][13] ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][12] ),
        .O(\r[mdioo]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r[mdioo]_i_19 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [1]),
        .I1(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [2]),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [3]),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][regadr]__0 [4]),
        .O(\r[mdioo]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F008F8F0F008080)) 
    \r[mdioo]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I1(\r[mdioo]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I3(\r_reg[mdioo]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I5(\r[mdioo]_i_6_n_0 ),
        .O(\r[mdioo]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r[mdioo]_i_20 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][phyadr_n_0_][1] ),
        .I1(\m100.u0/ethc0/data2 ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/data1 ),
        .I4(\m100.u0/ethc0/r_reg[cnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][phyadr_n_0_][4] ),
        .O(\r[mdioo]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \r[mdioo]_i_3 
       (.I0(\r[mdioo]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [3]),
        .I2(\r[mdioo]_i_8_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [2]),
        .I4(\r[mdioo]_i_9_n_0 ),
        .O(\m100.u0/ethc0/v[mdioo] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF11100100)) 
    \r[mdioo]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[cnt_n_0_][2] ),
        .I3(\r[mdioo]_i_10_n_0 ),
        .I4(\r[mdioo]_i_11_n_0 ),
        .I5(\r[mdioo]_i_12_n_0 ),
        .O(\r[mdioo]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88B8333388B80000)) 
    \r[mdioo]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I2(\etho[mdc] ),
        .I3(\m100.u0/ethc0/p_1_in143_in ),
        .I4(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][busy]__0 ),
        .O(\r[mdioo]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000202220)) 
    \r[mdioo]_i_7 
       (.I0(\etho[mdc] ),
        .I1(\m100.u0/ethc0/p_1_in143_in ),
        .I2(\m100.u0/ethc0/r_reg[mdio_ctrl][write]__0 ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I4(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I5(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .O(\r[mdioo]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30C030C074F330C0)) 
    \r[mdioo]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][read]__0 ),
        .I1(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I2(\m100.u0/ethc0/v[mdioo]5_out ),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I4(\etho[mdc] ),
        .I5(\m100.u0/ethc0/p_1_in143_in ),
        .O(\r[mdioo]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF8FFF8000000000)) 
    \r[mdioo]_i_9 
       (.I0(\r[mdioo]_i_16_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[cnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[mdio_state] [0]),
        .I3(\m100.u0/ethc0/r_reg[mdio_state] [1]),
        .I4(\m100.u0/ethc0/r_reg[mdio_ctrl][busy]__0 ),
        .I5(\m100.u0/ethc0/v[mdio_ctrl][write]1 ),
        .O(\r[mdioo]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[msbgood]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [21]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][37] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [22]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][38] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][39] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [23]),
        .O(\r[msbgood]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[msbgood]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [20]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][36] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [18]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][34] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][35] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [19]),
        .O(\r[msbgood]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[msbgood]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][33] ),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [17]),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [15]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][31] ),
        .I4(\m100.u0/ethc0/r_reg[checkdata]__0 [16]),
        .I5(\m100.u0/ethc0/r_reg[mac_addr_n_0_][32] ),
        .O(\r[msbgood]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[msbgood]_i_14 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [12]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][28] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [13]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][29] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][30] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [14]),
        .O(\r[msbgood]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[msbgood]_i_15 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [10]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][26] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [9]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][25] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][27] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [11]),
        .O(\r[msbgood]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[msbgood]_i_16 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [7]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][23] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [6]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][22] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][24] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [8]),
        .O(\r[msbgood]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[msbgood]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [5]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][21] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [3]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][19] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][20] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [4]),
        .O(\r[msbgood]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[msbgood]_i_18 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [0]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][16] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][17] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][18] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [2]),
        .O(\r[msbgood]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFD)) 
    \r[msbgood]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I2(\r[msbgood]_i_4_n_0 ),
        .O(\r[msbgood]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \r[msbgood]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .I1(\r[msbgood]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .O(\r[msbgood]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[msbgood]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[mac_addr_n_0_][47] ),
        .I1(\m100.u0/ethc0/r_reg[checkdata]__0 [31]),
        .I2(\m100.u0/ethc0/r_reg[mac_addr_n_0_][46] ),
        .I3(\m100.u0/ethc0/r_reg[checkdata]__0 [30]),
        .O(\r[msbgood]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[msbgood]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [27]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][43] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [28]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][44] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][45] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [29]),
        .O(\r[msbgood]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[msbgood]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[checkdata]__0 [24]),
        .I1(\m100.u0/ethc0/r_reg[mac_addr_n_0_][40] ),
        .I2(\m100.u0/ethc0/r_reg[checkdata]__0 [25]),
        .I3(\m100.u0/ethc0/r_reg[mac_addr_n_0_][41] ),
        .I4(\m100.u0/ethc0/r_reg[mac_addr_n_0_][42] ),
        .I5(\m100.u0/ethc0/r_reg[checkdata]__0 [26]),
        .O(\r[msbgood]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    \r[msbgood]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[check]__0 ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .O(\r[msbgood]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \r[nak]_i_1 
       (.I0(\m100.u0/ethc0/v[nak]1 ),
        .O(\r[nak]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[nak]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[seq] [13]),
        .I1(\m100.u0/rxwdata [31]),
        .I2(\m100.u0/ethc0/r_reg[seq] [12]),
        .I3(\m100.u0/rxwdata [30]),
        .O(\r[nak]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[nak]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[seq] [11]),
        .I1(\m100.u0/rxwdata [29]),
        .I2(\m100.u0/rxwdata [27]),
        .I3(\m100.u0/ethc0/r_reg[seq] [9]),
        .I4(\m100.u0/rxwdata [28]),
        .I5(\m100.u0/ethc0/r_reg[seq] [10]),
        .O(\r[nak]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[nak]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[seq] [8]),
        .I1(\m100.u0/rxwdata [26]),
        .I2(\m100.u0/rxwdata [25]),
        .I3(\m100.u0/ethc0/r_reg[seq] [7]),
        .I4(\m100.u0/rxwdata [24]),
        .I5(\m100.u0/ethc0/r_reg[seq] [6]),
        .O(\r[nak]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[nak]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[seq] [5]),
        .I1(\m100.u0/rxwdata [23]),
        .I2(\m100.u0/rxwdata [22]),
        .I3(\m100.u0/ethc0/r_reg[seq] [4]),
        .I4(\m100.u0/rxwdata [21]),
        .I5(\m100.u0/ethc0/r_reg[seq] [3]),
        .O(\r[nak]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[nak]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[seq] [0]),
        .I1(\m100.u0/rxwdata [18]),
        .I2(\m100.u0/rxwdata [20]),
        .I3(\m100.u0/ethc0/r_reg[seq] [2]),
        .I4(\m100.u0/rxwdata [19]),
        .I5(\m100.u0/ethc0/r_reg[seq] [1]),
        .O(\r[nak]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5545)) 
    \r[phywr]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I1(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I2(\m100.u0/ethc0/r_reg[rstaneg_n_0_] ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .O(\r[phywr]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000555400555554)) 
    \r[phywr]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[regaddr] [2]),
        .I1(\m100.u0/ethc0/r_reg[rstaneg_n_0_] ),
        .I2(\r[phywr]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[regaddr] [1]),
        .I4(\m100.u0/ethc0/r_reg[regaddr] [0]),
        .I5(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][0] ),
        .O(\m100.u0/ethc0/v[phywr] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0051)) 
    \r[phywr]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][12] ),
        .I1(\m100.u0/ethc0/r_reg[phywr]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rstaneg_n_0_] ),
        .I3(\m100.u0/ethc0/r_reg[mdio_ctrl][data_n_0_][15] ),
        .O(\r[phywr]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAEEEAAAA)) 
    \r[rcntl][0]_i_1 
       (.I0(\r[rcntl][0]_i_2_n_0 ),
        .I1(\r[rcntl][0]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\m100.u0/ethc0/v[rcntl] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4000555573114055)) 
    \r[rcntl][0]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\r[rcntl][0]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ewaddressl [0]),
        .O(\r[rcntl][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8888FFFF8C88FBFF)) 
    \r[rcntl][0]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I4(\m100.u0/ewaddressl [0]),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\r[rcntl][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000038CF)) 
    \r[rcntl][0]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/ewaddressl [0]),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\r[rcntl][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAEBFBFAEAEAEAEAE)) 
    \r[rcntl][1]_i_1 
       (.I0(\r[rcntl][1]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ewaddressl [1]),
        .I4(\m100.u0/ewaddressl [0]),
        .I5(\r[rcntl][1]_i_3_n_0 ),
        .O(\m100.u0/ethc0/v[rcntl] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40FF4000)) 
    \r[rcntl][1]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\r[rcntl][1]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I4(\r[rcntl][1]_i_5_n_0 ),
        .O(\r[rcntl][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[rcntl][1]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\r[rcntl][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h01FEFC0300FFFD02)) 
    \r[rcntl][1]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ewaddressl [1]),
        .I4(\m100.u0/ewaddressl [0]),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\r[rcntl][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB88B8BB88F8F8888)) 
    \r[rcntl][1]_i_5 
       (.I0(\r[rcntl][1]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ewaddressl [1]),
        .I3(\m100.u0/ewaddressl [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\r[rcntl][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1101221333130000)) 
    \r[rcntl][1]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I4(\m100.u0/ewaddressl [1]),
        .I5(\m100.u0/ewaddressl [0]),
        .O(\r[rcntl][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \r[rcntl][2]_i_1 
       (.I0(\r[rcntm][2]_i_2_n_0 ),
        .I1(\r[rcntl][2]_i_2_n_0 ),
        .I2(\r[rcntl][6]_i_8_n_0 ),
        .I3(\r[rcntl][2]_i_3_n_0 ),
        .I4(\r[rcntl][2]_i_4_n_0 ),
        .I5(\r[rcntl][6]_i_12_n_0 ),
        .O(\m100.u0/ethc0/v[rcntl] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF636900006369)) 
    \r[rcntl][2]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I1(\m100.u0/ewaddressl [2]),
        .I2(\m100.u0/ewaddressl [1]),
        .I3(\m100.u0/ewaddressl [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\r[rcntl][2]_i_5_n_0 ),
        .O(\r[rcntl][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    \r[rcntl][2]_i_3 
       (.I0(\m100.u0/ewaddressl [2]),
        .I1(\m100.u0/ewaddressl [0]),
        .I2(\m100.u0/ewaddressl [1]),
        .O(\r[rcntl][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h08F75FA0FF00F708)) 
    \r[rcntl][2]_i_4 
       (.I0(\r[rcntl][5]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/ewaddressl [2]),
        .I4(\m100.u0/ewaddressl [0]),
        .I5(\m100.u0/ewaddressl [1]),
        .O(\r[rcntl][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000051050000A2FB)) 
    \r[rcntl][2]_i_5 
       (.I0(\r[rcntl][2]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/ewaddressl [2]),
        .O(\r[rcntl][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[rcntl][2]_i_6 
       (.I0(\m100.u0/ewaddressl [1]),
        .I1(\m100.u0/ewaddressl [0]),
        .O(\r[rcntl][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEEEFEEEEEFEEE)) 
    \r[rcntl][3]_i_1 
       (.I0(\r[rcntl][3]_i_2_n_0 ),
        .I1(\r[rcntl][3]_i_3_n_0 ),
        .I2(\r[rcntl][3]_i_4_n_0 ),
        .I3(\m100.u0/ewaddressl [2]),
        .I4(\r[rcntl][3]_i_5_n_0 ),
        .I5(\m100.u0/ewaddressl [3]),
        .O(\m100.u0/ethc0/v[rcntl] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[rcntl][3]_i_10 
       (.I0(\m100.u0/ewaddressl [1]),
        .I1(\m100.u0/ewaddressl [2]),
        .O(\r[rcntl][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE00040F040F0E000)) 
    \r[rcntl][3]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\r[rcntl][3]_i_6_n_0 ),
        .I2(\r[rcntl][5]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\m100.u0/ewaddressl [2]),
        .I5(\m100.u0/ewaddressl [3]),
        .O(\r[rcntl][3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5454FCAC50500000)) 
    \r[rcntl][3]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\r[rcntl][3]_i_6_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\r[rcntl][3]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntl][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFA802)) 
    \r[rcntl][3]_i_3 
       (.I0(\r[rcntm][3]_i_8_n_0 ),
        .I1(\m100.u0/ewaddressl [1]),
        .I2(\m100.u0/ewaddressl [2]),
        .I3(\m100.u0/ewaddressl [3]),
        .I4(\r[rcntl][3]_i_8_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntl][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \r[rcntl][3]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\r[rcntl][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[rcntl][3]_i_5 
       (.I0(\m100.u0/ewaddressl [1]),
        .I1(\m100.u0/ewaddressl [0]),
        .O(\r[rcntl][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \r[rcntl][3]_i_6 
       (.I0(\m100.u0/ewaddressl [3]),
        .I1(\m100.u0/ewaddressl [0]),
        .I2(\m100.u0/ewaddressl [1]),
        .I3(\m100.u0/ewaddressl [2]),
        .O(\r[rcntl][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCECEECEC0FF0F0F0)) 
    \r[rcntl][3]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\r[rcntl][3]_i_9_n_0 ),
        .I2(\m100.u0/ewaddressl [3]),
        .I3(\m100.u0/ewaddressl [0]),
        .I4(\r[rcntl][3]_i_10_n_0 ),
        .I5(\r[rcntl][5]_i_5_n_0 ),
        .O(\r[rcntl][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF2F2F0F0F2220000)) 
    \r[rcntl][3]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\r[rcntl][5]_i_10_n_0 ),
        .I4(\r[rcntl][3]_i_6_n_0 ),
        .I5(\r[rcntl][3]_i_11_n_0 ),
        .O(\r[rcntl][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4444444114444444)) 
    \r[rcntl][3]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\m100.u0/ewaddressl [3]),
        .I2(\m100.u0/ewaddressl [2]),
        .I3(\m100.u0/ewaddressl [1]),
        .I4(\m100.u0/ewaddressl [0]),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\r[rcntl][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFAFAEEEEAAAA)) 
    \r[rcntl][4]_i_1 
       (.I0(\r[rcntl][4]_i_2_n_0 ),
        .I1(\r[rcntl][6]_i_8_n_0 ),
        .I2(\r[rcntl][4]_i_3_n_0 ),
        .I3(\r[rcntl][6]_i_10_n_0 ),
        .I4(\r[rcntl][4]_i_4_n_0 ),
        .I5(\r[rcntl][6]_i_12_n_0 ),
        .O(\m100.u0/ethc0/v[rcntl] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44444000)) 
    \r[rcntl][4]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\r[rcntl][4]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\r[rcntl][4]_i_6_n_0 ),
        .O(\r[rcntl][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0020A88888A82000)) 
    \r[rcntl][4]_i_3 
       (.I0(\r[rcntl][5]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\r[rcntl][5]_i_8_n_0 ),
        .I4(\m100.u0/ewaddressl [4]),
        .I5(\r[rcntl][5]_i_7_n_0 ),
        .O(\r[rcntl][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \r[rcntl][4]_i_4 
       (.I0(\m100.u0/ewaddressl [4]),
        .I1(\m100.u0/ewaddressl [1]),
        .I2(\m100.u0/ewaddressl [0]),
        .I3(\m100.u0/ewaddressl [3]),
        .I4(\m100.u0/ewaddressl [2]),
        .O(\r[rcntl][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF0FF20230000)) 
    \r[rcntl][4]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\r[rcntl][4]_i_4_n_0 ),
        .I5(\r[rcntl][4]_i_7_n_0 ),
        .O(\r[rcntl][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1320102313201320)) 
    \r[rcntl][4]_i_6 
       (.I0(\r[rcntl][4]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ewaddressl [4]),
        .I4(\m100.u0/ewaddressl [3]),
        .I5(\r[rcntl][4]_i_9_n_0 ),
        .O(\r[rcntl][4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC4C4C44C0CC0C0C0)) 
    \r[rcntl][4]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\r[rcntl][5]_i_5_n_0 ),
        .I2(\m100.u0/ewaddressl [4]),
        .I3(\m100.u0/ewaddressl [2]),
        .I4(\m100.u0/ewaddressl [3]),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\r[rcntl][4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8880)) 
    \r[rcntl][4]_i_8 
       (.I0(\m100.u0/ewaddressl [2]),
        .I1(\m100.u0/ewaddressl [3]),
        .I2(\m100.u0/ewaddressl [0]),
        .I3(\m100.u0/ewaddressl [1]),
        .O(\r[rcntl][4]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[rcntl][4]_i_9 
       (.I0(\m100.u0/ewaddressl [1]),
        .I1(\m100.u0/ewaddressl [2]),
        .O(\r[rcntl][4]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBAFFBABAAAAAAAAA)) 
    \r[rcntl][5]_i_1 
       (.I0(\r[rcntl][5]_i_2_n_0 ),
        .I1(\r[rcntl][6]_i_10_n_0 ),
        .I2(\r[rcntl][5]_i_3_n_0 ),
        .I3(\r[rcntl][5]_i_4_n_0 ),
        .I4(\r[rcntl][5]_i_5_n_0 ),
        .I5(\r[rcntl][6]_i_12_n_0 ),
        .O(\m100.u0/ethc0/v[rcntl] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00D1)) 
    \r[rcntl][5]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\r[rcntl][5]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h70D070D000F0F000)) 
    \r[rcntl][5]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\r[rcntl][5]_i_13_n_0 ),
        .I2(\r[rcntl][5]_i_5_n_0 ),
        .I3(\m100.u0/ewaddressl [5]),
        .I4(\r[rcntl][5]_i_14_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\r[rcntl][5]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \r[rcntl][5]_i_12 
       (.I0(\m100.u0/ewaddressl [2]),
        .I1(\m100.u0/ewaddressl [1]),
        .I2(\m100.u0/ewaddressl [3]),
        .O(\r[rcntl][5]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \r[rcntl][5]_i_13 
       (.I0(\m100.u0/ewaddressl [2]),
        .I1(\m100.u0/ewaddressl [3]),
        .I2(\m100.u0/ewaddressl [4]),
        .O(\r[rcntl][5]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \r[rcntl][5]_i_14 
       (.I0(\m100.u0/ewaddressl [2]),
        .I1(\m100.u0/ewaddressl [3]),
        .I2(\m100.u0/ewaddressl [4]),
        .O(\r[rcntl][5]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h02020202FF000808)) 
    \r[rcntl][5]_i_2 
       (.I0(\r[rcntl][5]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\r[rcntl][5]_i_6_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntl][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    \r[rcntl][5]_i_3 
       (.I0(\m100.u0/ewaddressl [5]),
        .I1(\m100.u0/ewaddressl [1]),
        .I2(\m100.u0/ewaddressl [0]),
        .I3(\m100.u0/ewaddressl [2]),
        .I4(\m100.u0/ewaddressl [3]),
        .I5(\m100.u0/ewaddressl [4]),
        .O(\r[rcntl][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h939393933C33FFFF)) 
    \r[rcntl][5]_i_4 
       (.I0(\r[rcntl][5]_i_7_n_0 ),
        .I1(\m100.u0/ewaddressl [5]),
        .I2(\m100.u0/ewaddressl [4]),
        .I3(\r[rcntl][5]_i_8_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\r[rcntl][5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[rcntl][5]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .O(\r[rcntl][5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEAAEEEAEAAAAA)) 
    \r[rcntl][5]_i_6 
       (.I0(\r[rcntl][5]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\r[rcntl][5]_i_10_n_0 ),
        .I3(\FSM_sequential_r[edclrstate][3]_i_20_n_0 ),
        .I4(\r[rcntl][5]_i_3_n_0 ),
        .I5(\r[rcntl][5]_i_11_n_0 ),
        .O(\r[rcntl][5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \r[rcntl][5]_i_7 
       (.I0(\m100.u0/ewaddressl [2]),
        .I1(\m100.u0/ewaddressl [1]),
        .I2(\m100.u0/ewaddressl [3]),
        .O(\r[rcntl][5]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \r[rcntl][5]_i_8 
       (.I0(\m100.u0/ewaddressl [0]),
        .I1(\m100.u0/ewaddressl [1]),
        .I2(\m100.u0/ewaddressl [2]),
        .I3(\m100.u0/ewaddressl [3]),
        .O(\r[rcntl][5]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1320300313203300)) 
    \r[rcntl][5]_i_9 
       (.I0(\r[rcntl][4]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ewaddressl [5]),
        .I4(\m100.u0/ewaddressl [4]),
        .I5(\r[rcntl][5]_i_12_n_0 ),
        .O(\r[rcntl][5]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF2F000000)) 
    \r[rcntl][6]_i_1 
       (.I0(\r[rcntl][6]_i_3_n_0 ),
        .I1(\r[rcntl][6]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\r[rcntl][6]_i_5_n_0 ),
        .I5(\r[rcntl][6]_i_6_n_0 ),
        .O(\r[rcntl][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1110)) 
    \r[rcntl][6]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\r[rcntl][6]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \r[rcntl][6]_i_11 
       (.I0(\m100.u0/ewaddressl [6]),
        .I1(\m100.u0/ewaddressl [1]),
        .I2(\m100.u0/ewaddressl [0]),
        .I3(\r[rcntl][6]_i_18_n_0 ),
        .O(\r[rcntl][6]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \r[rcntl][6]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntl][6]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000888B8B88)) 
    \r[rcntl][6]_i_13 
       (.I0(\m100.u0/ethc0/v[writeok]1 ),
        .I1(\r[erxidle]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/p_6_in [14]),
        .I3(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I4(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntl][6]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2800222228008888)) 
    \r[rcntl][6]_i_14 
       (.I0(\r[rcntl][5]_i_5_n_0 ),
        .I1(\m100.u0/ewaddressl [6]),
        .I2(\r[rcntl][6]_i_19_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I5(\r[rcntl][6]_i_18_n_0 ),
        .O(\r[rcntl][6]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBEBA)) 
    \r[rcntl][6]_i_15 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\r[rcntl][6]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1320102313201320)) 
    \r[rcntl][6]_i_16 
       (.I0(\r[rcntl][6]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ewaddressl [6]),
        .I4(\m100.u0/ewaddressl [1]),
        .I5(\r[rcntl][6]_i_19_n_0 ),
        .O(\r[rcntl][6]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4440444400040000)) 
    \r[rcntl][6]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ewaddressl [0]),
        .I3(\m100.u0/ewaddressl [1]),
        .I4(\r[rcntl][6]_i_19_n_0 ),
        .I5(\m100.u0/ewaddressl [6]),
        .O(\r[rcntl][6]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \r[rcntl][6]_i_18 
       (.I0(\m100.u0/ewaddressl [4]),
        .I1(\m100.u0/ewaddressl [3]),
        .I2(\m100.u0/ewaddressl [2]),
        .I3(\m100.u0/ewaddressl [5]),
        .O(\r[rcntl][6]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \r[rcntl][6]_i_19 
       (.I0(\m100.u0/ewaddressl [4]),
        .I1(\m100.u0/ewaddressl [3]),
        .I2(\m100.u0/ewaddressl [2]),
        .I3(\m100.u0/ewaddressl [5]),
        .O(\r[rcntl][6]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFAFAEEEEAAAA)) 
    \r[rcntl][6]_i_2 
       (.I0(\r[rcntl][6]_i_7_n_0 ),
        .I1(\r[rcntl][6]_i_8_n_0 ),
        .I2(\r[rcntl][6]_i_9_n_0 ),
        .I3(\r[rcntl][6]_i_10_n_0 ),
        .I4(\r[rcntl][6]_i_11_n_0 ),
        .I5(\r[rcntl][6]_i_12_n_0 ),
        .O(\m100.u0/ethc0/v[rcntl] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000800080000000)) 
    \r[rcntl][6]_i_20 
       (.I0(\m100.u0/ewaddressl [5]),
        .I1(\m100.u0/ewaddressl [2]),
        .I2(\m100.u0/ewaddressl [3]),
        .I3(\m100.u0/ewaddressl [4]),
        .I4(\m100.u0/ewaddressl [0]),
        .I5(\m100.u0/ewaddressl [1]),
        .O(\r[rcntl][6]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \r[rcntl][6]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I1(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\r[rcntl][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \r[rcntl][6]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\r[rcntl][6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[rcntl][6]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntl][6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFAAEAAA)) 
    \r[rcntl][6]_i_6 
       (.I0(\r[rcntl][6]_i_13_n_0 ),
        .I1(\m100.u0/ethc0/v[rcntm]0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I4(\r[rcntm][6]_i_4_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\r[rcntl][6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA88A80000)) 
    \r[rcntl][6]_i_7 
       (.I0(\r[rcntm][2]_i_2_n_0 ),
        .I1(\r[rcntl][6]_i_14_n_0 ),
        .I2(\r[rcntl][6]_i_11_n_0 ),
        .I3(\r[rcntl][6]_i_15_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\r[rcntl][6]_i_16_n_0 ),
        .O(\r[rcntl][6]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0034)) 
    \r[rcntl][6]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\r[rcntl][6]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8AAAA88888888888)) 
    \r[rcntl][6]_i_9 
       (.I0(\r[rcntl][5]_i_5_n_0 ),
        .I1(\r[rcntl][6]_i_17_n_0 ),
        .I2(\r[rcntl][6]_i_18_n_0 ),
        .I3(\m100.u0/ewaddressl [1]),
        .I4(\m100.u0/ewaddressl [6]),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\r[rcntl][6]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAEAEAEAEEEAEAEA)) 
    \r[rcntm][0]_i_1 
       (.I0(\r[rcntm][0]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\r[rcntm][0]_i_3_n_0 ),
        .I3(\r[rcntm][0]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\m100.u0/ethc0/v[rcntm] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h080B0000040400CC)) 
    \r[rcntm][0]_i_2 
       (.I0(\r[rcntm][0]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ewaddressm [0]),
        .O(\r[rcntm][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555000044447337)) 
    \r[rcntm][0]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[rxdone] ),
        .I3(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ewaddressm [0]),
        .O(\r[rcntm][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11012156)) 
    \r[rcntm][0]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ewaddressm [0]),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .O(\r[rcntm][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0110)) 
    \r[rcntm][0]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\r[rcntm][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAEAEFEAE)) 
    \r[rcntm][1]_i_1 
       (.I0(\r[rcntm][1]_i_2_n_0 ),
        .I1(\r[rcntm][1]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\r[rcntm][1]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\m100.u0/ethc0/v[rcntm] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FA004400AA0044)) 
    \r[rcntm][1]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\r[rcntm][1]_i_5_n_0 ),
        .I2(\r[rcntm][1]_i_6_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntm][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F807FB043807FB)) 
    \r[rcntm][1]_i_3 
       (.I0(\m100.u0/ewaddressm [0]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ewaddressm [1]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\r[rcntm][1]_i_7_n_0 ),
        .O(\r[rcntm][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0440444444440440)) 
    \r[rcntm][1]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\m100.u0/ewaddressm [0]),
        .I3(\m100.u0/ewaddressm [1]),
        .I4(\m100.u0/ethc0/r_reg[rxdone] ),
        .I5(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\r[rcntm][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[rcntm][1]_i_5 
       (.I0(\m100.u0/ewaddressm [0]),
        .I1(\m100.u0/ewaddressm [1]),
        .O(\r[rcntm][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6666666669666556)) 
    \r[rcntm][1]_i_6 
       (.I0(\m100.u0/ewaddressm [1]),
        .I1(\m100.u0/ewaddressm [0]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\r[rcntm][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F0F0A060006060A)) 
    \r[rcntm][1]_i_7 
       (.I0(\m100.u0/ewaddressm [1]),
        .I1(\m100.u0/ewaddressm [0]),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\r[rcntm][1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF8F8F888)) 
    \r[rcntm][2]_i_1 
       (.I0(\r[rcntm][2]_i_2_n_0 ),
        .I1(\r[rcntm][2]_i_3_n_0 ),
        .I2(\r[rcntm][6]_i_10_n_0 ),
        .I3(\r[rcntm][2]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/v[rxstatus]2 ),
        .I5(\r[rcntm][2]_i_5_n_0 ),
        .O(\m100.u0/ethc0/v[rcntm] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \r[rcntm][2]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\r[rcntm][2]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFDF)) 
    \r[rcntm][2]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\r[rcntm][2]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[rcntm][2]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntm][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF3C7800003C78)) 
    \r[rcntm][2]_i_3 
       (.I0(\m100.u0/ewaddressm [0]),
        .I1(\m100.u0/ewaddressm [1]),
        .I2(\m100.u0/ewaddressm [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\r[rcntm][2]_i_6_n_0 ),
        .O(\r[rcntm][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    \r[rcntm][2]_i_4 
       (.I0(\m100.u0/ewaddressm [2]),
        .I1(\m100.u0/ewaddressm [1]),
        .I2(\m100.u0/ewaddressm [0]),
        .O(\r[rcntm][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h445444444444FF44)) 
    \r[rcntm][2]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\r[rcntm][2]_i_7_n_0 ),
        .I2(\r[rcntm][2]_i_8_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntm][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0005544800055E4D)) 
    \r[rcntm][2]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\r[rcntm][2]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/ewaddressm [2]),
        .O(\r[rcntm][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000787800C30000)) 
    \r[rcntm][2]_i_7 
       (.I0(\m100.u0/ewaddressm [0]),
        .I1(\m100.u0/ewaddressm [1]),
        .I2(\m100.u0/ewaddressm [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntm][2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFEBB0000)) 
    \r[rcntm][2]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\r[rcntm][2]_i_4_n_0 ),
        .I5(\r[rcntm][2]_i_9_n_0 ),
        .O(\r[rcntm][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F444F000F44440F)) 
    \r[rcntm][2]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\r[rcntm][2]_i_10_n_0 ),
        .I2(\r[rcntm][2]_i_11_n_0 ),
        .I3(\m100.u0/ewaddressm [2]),
        .I4(\m100.u0/ewaddressm [1]),
        .I5(\m100.u0/ewaddressm [0]),
        .O(\r[rcntm][2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF2E0C2A00)) 
    \r[rcntm][3]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I3(\r[rcntm][3]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\r[rcntm][3]_i_3_n_0 ),
        .O(\m100.u0/ethc0/v[rcntm] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \r[rcntm][3]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\r[rcntm][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0155)) 
    \r[rcntm][3]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .O(\r[rcntm][3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \r[rcntm][3]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\r[rcntm][3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000074000030E2)) 
    \r[rcntm][3]_i_13 
       (.I0(\r[rcntm][3]_i_15_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\r[rcntm][3]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\r[rcntm][3]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[rcntm][3]_i_14 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\r[rcntm][3]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[rcntm][3]_i_15 
       (.I0(\m100.u0/ewaddressm [2]),
        .I1(\m100.u0/ewaddressm [3]),
        .O(\r[rcntm][3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF82AAFF0082AA)) 
    \r[rcntm][3]_i_2 
       (.I0(\r[rcntm][3]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdone] ),
        .I2(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\r[rcntm][3]_i_5_n_0 ),
        .O(\r[rcntm][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F8F8F888F888F88)) 
    \r[rcntm][3]_i_3 
       (.I0(\r[rcntm][3]_i_6_n_0 ),
        .I1(\r[rcntl][3]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\r[rcntm][3]_i_7_n_0 ),
        .I4(\r[rcntm][3]_i_4_n_0 ),
        .I5(\r[rcntm][3]_i_8_n_0 ),
        .O(\r[rcntm][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \r[rcntm][3]_i_4 
       (.I0(\m100.u0/ewaddressm [3]),
        .I1(\m100.u0/ewaddressm [2]),
        .I2(\m100.u0/ewaddressm [0]),
        .I3(\m100.u0/ewaddressm [1]),
        .O(\r[rcntm][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF444F444FFFFF444)) 
    \r[rcntm][3]_i_5 
       (.I0(\r[rcntm][3]_i_9_n_0 ),
        .I1(\r[rcntl][5]_i_5_n_0 ),
        .I2(\r[rcntm][3]_i_10_n_0 ),
        .I3(\r[rcntm][3]_i_6_n_0 ),
        .I4(\r[rcntm][3]_i_4_n_0 ),
        .I5(\r[rcntm][3]_i_11_n_0 ),
        .O(\r[rcntm][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    \r[rcntm][3]_i_6 
       (.I0(\m100.u0/ewaddressm [3]),
        .I1(\m100.u0/ewaddressm [2]),
        .I2(\m100.u0/ewaddressm [1]),
        .O(\r[rcntm][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F4F44F44444444)) 
    \r[rcntm][3]_i_7 
       (.I0(\r[rcntm][3]_i_12_n_0 ),
        .I1(\r[rcntm][3]_i_13_n_0 ),
        .I2(\m100.u0/ewaddressm [3]),
        .I3(\m100.u0/ewaddressm [2]),
        .I4(\m100.u0/ewaddressm [1]),
        .I5(\r[rcntm][3]_i_14_n_0 ),
        .O(\r[rcntm][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[rcntm][3]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .O(\r[rcntm][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h704000088FBFFFF7)) 
    \r[rcntm][3]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ewaddressm [1]),
        .I3(\m100.u0/ewaddressm [0]),
        .I4(\m100.u0/ewaddressm [2]),
        .I5(\m100.u0/ewaddressm [3]),
        .O(\r[rcntm][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF2F2FFF2F2F2F2F2)) 
    \r[rcntm][4]_i_1 
       (.I0(\r[rcntm][4]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\r[rcntm][4]_i_3_n_0 ),
        .I3(\r[rcntm][4]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/v[rxstatus]2 ),
        .I5(\r[rcntm][6]_i_10_n_0 ),
        .O(\m100.u0/ethc0/v[rcntm] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3F0F0F0F0F0F0B4)) 
    \r[rcntm][4]_i_10 
       (.I0(\m100.u0/ewaddressm [0]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\m100.u0/ewaddressm [4]),
        .I3(\m100.u0/ewaddressm [2]),
        .I4(\m100.u0/ewaddressm [3]),
        .I5(\m100.u0/ewaddressm [1]),
        .O(\r[rcntm][4]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h008A00208A882022)) 
    \r[rcntm][4]_i_11 
       (.I0(\r[rcntm][6]_i_28_n_0 ),
        .I1(\r[rcntm][5]_i_13_n_0 ),
        .I2(\r[rcntm][6]_i_21_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ewaddressm [4]),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\r[rcntm][4]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r[rcntm][4]_i_12 
       (.I0(\m100.u0/ewaddressm [2]),
        .I1(\m100.u0/ewaddressm [3]),
        .O(\r[rcntm][4]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFAFFFAEAEAEAEAEA)) 
    \r[rcntm][4]_i_2 
       (.I0(\r[rcntm][4]_i_5_n_0 ),
        .I1(\r[rcntl][1]_i_3_n_0 ),
        .I2(\r[rcntm][4]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I4(\r[rcntm][4]_i_6_n_0 ),
        .I5(\r[rcntm][6]_i_18_n_0 ),
        .O(\r[rcntm][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8A808A8A8A808080)) 
    \r[rcntm][4]_i_3 
       (.I0(\r[rcntm][2]_i_2_n_0 ),
        .I1(\r[rcntm][4]_i_7_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\r[rcntm][4]_i_8_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\r[rcntm][4]_i_4_n_0 ),
        .O(\r[rcntm][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \r[rcntm][4]_i_4 
       (.I0(\m100.u0/ewaddressm [4]),
        .I1(\m100.u0/ewaddressm [2]),
        .I2(\m100.u0/ewaddressm [3]),
        .I3(\m100.u0/ewaddressm [0]),
        .I4(\m100.u0/ewaddressm [1]),
        .O(\r[rcntm][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4444444000000004)) 
    \r[rcntm][4]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\r[rcntm][4]_i_9_n_0 ),
        .I2(\m100.u0/ewaddressm [1]),
        .I3(\m100.u0/ewaddressm [3]),
        .I4(\m100.u0/ewaddressm [2]),
        .I5(\m100.u0/ewaddressm [4]),
        .O(\r[rcntm][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF0EFEF0F004040)) 
    \r[rcntm][4]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\r[rcntm][4]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\r[rcntm][4]_i_10_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I5(\r[rcntm][4]_i_4_n_0 ),
        .O(\r[rcntm][4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAAEEEEEEAAEAAAA)) 
    \r[rcntm][4]_i_7 
       (.I0(\r[rcntm][4]_i_11_n_0 ),
        .I1(\r[rcntm][6]_i_27_n_0 ),
        .I2(\m100.u0/ewaddressm [4]),
        .I3(\r[rcntm][4]_i_12_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I5(\r[rcntm][4]_i_4_n_0 ),
        .O(\r[rcntm][4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \r[rcntm][4]_i_8 
       (.I0(\m100.u0/ewaddressm [4]),
        .I1(\m100.u0/ewaddressm [2]),
        .I2(\m100.u0/ewaddressm [3]),
        .I3(\m100.u0/ewaddressm [1]),
        .O(\r[rcntm][4]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[rcntm][4]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\r[rcntm][4]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF2F2FFF2F2F2F2F2)) 
    \r[rcntm][5]_i_1 
       (.I0(\r[rcntm][5]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\r[rcntm][5]_i_3_n_0 ),
        .I3(\r[rcntm][5]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/v[rxstatus]2 ),
        .I5(\r[rcntm][6]_i_10_n_0 ),
        .O(\m100.u0/ethc0/v[rcntm] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF2FEF000020200)) 
    \r[rcntm][5]_i_10 
       (.I0(\r[rcntm][5]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I5(\r[rcntm][5]_i_4_n_0 ),
        .O(\r[rcntm][5]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3333333C55555555)) 
    \r[rcntm][5]_i_11 
       (.I0(\r[rcntm][5]_i_4_n_0 ),
        .I1(\m100.u0/ewaddressm [5]),
        .I2(\m100.u0/ewaddressm [2]),
        .I3(\m100.u0/ewaddressm [3]),
        .I4(\m100.u0/ewaddressm [4]),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\r[rcntm][5]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDEDDDDD55A65555)) 
    \r[rcntm][5]_i_12 
       (.I0(\m100.u0/ewaddressm [5]),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I2(\r[rcntm][6]_i_21_n_0 ),
        .I3(\r[rcntm][5]_i_13_n_0 ),
        .I4(\m100.u0/ewaddressm [4]),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\r[rcntm][5]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \r[rcntm][5]_i_13 
       (.I0(\m100.u0/ewaddressm [2]),
        .I1(\m100.u0/ewaddressm [3]),
        .O(\r[rcntm][5]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00F0CCCC00AA0000)) 
    \r[rcntm][5]_i_2 
       (.I0(\r[rcntm][5]_i_5_n_0 ),
        .I1(\r[rcntm][5]_i_4_n_0 ),
        .I2(\r[rcntm][5]_i_6_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntm][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88A888AA88A88888)) 
    \r[rcntm][5]_i_3 
       (.I0(\r[rcntm][2]_i_2_n_0 ),
        .I1(\r[rcntm][5]_i_7_n_0 ),
        .I2(\r[rcntm][5]_i_8_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\r[rcntm][5]_i_4_n_0 ),
        .O(\r[rcntm][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    \r[rcntm][5]_i_4 
       (.I0(\m100.u0/ewaddressm [5]),
        .I1(\m100.u0/ewaddressm [4]),
        .I2(\m100.u0/ewaddressm [1]),
        .I3(\m100.u0/ewaddressm [0]),
        .I4(\m100.u0/ewaddressm [3]),
        .I5(\m100.u0/ewaddressm [2]),
        .O(\r[rcntm][5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAAAA9)) 
    \r[rcntm][5]_i_5 
       (.I0(\m100.u0/ewaddressm [5]),
        .I1(\m100.u0/ewaddressm [4]),
        .I2(\m100.u0/ewaddressm [1]),
        .I3(\m100.u0/ewaddressm [3]),
        .I4(\m100.u0/ewaddressm [2]),
        .O(\r[rcntm][5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF30AA0000)) 
    \r[rcntm][5]_i_6 
       (.I0(\r[rcntm][5]_i_4_n_0 ),
        .I1(\r[rcntm][5]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\r[rcntl][5]_i_5_n_0 ),
        .I5(\r[rcntm][5]_i_10_n_0 ),
        .O(\r[rcntm][5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0002111300000000)) 
    \r[rcntm][5]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\r[rcntm][5]_i_11_n_0 ),
        .I4(\r[rcntm][5]_i_12_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\r[rcntm][5]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \r[rcntm][5]_i_8 
       (.I0(\m100.u0/ewaddressm [5]),
        .I1(\m100.u0/ewaddressm [3]),
        .I2(\m100.u0/ewaddressm [2]),
        .I3(\m100.u0/ewaddressm [4]),
        .I4(\m100.u0/ewaddressm [1]),
        .O(\r[rcntm][5]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555555555555556)) 
    \r[rcntm][5]_i_9 
       (.I0(\m100.u0/ewaddressm [5]),
        .I1(\m100.u0/ewaddressm [1]),
        .I2(\m100.u0/ewaddressm [0]),
        .I3(\m100.u0/ewaddressm [3]),
        .I4(\m100.u0/ewaddressm [2]),
        .I5(\m100.u0/ewaddressm [4]),
        .O(\r[rcntm][5]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF2E22)) 
    \r[rcntm][6]_i_1 
       (.I0(\r[rcntm][6]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\r[rcntm][6]_i_4_n_0 ),
        .I4(\r[rcntm][6]_i_5_n_0 ),
        .O(\r[rcntm][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \r[rcntm][6]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\r[rcntm][6]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h140014141414143C)) 
    \r[rcntm][6]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I2(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .O(\r[rcntm][6]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[rcntm][6]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .O(\r[rcntm][6]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000007000700000)) 
    \r[rcntm][6]_i_13 
       (.I0(\r[rcntm][6]_i_22_n_0 ),
        .I1(\m100.u0/ewaddressm [6]),
        .I2(\m100.u0/ethc0/r_reg[ewr]__0 ),
        .I3(\m100.u0/ethc0/r_reg[nak_n_0_] ),
        .I4(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I5(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .O(\m100.u0/ethc0/v[rcntm]0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF88FF8F888888888)) 
    \r[rcntm][6]_i_14 
       (.I0(\r[rcntm][6]_i_8_n_0 ),
        .I1(\r[rcntl][1]_i_3_n_0 ),
        .I2(\m100.u0/ewaddressm [6]),
        .I3(\m100.u0/ewaddressm [1]),
        .I4(\r[rcntm][6]_i_23_n_0 ),
        .I5(\r[rcntm][6]_i_24_n_0 ),
        .O(\r[rcntm][6]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FD010000)) 
    \r[rcntm][6]_i_15 
       (.I0(\r[rcntm][6]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I3(\r[rcntm][6]_i_8_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\r[rcntm][6]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AA00AA00AA0C)) 
    \r[rcntm][6]_i_16 
       (.I0(\r[rcntm][6]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I5(\r[rcntm][6]_i_20_n_0 ),
        .O(\r[rcntm][6]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h333CFFFF55555555)) 
    \r[rcntm][6]_i_17 
       (.I0(\r[rcntm][6]_i_8_n_0 ),
        .I1(\m100.u0/ewaddressm [6]),
        .I2(\r[rcntm][6]_i_25_n_0 ),
        .I3(\m100.u0/ewaddressm [5]),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .O(\r[rcntm][6]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \r[rcntm][6]_i_18 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntm][6]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAEEAEEEEAEEAAAAA)) 
    \r[rcntm][6]_i_19 
       (.I0(\r[rcntm][6]_i_26_n_0 ),
        .I1(\r[rcntm][6]_i_27_n_0 ),
        .I2(\m100.u0/ewaddressm [6]),
        .I3(\r[rcntm][6]_i_23_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I5(\r[rcntm][6]_i_8_n_0 ),
        .O(\r[rcntm][6]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF2F2FFF2F2F2F2F2)) 
    \r[rcntm][6]_i_2 
       (.I0(\r[rcntm][6]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\r[rcntm][6]_i_7_n_0 ),
        .I3(\r[rcntm][6]_i_8_n_0 ),
        .I4(\m100.u0/ethc0/v[rxstatus]2 ),
        .I5(\r[rcntm][6]_i_10_n_0 ),
        .O(\m100.u0/ethc0/v[rcntm] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9555555555555555)) 
    \r[rcntm][6]_i_20 
       (.I0(\m100.u0/ewaddressm [6]),
        .I1(\m100.u0/ewaddressm [4]),
        .I2(\m100.u0/ewaddressm [2]),
        .I3(\m100.u0/ewaddressm [3]),
        .I4(\m100.u0/ewaddressm [5]),
        .I5(\m100.u0/ewaddressm [1]),
        .O(\r[rcntm][6]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[rcntm][6]_i_21 
       (.I0(\m100.u0/ewaddressm [0]),
        .I1(\m100.u0/ewaddressm [1]),
        .O(\r[rcntm][6]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \r[rcntm][6]_i_22 
       (.I0(\m100.u0/ewaddressm [1]),
        .I1(\m100.u0/ewaddressm [0]),
        .I2(\m100.u0/ewaddressm [5]),
        .I3(\m100.u0/ewaddressm [3]),
        .I4(\m100.u0/ewaddressm [2]),
        .I5(\m100.u0/ewaddressm [4]),
        .O(\r[rcntm][6]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \r[rcntm][6]_i_23 
       (.I0(\m100.u0/ewaddressm [2]),
        .I1(\m100.u0/ewaddressm [3]),
        .I2(\m100.u0/ewaddressm [4]),
        .I3(\m100.u0/ewaddressm [5]),
        .O(\r[rcntm][6]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \r[rcntm][6]_i_24 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[rcntm][6]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \r[rcntm][6]_i_25 
       (.I0(\m100.u0/ewaddressm [4]),
        .I1(\m100.u0/ewaddressm [2]),
        .I2(\m100.u0/ewaddressm [3]),
        .I3(\m100.u0/ewaddressm [0]),
        .I4(\m100.u0/ewaddressm [1]),
        .O(\r[rcntm][6]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h088A08800880088A)) 
    \r[rcntm][6]_i_26 
       (.I0(\r[rcntm][6]_i_28_n_0 ),
        .I1(\r[rcntm][6]_i_8_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I4(\r[rcntm][6]_i_29_n_0 ),
        .I5(\m100.u0/ewaddressm [6]),
        .O(\r[rcntm][6]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \r[rcntm][6]_i_27 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\r[rcntm][6]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[rcntm][6]_i_28 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .O(\r[rcntm][6]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \r[rcntm][6]_i_29 
       (.I0(\m100.u0/ewaddressm [4]),
        .I1(\m100.u0/ewaddressm [2]),
        .I2(\m100.u0/ewaddressm [3]),
        .I3(\m100.u0/ewaddressm [5]),
        .O(\r[rcntm][6]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAF0FA000FFFCF0FC)) 
    \r[rcntm][6]_i_3 
       (.I0(\r[rcntm][6]_i_11_n_0 ),
        .I1(\m100.u0/ethc0/v[edclrstate]0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\m100.u0/ethc0/v[writeok]1 ),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\r[rcntm][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF7500FFFF000000)) 
    \r[rcntm][6]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .I2(\r[rcntm][6]_i_12_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\m100.u0/ethc0/v[writeok]1 ),
        .O(\r[rcntm][6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F60000000000)) 
    \r[rcntm][6]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdone] ),
        .I2(\m100.u0/ethc0/v[rcntm]0 ),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\r[rcntm][6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFFFEAAAAAAAA)) 
    \r[rcntm][6]_i_6 
       (.I0(\r[rcntm][6]_i_14_n_0 ),
        .I1(\r[rcntm][6]_i_15_n_0 ),
        .I2(\r[rcntm][6]_i_16_n_0 ),
        .I3(\r[rcntl][5]_i_5_n_0 ),
        .I4(\r[rcntm][6]_i_17_n_0 ),
        .I5(\r[rcntm][6]_i_18_n_0 ),
        .O(\r[rcntm][6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h808A8A8A808A8080)) 
    \r[rcntm][6]_i_7 
       (.I0(\r[rcntm][2]_i_2_n_0 ),
        .I1(\r[rcntm][6]_i_19_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I3(\r[rcntm][6]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I5(\r[rcntm][6]_i_8_n_0 ),
        .O(\r[rcntm][6]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    \r[rcntm][6]_i_8 
       (.I0(\m100.u0/ewaddressm [6]),
        .I1(\m100.u0/ewaddressm [4]),
        .I2(\m100.u0/ewaddressm [2]),
        .I3(\m100.u0/ewaddressm [3]),
        .I4(\m100.u0/ewaddressm [5]),
        .I5(\r[rcntm][6]_i_21_n_0 ),
        .O(\r[rcntm][6]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[rcntm][6]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[rxdone] ),
        .I1(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\m100.u0/ethc0/v[rxstatus]2 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \r[retry]_i_1 
       (.I0(\m100.u0/ethc0/ahb0/r_reg ),
        .I1(\ahbmi[hresp] [1]),
        .I2(\ahbmi[hready] ),
        .O(\r[retry]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT4 #(
    .INIT(16'hA99A)) 
    \r[rfcnt][0]_i_1 
       (.I0(\m100.u0/ethc0/v[rfcnt] [0]),
        .I1(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I3(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .O(\m100.u0/ethc0/v[rfcnt]__0 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT5 #(
    .INIT(32'hAA96AAAA)) 
    \r[rfcnt][1]_i_1 
       (.I0(\m100.u0/ethc0/v[rfcnt] [1]),
        .I1(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I2(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I3(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/v[rfcnt] [0]),
        .O(\m100.u0/ethc0/v[rfcnt]__0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAA6A6AAAAAAAAAA)) 
    \r[rfcnt][2]_i_1 
       (.I0(\m100.u0/ethc0/v[rfcnt] [2]),
        .I1(\m100.u0/ethc0/v[rfcnt] [0]),
        .I2(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I4(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I5(\m100.u0/ethc0/v[rfcnt] [1]),
        .O(\m100.u0/ethc0/v[rfcnt]__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFFFFFF40000000)) 
    \r[rfcnt][2]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[rfcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/rmsti[ready] ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rfcnt_n_0_][1] ),
        .O(\r[rfcnt][2]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[rfcnt][2]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[rfcnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[rfcnt_n_0_][0] ),
        .O(\r[rfcnt][2]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r[rfcnt][2]_i_2 
       (.I0(\r[rfcnt][2]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I2(\r[rfcnt][2]_i_6_n_0 ),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .O(\m100.u0/ethc0/v[rfcnt] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8BBBFFFFB8880000)) 
    \r[rfcnt][2]_i_3 
       (.I0(\r[rfcnt][2]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I2(\r[rfcnt][2]_i_8_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rfcnt_n_0_][0] ),
        .O(\m100.u0/ethc0/v[rfcnt] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r[rfcnt][2]_i_4 
       (.I0(\r[rfcnt][2]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rfcnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\r[rfcnt][2]_i_10_n_0 ),
        .O(\m100.u0/ethc0/v[rfcnt] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30B830FF00030000)) 
    \r[rfcnt][2]_i_5 
       (.I0(\r[rfrpnt][0]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\r[rfrpnt][1]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]154_out ),
        .I4(\r[rfcnt][2]_i_11_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .O(\r[rfcnt][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF10000000)) 
    \r[rfcnt][2]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rfcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[rfcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/rmsti[ready] ),
        .I3(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I5(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .O(\r[rfcnt][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r[rfcnt][2]_i_7 
       (.I0(\m100.u0/ethc0/v[ctrlpkt]69_out ),
        .I1(\r[rxcnt][10]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\r[rfrpnt][1]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[rfcnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/v[rmsto][req]57_out ),
        .O(\r[rfcnt][2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r[rfcnt][2]_i_8 
       (.I0(\m100.u0/ethc0/ahb0/r_reg ),
        .I1(\ahbmi[hready] ),
        .I2(\ahbmi[hresp] [1]),
        .I3(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I4(\ahbmi[hresp] [0]),
        .I5(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .O(\r[rfcnt][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30FF30740000008B)) 
    \r[rfcnt][2]_i_9 
       (.I0(\r[rfrpnt][1]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\r[rfrpnt][1]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/v[writeok]154_out ),
        .I4(\m100.u0/ethc0/r_reg[rfcnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[rfcnt_n_0_][1] ),
        .O(\r[rfcnt][2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    \r[rfrpnt][0]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I1(\m100.u0/ethc0/rmsti[ready] ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rfrpnt_n_0_][0] ),
        .O(\r[rfrpnt][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8FFFFBB880000)) 
    \r[rfrpnt][0]_i_3 
       (.I0(\r[rfrpnt][0]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\r[rfrpnt][1]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/v[rmsto][req]57_out ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rfrpnt_n_0_][0] ),
        .O(\r[rfrpnt][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h090909090909090A)) 
    \r[rfrpnt][0]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[rfrpnt_n_0_][0] ),
        .I1(\r[rfrpnt][0]_i_6_n_0 ),
        .I2(\m100.u0/ethc0/v[writeok]154_out ),
        .I3(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[rfcnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[rfcnt_n_0_][0] ),
        .O(\r[rfrpnt][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000004440404040)) 
    \r[rfrpnt][0]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[edclactive_n_0_] ),
        .I1(\r[status][toosmall]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxburstav]__0 ),
        .I3(\m100.u0/ethc0/v[status][toosmall]2 ),
        .I4(\m100.u0/ethc0/p_0_in153_in ),
        .I5(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .O(\m100.u0/ethc0/v[rmsto][req]57_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[rfrpnt][0]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I1(\r_reg[rxcnt][10]_i_8_n_2 ),
        .O(\r[rfrpnt][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r[rfrpnt][1]_i_1 
       (.I0(\r[rfrpnt][1]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rfrpnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\r[rfrpnt][1]_i_3_n_0 ),
        .O(\m100.u0/rxraddress [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3030000074FF8B00)) 
    \r[rfrpnt][1]_i_2 
       (.I0(\r[rfrpnt][1]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\r[rfrpnt][1]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rfrpnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[rfrpnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/v[writeok]154_out ),
        .O(\r[rfrpnt][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7FFFFFFF80000000)) 
    \r[rfrpnt][1]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rfrpnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/rmsti[ready] ),
        .I2(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rfrpnt_n_0_][1] ),
        .O(\r[rfrpnt][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBBBB0)) 
    \r[rfrpnt][1]_i_4 
       (.I0(\r_reg[rxcnt][10]_i_8_n_2 ),
        .I1(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I2(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[rfcnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[rfcnt_n_0_][0] ),
        .O(\r[rfrpnt][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDDDCDCDCFFFCFFF)) 
    \r[rfrpnt][1]_i_5 
       (.I0(\m100.u0/ethc0/p_0_in153_in ),
        .I1(\m100.u0/ethc0/r_reg[edclactive_n_0_] ),
        .I2(\r[status][toosmall]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxburstav]__0 ),
        .I4(\m100.u0/ethc0/v[status][toosmall]2 ),
        .I5(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .O(\r[rfrpnt][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h54450330)) 
    \r[rfwpnt][0]_i_1 
       (.I0(\m100.u0/ethc0/v[rxlength] ),
        .I1(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I3(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I4(\m100.u0/rxwaddress [0]),
        .O(\r[rfwpnt][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h33353533000A0A00)) 
    \r[rfwpnt][1]_i_1 
       (.I0(\m100.u0/rxwaddress [0]),
        .I1(\m100.u0/ethc0/v[rxlength] ),
        .I2(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I4(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I5(\m100.u0/rxwaddress [1]),
        .O(\r[rfwpnt][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000A00000000000)) 
    \r[rfwpnt][1]_i_2 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/p_0_in153_in ),
        .I3(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I4(\m100.u0/ethc0/r_reg[edclactive_n_0_] ),
        .I5(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .O(\m100.u0/ethc0/v[rxlength] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][13]_i_2 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [16]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [16]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][13]_i_3 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [15]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [15]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][13]_i_4 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [14]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [14]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][13]_i_5 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [13]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [13]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][13]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][13]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][13]_i_10_n_4 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][16] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][16] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][13]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][13]_i_10_n_5 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][15] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][15] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][13]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][13]_i_10_n_6 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][14] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][14] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][13]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][13]_i_10_n_7 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][13] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][13] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][17]_i_2 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [20]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [20]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][17]_i_3 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [19]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [19]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][17]_i_4 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [18]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [18]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][17]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][17]_i_5 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [17]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [17]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][17]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][17]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][17]_i_10_n_4 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][20] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][20] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][17]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][17]_i_10_n_5 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][19] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][19] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][17]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][17]_i_10_n_6 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][18] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][18] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][17]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][17]_i_10_n_7 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][17] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][17] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAFFAAAAFFFEBBFE)) 
    \r[rmsto][addr][1]_i_1 
       (.I0(\m100.u0/ethc0/rmsti[retry] ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/p_6_in [1]),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/rmsti[grant] ),
        .I5(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .O(\r[rmsto][addr][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \r[rmsto][addr][1]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[rmsto][addr] [2]),
        .O(\r[rmsto][addr][1]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][1]_i_3 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [4]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [4]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][1]_i_4 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [3]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [3]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][1]_i_5 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [2]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [2]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8B8B888888888)) 
    \r[rmsto][addr][1]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rmsto][addr] [1]),
        .I1(\m100.u0/ethc0/rmsti[retry] ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\r_reg[rmsto][addr][1]_i_10_n_7 ),
        .O(\r[rmsto][addr][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][1]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][1]_i_10_n_4 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][4] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdsel_n_0_][4] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][1]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][1]_i_10_n_5 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][3] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdsel_n_0_][3] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFE30AA00)) 
    \r[rmsto][addr][1]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/r_reg[rxaddr_n_0_][2] ),
        .I3(\r_reg[rmsto][addr][1]_i_10_n_6 ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][21]_i_2 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [24]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [24]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][21]_i_3 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [23]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [23]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][21]_i_4 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [22]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [22]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][21]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][21]_i_5 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [21]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [21]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][21]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][21]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][21]_i_10_n_4 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][24] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][24] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][21]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][21]_i_10_n_5 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][23] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][23] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][21]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][21]_i_10_n_6 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][22] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][22] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][21]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][21]_i_10_n_7 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][21] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][21] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][25]_i_2 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [28]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [28]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][25]_i_3 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [27]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [27]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][25]_i_4 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [26]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [26]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][25]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][25]_i_5 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [25]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [25]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][25]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][25]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][25]_i_10_n_4 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][28] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][28] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][25]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][25]_i_10_n_5 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][27] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][27] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][25]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][25]_i_10_n_6 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][26] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][26] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][25]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][25]_i_10_n_7 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][25] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][25] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC5CCCCCCCCCCCCCC)) 
    \r[rmsto][addr][29]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rmsto][addr] [31]),
        .I1(\m100.u0/ethc0/v[rmsto][addr] [31]),
        .I2(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I3(\ahbmi[hresp] [1]),
        .I4(\m100.u0/ethc0/ahb0/r_reg ),
        .I5(\ahbmi[hready] ),
        .O(\r[rmsto][addr][29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][29]_i_3 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [30]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [30]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][29]_i_4 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [29]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [29]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][29]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][29]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][29]_i_8_n_5 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][31] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][31] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][29]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][29]_i_8_n_6 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][30] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][30] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][29]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][29]_i_8_n_7 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][29] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][29] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][5]_i_2 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [8]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [8]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][5]_i_3 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [7]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [7]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][5]_i_4 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [6]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [6]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][5]_i_5 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [5]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [5]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][5]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][5]_i_10_n_4 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][8] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdsel_n_0_][8] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][5]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][5]_i_10_n_5 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][7] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdsel_n_0_][7] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][5]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][5]_i_10_n_6 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][6] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdsel_n_0_][6] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][5]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][5]_i_10_n_7 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][5] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdsel_n_0_][5] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][9]_i_2 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [12]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [12]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][9]_i_3 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [11]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [11]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][9]_i_4 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [10]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [10]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA3AAAAAAA)) 
    \r[rmsto][addr][9]_i_5 
       (.I0(\m100.u0/ethc0/v[rmsto][addr] [9]),
        .I1(\m100.u0/ethc0/r_reg[rmsto][addr] [9]),
        .I2(\ahbmi[hready] ),
        .I3(\m100.u0/ethc0/ahb0/r_reg ),
        .I4(\ahbmi[hresp] [1]),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[rmsto][addr][9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][9]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][9]_i_10_n_4 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][12] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][12] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][9]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][9]_i_10_n_5 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][11] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][11] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][9]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][9]_i_10_n_6 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][10] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdesc_n_0_][10] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCDC8DDDDCDC88888)) 
    \r[rmsto][addr][9]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\r_reg[rmsto][addr][9]_i_10_n_7 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxaddr_n_0_][9] ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdsel_n_0_][9] ),
        .O(\m100.u0/ethc0/v[rmsto][addr] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[rmsto][data][0]_i_1 
       (.I0(\m100.u0/rxrdata [0]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][0] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[rmsto][data][10]_i_1 
       (.I0(\m100.u0/rxrdata [10]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][10] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r[rmsto][data][14]_i_1 
       (.I0(\m100.u0/rxrdata [14]),
        .I1(\m100.u0/ethc0/r_reg[rxstatus_n_0_][0] ),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r[rmsto][data][15]_i_1 
       (.I0(\m100.u0/rxrdata [15]),
        .I1(\m100.u0/ethc0/r_reg[rxstatus_n_0_][1] ),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r[rmsto][data][16]_i_1 
       (.I0(\m100.u0/rxrdata [16]),
        .I1(\m100.u0/ethc0/r_reg[rxstatus_n_0_][2] ),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[rmsto][data][17]_i_1 
       (.I0(\m100.u0/rxrdata [17]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/p_0_in153_in ),
        .O(\m100.u0/ethc0/v[rmsto][data] [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h45A0)) 
    \r[rmsto][data][18]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/rmsti[ready] ),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .O(\r[rmsto][data][18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r[rmsto][data][18]_i_2 
       (.I0(\m100.u0/rxrdata [18]),
        .I1(\m100.u0/ethc0/p_1_in4_in ),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[rmsto][data][1]_i_1 
       (.I0(\m100.u0/rxrdata [1]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][1] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[rmsto][data][2]_i_1 
       (.I0(\m100.u0/rxrdata [2]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \r[rmsto][data][31]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .O(\r[rmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[rmsto][data][3]_i_1 
       (.I0(\m100.u0/rxrdata [3]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[rmsto][data][4]_i_1 
       (.I0(\m100.u0/rxrdata [4]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][4] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[rmsto][data][5]_i_1 
       (.I0(\m100.u0/rxrdata [5]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][5] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[rmsto][data][6]_i_1 
       (.I0(\m100.u0/rxrdata [6]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][6] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[rmsto][data][7]_i_1 
       (.I0(\m100.u0/rxrdata [7]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][7] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[rmsto][data][8]_i_1 
       (.I0(\m100.u0/rxrdata [8]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][8] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[rmsto][data][9]_i_1 
       (.I0(\m100.u0/rxrdata [9]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][9] ),
        .O(\m100.u0/ethc0/v[rmsto][data] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFABFBFFFFA808)) 
    \r[rmsto][req]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][req] ),
        .I1(\r[rmsto][req]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I3(\r[rmsto][req]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/rmsti[retry] ),
        .I5(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .O(\r[rmsto][req]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h2222222B)) 
    \r[rmsto][req]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][10] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][9] ),
        .I3(\r[rmsto][req]_i_28_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .O(\r[rmsto][req]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h02AAABFC0002AAA8)) 
    \r[rmsto][req]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .I2(\r[rmsto][req]_i_29_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][8] ),
        .I4(\m100.u0/ethc0/r_reg[rxlength_n_0_][9] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .O(\r[rmsto][req]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAA85556)) 
    \r[rmsto][req]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][10] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][9] ),
        .I2(\r[rmsto][req]_i_28_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ),
        .O(\r[rmsto][req]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9090900609090990)) 
    \r[rmsto][req]_i_14 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][9] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][8] ),
        .I3(\r[rmsto][req]_i_29_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .O(\r[rmsto][req]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5701)) 
    \r[rmsto][req]_i_16 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][10] ),
        .I1(\r[rmsto][req]_i_28_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][9] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ),
        .O(\r[rmsto][req]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h2ABC02A8)) 
    \r[rmsto][req]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][8] ),
        .I2(\r[rmsto][req]_i_29_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][9] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .O(\r[rmsto][req]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA856)) 
    \r[rmsto][req]_i_18 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][10] ),
        .I1(\r[rmsto][req]_i_28_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][9] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ),
        .O(\r[rmsto][req]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h90060990)) 
    \r[rmsto][req]_i_19 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][9] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][8] ),
        .I3(\r[rmsto][req]_i_29_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .O(\r[rmsto][req]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00550055FC55FC00)) 
    \r[rmsto][req]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I2(\m100.u0/ethc0/r_reg[rxburstav]__0 ),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/p_6_in [1]),
        .I5(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .O(\m100.u0/ethc0/v[rmsto][req] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h02AAABFC0002AAA8)) 
    \r[rmsto][req]_i_20 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .I2(\r[rmsto][req]_i_38_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][6] ),
        .I4(\m100.u0/ethc0/r_reg[rxlength_n_0_][7] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .O(\r[rmsto][req]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0A2AAFBC0002AAA8)) 
    \r[rmsto][req]_i_21 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[rxlength_n_0_][5] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .O(\r[rmsto][req]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB288)) 
    \r[rmsto][req]_i_22 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .O(\r[rmsto][req]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    \r[rmsto][req]_i_23 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][0] ),
        .O(\r[rmsto][req]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9090900609090990)) 
    \r[rmsto][req]_i_24 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][6] ),
        .I3(\r[rmsto][req]_i_38_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .O(\r[rmsto][req]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9090900609090990)) 
    \r[rmsto][req]_i_25 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .O(\r[rmsto][req]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4218)) 
    \r[rmsto][req]_i_26 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .O(\r[rmsto][req]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[rmsto][req]_i_27 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .O(\r[rmsto][req]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r[rmsto][req]_i_28 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][8] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][6] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][4] ),
        .I4(\m100.u0/ethc0/r_reg[rxlength_n_0_][5] ),
        .I5(\m100.u0/ethc0/r_reg[rxlength_n_0_][7] ),
        .O(\r[rmsto][req]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \r[rmsto][req]_i_29 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[rxlength_n_0_][6] ),
        .O(\r[rmsto][req]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8A0A8A8FFFFFFFF)) 
    \r[rmsto][req]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/rmsti[grant] ),
        .I2(\m100.u0/ethc0/rmsti ),
        .I3(\r[rmsto][req]_i_6_n_0 ),
        .I4(\r[rmsto][req]_i_7_n_0 ),
        .I5(\m100.u0/ethc0/v[rmsto][write] ),
        .O(\r[rmsto][req]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h2ABC02A8)) 
    \r[rmsto][req]_i_30 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][6] ),
        .I2(\r[rmsto][req]_i_38_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][7] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .O(\r[rmsto][req]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h2ABC02A8)) 
    \r[rmsto][req]_i_31 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][5] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .O(\r[rmsto][req]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h88E8)) 
    \r[rmsto][req]_i_32 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .O(\r[rmsto][req]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    \r[rmsto][req]_i_33 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][0] ),
        .O(\r[rmsto][req]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h90060990)) 
    \r[rmsto][req]_i_34 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][6] ),
        .I3(\r[rmsto][req]_i_38_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .O(\r[rmsto][req]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h90060990)) 
    \r[rmsto][req]_i_35 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][4] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .O(\r[rmsto][req]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6006)) 
    \r[rmsto][req]_i_36 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .O(\r[rmsto][req]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[rmsto][req]_i_37 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .O(\r[rmsto][req]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r[rmsto][req]_i_38 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .O(\r[rmsto][req]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3B3B3B083B383B08)) 
    \r[rmsto][req]_i_4 
       (.I0(\m100.u0/ethc0/v[rmsto][req]57_out ),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/rmsti ),
        .I4(\m100.u0/ethc0/rmsti[grant] ),
        .I5(\m100.u0/ethc0/r_reg[rxburstcnt_n_0_][0] ),
        .O(\r[rmsto][req]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4000)) 
    \r[rmsto][req]_i_5 
       (.I0(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I1(\ahbmi[hresp] [1]),
        .I2(\m100.u0/ethc0/ahb0/r_reg ),
        .I3(\ahbmi[hready] ),
        .O(\m100.u0/ethc0/rmsti[retry] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[rmsto][req]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rxburstcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[rxburstcnt_n_0_][1] ),
        .O(\r[rmsto][req]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h57F7)) 
    \r[rmsto][req]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I1(\m100.u0/ethc0/v[rmsto][req]2136_in ),
        .I2(\m100.u0/ethc0/rmsti[ready] ),
        .I3(\m100.u0/ethc0/v[rmsto][req]2137_in ),
        .O(\r[rmsto][req]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[rpnt][0]_i_1 
       (.I0(\m100.u0/ethc0/v[rpnt] ),
        .I1(\m100.u0/ewaddressm [7]),
        .O(\r[rpnt][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT3 #(
    .INIT(8'h78)) 
    \r[rpnt][1]_i_1 
       (.I0(\m100.u0/ewaddressm [7]),
        .I1(\m100.u0/ethc0/v[rpnt] ),
        .I2(\m100.u0/ewaddressm [8]),
        .O(\r[rpnt][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0020002C00000000)) 
    \r[rpnt][1]_i_2 
       (.I0(\r[rpnt][1]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I4(\r[erxidle]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .O(\m100.u0/ethc0/v[rpnt] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \r[rpnt][1]_i_3 
       (.I0(\r[rxstatus][4]_i_1_n_0 ),
        .I1(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I2(\m100.u0/ethc0/rxo[status] [0]),
        .I3(\m100.u0/ethc0/rxo[gotframe] ),
        .I4(\FSM_sequential_r[edclrstate][2]_i_14_n_0 ),
        .I5(\r[rxstatus][1]_i_1_n_0 ),
        .O(\r[rpnt][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[rstaneg]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[duplexstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[duplexstate_n_0_][0] ),
        .O(\r[rstaneg]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \r[rxaddr][31]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/rmsti[ready] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .O(\m100.u0/ethc0/v[rxaddr] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBFBFBF00)) 
    \r[rxburstav]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rfcnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .O(\m100.u0/ethc0/v[rxburstav] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000CD6EFFFF1080)) 
    \r[rxburstcnt][0]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/rmsti[grant] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\m100.u0/ethc0/rmsti[retry] ),
        .I5(\m100.u0/ethc0/r_reg[rxburstcnt_n_0_][0] ),
        .O(\r[rxburstcnt][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0008000008080000)) 
    \r[rxburstcnt][0]_i_2 
       (.I0(\m100.u0/ethc0/ahb0/r_reg[bg]__0 ),
        .I1(\ahbmi[hready] ),
        .I2(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .O(\m100.u0/ethc0/rmsti[grant] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA14FFFF14AA0000)) 
    \r[rxburstcnt][1]_i_1 
       (.I0(\m100.u0/ethc0/rmsti[retry] ),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[rxburstcnt_n_0_][0] ),
        .I4(\r[rxburstcnt][1]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[rxburstcnt_n_0_][1] ),
        .O(\r[rxburstcnt][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF3291)) 
    \r[rxburstcnt][1]_i_2 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/rmsti[grant] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\m100.u0/ethc0/rmsti[retry] ),
        .O(\r[rxburstcnt][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00828200)) 
    \r[rxbytecount][0]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[rxdone] ),
        .I4(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\r[rxbytecount][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00828200)) 
    \r[rxbytecount][10]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [10]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[rxdone] ),
        .I4(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\r[rxbytecount][10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00828200)) 
    \r[rxbytecount][1]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[rxdone] ),
        .I4(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\r[rxbytecount][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00828200)) 
    \r[rxbytecount][2]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[rxdone] ),
        .I4(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\r[rxbytecount][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00828200)) 
    \r[rxbytecount][3]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[rxdone] ),
        .I4(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\r[rxbytecount][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00828200)) 
    \r[rxbytecount][4]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [4]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[rxdone] ),
        .I4(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\r[rxbytecount][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h09900000)) 
    \r[rxbytecount][5]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I2(\m100.u0/ethc0/r_reg[rxdone] ),
        .I3(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .I4(\m100.u0/ethc0/rxo[byte_count] [5]),
        .O(\r[rxbytecount][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00828200)) 
    \r[rxbytecount][6]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [6]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[rxdone] ),
        .I4(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\r[rxbytecount][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00828200)) 
    \r[rxbytecount][7]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [7]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[rxdone] ),
        .I4(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\r[rxbytecount][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00828200)) 
    \r[rxbytecount][8]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [8]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[rxdone] ),
        .I4(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\r[rxbytecount][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00828200)) 
    \r[rxbytecount][9]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [9]),
        .I1(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[rxdone] ),
        .I4(\m100.u0/ethc0/r_reg[rxdoneack]__0 ),
        .O(\r[rxbytecount][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8B88)) 
    \r[rxcnt][0]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .O(\m100.u0/ethc0/v[rxcnt] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB800003333F3F3)) 
    \r[rxcnt][10]_i_1 
       (.I0(\r[rxcnt][10]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I2(\m100.u0/ethc0/rmsti[ready] ),
        .I3(\m100.u0/ethc0/rmsti ),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .O(\r[rxcnt][10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[rxcnt][10]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[rxbytecount]__0 [10]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ),
        .O(\r[rxcnt][10]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h44D4)) 
    \r[rxcnt][10]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .I1(\m100.u0/ethc0/r_reg[rxbytecount]__0 [9]),
        .I2(\m100.u0/ethc0/r_reg[rxbytecount]__0 [8]),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .O(\r[rxcnt][10]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r[rxcnt][10]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ),
        .I1(\m100.u0/ethc0/r_reg[rxbytecount]__0 [10]),
        .O(\r[rxcnt][10]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[rxcnt][10]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[rxbytecount]__0 [9]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .I2(\m100.u0/ethc0/r_reg[rxbytecount]__0 [8]),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .O(\r[rxcnt][10]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h44D4)) 
    \r[rxcnt][10]_i_14 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[rxbytecount]__0 [7]),
        .I2(\m100.u0/ethc0/r_reg[rxbytecount]__0 [6]),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .O(\r[rxcnt][10]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h44D4)) 
    \r[rxcnt][10]_i_15 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[rxbytecount]__0 [5]),
        .I2(\m100.u0/ethc0/r_reg[rxbytecount]__0 [4]),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .O(\r[rxcnt][10]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h44D4)) 
    \r[rxcnt][10]_i_16 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[rxbytecount]__0 [3]),
        .I2(\m100.u0/ethc0/r_reg[rxbytecount]__0 [2]),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .O(\r[rxcnt][10]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    \r[rxcnt][10]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[rxbytecount]__0 [1]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[rxbytecount]__0 [0]),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .O(\r[rxcnt][10]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[rxcnt][10]_i_18 
       (.I0(\m100.u0/ethc0/r_reg[rxbytecount]__0 [7]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .I2(\m100.u0/ethc0/r_reg[rxbytecount]__0 [6]),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .O(\r[rxcnt][10]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[rxcnt][10]_i_19 
       (.I0(\m100.u0/ethc0/r_reg[rxbytecount]__0 [5]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[rxbytecount]__0 [4]),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .O(\r[rxcnt][10]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h283C282828EC2828)) 
    \r[rxcnt][10]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ),
        .I2(\r[rxcnt][10]_i_6_n_0 ),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\r[rxcnt][10]_i_7_n_0 ),
        .O(\m100.u0/ethc0/v[rxcnt] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[rxcnt][10]_i_20 
       (.I0(\m100.u0/ethc0/r_reg[rxbytecount]__0 [3]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[rxbytecount]__0 [2]),
        .O(\r[rxcnt][10]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[rxcnt][10]_i_21 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[rxbytecount]__0 [1]),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[rxbytecount]__0 [0]),
        .O(\r[rxcnt][10]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5D5D5D5D5D5D5D00)) 
    \r[rxcnt][10]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I1(\r_reg[rxcnt][10]_i_8_n_2 ),
        .I2(\m100.u0/ethc0/p_0_in153_in ),
        .I3(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[rfcnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[rfcnt_n_0_][0] ),
        .O(\r[rxcnt][10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h01000000)) 
    \r[rxcnt][10]_i_4 
       (.I0(\ahbmi[hresp] [0]),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\ahbmi[hresp] [1]),
        .I3(\ahbmi[hready] ),
        .I4(\m100.u0/ethc0/ahb0/r_reg ),
        .O(\m100.u0/ethc0/rmsti[ready] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h04000000)) 
    \r[rxcnt][10]_i_5 
       (.I0(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I1(\ahbmi[hresp] [0]),
        .I2(\ahbmi[hresp] [1]),
        .I3(\ahbmi[hready] ),
        .I4(\m100.u0/ethc0/ahb0/r_reg ),
        .O(\m100.u0/ethc0/rmsti ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \r[rxcnt][10]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .I1(\r[rxcnt][8]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .O(\r[rxcnt][10]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[rxcnt][10]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .O(\r[rxcnt][10]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8B888C88)) 
    \r[rxcnt][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .O(\m100.u0/ethc0/v[rxcnt] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5575757510202020)) 
    \r[rxcnt][2]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .O(\m100.u0/ethc0/v[rxcnt] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h66666E6606000A00)) 
    \r[rxcnt][3]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\r[rxcnt][10]_i_7_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .O(\m100.u0/ethc0/v[rxcnt] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h283C282828EC2828)) 
    \r[rxcnt][4]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .I2(\r[rxcnt][4]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\r[rxcnt][10]_i_7_n_0 ),
        .O(\m100.u0/ethc0/v[rxcnt] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[rxcnt][4]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .O(\r[rxcnt][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h28FF282828282828)) 
    \r[rxcnt][5]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I2(\r[rxcnt][5]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\r[rxcnt][5]_i_3_n_0 ),
        .O(\m100.u0/ethc0/v[rxcnt] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \r[rxcnt][5]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .O(\r[rxcnt][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6AAAAAAAAAAAAAAA)) 
    \r[rxcnt][5]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .O(\r[rxcnt][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h283B282828EC2828)) 
    \r[rxcnt][6]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .I2(\r[rxcnt][6]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\r[rxcnt][6]_i_3_n_0 ),
        .O(\m100.u0/ethc0/v[rxcnt] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \r[rxcnt][6]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .O(\r[rxcnt][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \r[rxcnt][6]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .O(\r[rxcnt][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h283B282828EC2828)) 
    \r[rxcnt][7]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .I2(\r[rxcnt][7]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\r[rxcnt][7]_i_3_n_0 ),
        .O(\m100.u0/ethc0/v[rxcnt] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \r[rxcnt][7]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .O(\r[rxcnt][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \r[rxcnt][7]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I3(\r[rxcnt][10]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .O(\r[rxcnt][7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h28FF282828282828)) 
    \r[rxcnt][8]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .I2(\r[rxcnt][8]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\r[rxcnt][8]_i_3_n_0 ),
        .O(\m100.u0/ethc0/v[rxcnt] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \r[rxcnt][8]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .O(\r[rxcnt][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6AAA)) 
    \r[rxcnt][8]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .I2(\r[rxcnt][6]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .O(\r[rxcnt][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h28FF282828282828)) 
    \r[rxcnt][9]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .I2(\r[rxcnt][9]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\r[rxcnt][9]_i_3_n_0 ),
        .O(\m100.u0/ethc0/v[rxcnt] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \r[rxcnt][9]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I2(\r[rxcnt][4]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .O(\r[rxcnt][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \r[rxcnt][9]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .I3(\r[rxcnt][6]_i_3_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .O(\r[rxcnt][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \r[rxdesc][31]_i_1 
       (.I0(\apbo[prdata][14]_INST_0_i_5_n_0 ),
        .I1(\apbi[pwrite] ),
        .I2(apbi[15]),
        .I3(\apbi[penable] ),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [2]),
        .O(\r[rxdesc][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFF00)) 
    \r[rxdoneold]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I4(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .O(\r[rxdoneold]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF40000000)) 
    \r[rxdsel][3]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\r[rxdsel][3]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/rmsti[ready] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\apbi[pwdata] [3]),
        .O(\m100.u0/ethc0/v[rxdsel] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[rxdsel][3]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxwrap_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][3] ),
        .O(\r[rxdsel][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF40000000)) 
    \r[rxdsel][4]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\r[rxdsel][4]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/rmsti[ready] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\apbi[pwdata] [4]),
        .O(\m100.u0/ethc0/v[rxdsel] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \r[rxdsel][4]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxdsel_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxwrap_n_0_] ),
        .O(\r[rxdsel][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF40000000)) 
    \r[rxdsel][5]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\r[rxdsel][5]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/rmsti[ready] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\apbi[pwdata] [5]),
        .O(\m100.u0/ethc0/v[rxdsel] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1540)) 
    \r[rxdsel][5]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxwrap_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxdsel_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[rxdsel_n_0_][5] ),
        .O(\r[rxdsel][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF40000000)) 
    \r[rxdsel][6]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\r[rxdsel][6]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/rmsti[ready] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\apbi[pwdata] [6]),
        .O(\m100.u0/ethc0/v[rxdsel] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h15554000)) 
    \r[rxdsel][6]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxwrap_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[rxdsel_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[rxdsel_n_0_][5] ),
        .I4(\m100.u0/ethc0/r_reg[rxdsel_n_0_][6] ),
        .O(\r[rxdsel][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFF40000000)) 
    \r[rxdsel][7]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\r[rxdsel][7]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/rmsti[ready] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\apbi[pwdata] [7]),
        .O(\m100.u0/ethc0/v[rxdsel] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1555555540000000)) 
    \r[rxdsel][7]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxwrap_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[rxdsel_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[rxdsel_n_0_][4] ),
        .I4(\m100.u0/ethc0/r_reg[rxdsel_n_0_][6] ),
        .I5(\m100.u0/ethc0/r_reg[rxdsel_n_0_][7] ),
        .O(\r[rxdsel][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEF40)) 
    \r[rxdsel][8]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\r[rxdsel][8]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I3(\apbi[pwdata] [8]),
        .O(\m100.u0/ethc0/v[rxdsel] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h06FFFFFF06000000)) 
    \r[rxdsel][8]_i_2 
       (.I0(\r[rxdsel][9]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][8] ),
        .I2(\m100.u0/ethc0/r_reg[rxwrap_n_0_] ),
        .I3(\m100.u0/ethc0/rmsti[ready] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I5(\apbi[pwdata] [8]),
        .O(\r[rxdsel][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF4000)) 
    \r[rxdsel][9]_i_1 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\m100.u0/ethc0/rmsti[ready] ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\r[rxdesc][31]_i_1_n_0 ),
        .O(\r[rxdsel][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF4000)) 
    \r[rxdsel][9]_i_2 
       (.I0(\m100.u0/ethc0/v[rmsto][write] ),
        .I1(\r[rxdsel][9]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I4(\apbi[pwdata] [9]),
        .O(\m100.u0/ethc0/v[rxdsel] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1540FFFF15400000)) 
    \r[rxdsel][9]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxwrap_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][8] ),
        .I2(\r[rxdsel][9]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[rxdsel_n_0_][9] ),
        .I4(\m100.u0/ethc0/rmsti[ready] ),
        .I5(\apbi[pwdata] [9]),
        .O(\r[rxdsel][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \r[rxdsel][9]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[rxdsel_n_0_][6] ),
        .I1(\m100.u0/ethc0/r_reg[rxdsel_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[rxdsel_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[rxdsel_n_0_][5] ),
        .I4(\m100.u0/ethc0/r_reg[rxdsel_n_0_][7] ),
        .O(\r[rxdsel][9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \r[rxirq]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/rmsti[ready] ),
        .I5(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .O(\m100.u0/ethc0/v[rxwrap] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \r[rxlength][0]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I1(\r[rxlength][10]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/rxo[lentype] [0]),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[rxlength][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFA0200000)) 
    \r[rxlength][10]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/r_reg[edclactive_n_0_] ),
        .I2(\m100.u0/ethc0/v[writeok]154_out ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/v[rmsto][write] ),
        .I5(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\m100.u0/ethc0/v[rxbytecount] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \r[rxlength][10]_i_10 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [8]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [10]),
        .O(\r[rxlength][10]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \r[rxlength][10]_i_2 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [10]),
        .I1(\r[rxlength][10]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/rxo[lentype] [10]),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[rxlength][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[rxlength][10]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I1(\m100.u0/ethc0/p_0_in153_in ),
        .O(\m100.u0/ethc0/v[writeok]154_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000055D1)) 
    \r[rxlength][10]_i_4 
       (.I0(\m100.u0/ethc0/v[rxstatus]2130_in ),
        .I1(\r[rxlength][10]_i_5_n_0 ),
        .I2(\r[rxlength][10]_i_6_n_0 ),
        .I3(\r[rxlength][10]_i_7_n_0 ),
        .I4(\r[rxlength][10]_i_8_n_0 ),
        .O(\r[rxlength][10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \r[rxlength][10]_i_5 
       (.I0(\m100.u0/ethc0/rxo[lentype] [10]),
        .I1(\m100.u0/ethc0/rxo[lentype] [6]),
        .I2(\m100.u0/ethc0/rxo[lentype] [8]),
        .I3(\m100.u0/ethc0/rxo[lentype] [9]),
        .I4(\m100.u0/ethc0/rxo[lentype] [7]),
        .O(\r[rxlength][10]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    \r[rxlength][10]_i_6 
       (.I0(\r[rxlength][10]_i_9_n_0 ),
        .I1(\r[rxlength][10]_i_10_n_0 ),
        .I2(\m100.u0/ethc0/rxo[byte_count] [5]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [2]),
        .O(\r[rxlength][10]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE000000000000000)) 
    \r[rxlength][10]_i_7 
       (.I0(\m100.u0/ethc0/rxo[lentype] [1]),
        .I1(\m100.u0/ethc0/rxo[lentype] [0]),
        .I2(\m100.u0/ethc0/rxo[lentype] [2]),
        .I3(\m100.u0/ethc0/rxo[lentype] [3]),
        .I4(\m100.u0/ethc0/rxo[lentype] [4]),
        .I5(\m100.u0/ethc0/rxo[lentype] [5]),
        .O(\r[rxlength][10]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFFEFEF)) 
    \r[rxlength][10]_i_8 
       (.I0(\r[rxstatus][4]_i_11_n_0 ),
        .I1(\r[rxstatus][4]_i_10_n_0 ),
        .I2(\r[rxstatus][4]_i_5_n_0 ),
        .I3(\r[rxstatus][4]_i_9_n_0 ),
        .I4(\r[rxstatus][4]_i_8_n_0 ),
        .O(\r[rxlength][10]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    \r[rxlength][10]_i_9 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [6]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [7]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [4]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [9]),
        .O(\r[rxlength][10]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \r[rxlength][1]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I1(\r[rxlength][10]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/rxo[lentype] [1]),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[rxlength][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \r[rxlength][2]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I1(\r[rxlength][10]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/rxo[lentype] [2]),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[rxlength][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \r[rxlength][3]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I1(\r[rxlength][10]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/rxo[lentype] [3]),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[rxlength][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \r[rxlength][4]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [4]),
        .I1(\r[rxlength][10]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/rxo[lentype] [4]),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[rxlength][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \r[rxlength][5]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [5]),
        .I1(\r[rxlength][10]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/rxo[lentype] [5]),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[rxlength][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \r[rxlength][6]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [6]),
        .I1(\r[rxlength][10]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/rxo[lentype] [6]),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[rxlength][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \r[rxlength][7]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [7]),
        .I1(\r[rxlength][10]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/rxo[lentype] [7]),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[rxlength][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \r[rxlength][8]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [8]),
        .I1(\r[rxlength][10]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/rxo[lentype] [8]),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[rxlength][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \r[rxlength][9]_i_1 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [9]),
        .I1(\r[rxlength][10]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/rxo[lentype] [9]),
        .I3(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[rxlength][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    \r[rxstart][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I1(\r[rxstart][1]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .O(\r[rxstart][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000008B8B00)) 
    \r[rxstart][1]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxden]__0 ),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/p_6_in [1]),
        .I3(\m100.u0/ethc0/r_reg[rxstart]__0 [0]),
        .I4(\m100.u0/ethc0/r_reg[rxstart]__0 [1]),
        .I5(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .O(\r[rxstart][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBBB8B88888888)) 
    \r[rxstatus][0]_i_1 
       (.I0(\m100.u0/ethc0/rxo[status] [0]),
        .I1(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I5(\m100.u0/ethc0/r_reg[rxstatus_n_0_][0] ),
        .O(\r[rxstatus][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBBB8B88888888)) 
    \r[rxstatus][1]_i_1 
       (.I0(\m100.u0/ethc0/rxo[status] [1]),
        .I1(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I5(\m100.u0/ethc0/r_reg[rxstatus_n_0_][1] ),
        .O(\r[rxstatus][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBBB8B88888888)) 
    \r[rxstatus][2]_i_1 
       (.I0(\m100.u0/ethc0/rxo[status] [2]),
        .I1(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I3(\m100.u0/ethc0/v[rmsto][write] ),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I5(\m100.u0/ethc0/r_reg[rxstatus_n_0_][2] ),
        .O(\r[rxstatus][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8BBBB88888888)) 
    \r[rxstatus][3]_i_1 
       (.I0(\m100.u0/ethc0/rxo[status] [3]),
        .I1(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .I2(\m100.u0/ethc0/v[rmsto][write] ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I5(\m100.u0/ethc0/p_0_in153_in ),
        .O(\r[rxstatus][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBAAAAAABAAABAAA)) 
    \r[rxstatus][4]_i_1 
       (.I0(\m100.u0/ethc0/v[rxstatus] ),
        .I1(\r[rxstatus][4]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/v[rxstatus]2130_in ),
        .I3(\r[rxstatus][4]_i_5_n_0 ),
        .I4(\r[rxstatus][4]_i_6_n_0 ),
        .I5(\r[rxstatus][4]_i_7_n_0 ),
        .O(\r[rxstatus][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF8)) 
    \r[rxstatus][4]_i_10 
       (.I0(\m100.u0/ethc0/rxo[lentype] [10]),
        .I1(\m100.u0/ethc0/rxo[lentype] [9]),
        .I2(\m100.u0/ethc0/rxo[lentype] [12]),
        .I3(\m100.u0/ethc0/rxo[status] [3]),
        .O(\r[rxstatus][4]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r[rxstatus][4]_i_11 
       (.I0(\m100.u0/ethc0/rxo[lentype] [14]),
        .I1(\m100.u0/ethc0/rxo[lentype] [15]),
        .I2(\m100.u0/ethc0/rxo[lentype] [13]),
        .I3(\m100.u0/ethc0/rxo[lentype] [11]),
        .O(\r[rxstatus][4]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[rxstatus][4]_i_12 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [9]),
        .I1(\m100.u0/ethc0/rxo[lentype] [9]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [10]),
        .I3(\m100.u0/ethc0/rxo[lentype] [10]),
        .O(\r[rxstatus][4]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[rxstatus][4]_i_13 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [7]),
        .I1(\m100.u0/ethc0/rxo[lentype] [7]),
        .I2(\m100.u0/ethc0/rxo[lentype] [8]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [8]),
        .I4(\m100.u0/ethc0/rxo[lentype] [6]),
        .I5(\m100.u0/ethc0/rxo[byte_count] [6]),
        .O(\r[rxstatus][4]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[rxstatus][4]_i_14 
       (.I0(\m100.u0/ethc0/rxo[lentype] [5]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [5]),
        .I2(\m100.u0/ethc0/rxo[lentype] [4]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [4]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [3]),
        .I5(\m100.u0/ethc0/rxo[lentype] [3]),
        .O(\r[rxstatus][4]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \r[rxstatus][4]_i_15 
       (.I0(\m100.u0/ethc0/rxo[lentype] [2]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [2]),
        .I2(\m100.u0/ethc0/rxo[lentype] [1]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I5(\m100.u0/ethc0/rxo[lentype] [0]),
        .O(\r[rxstatus][4]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r[rxstatus][4]_i_16 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [7]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [6]),
        .O(\r[rxstatus][4]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFEFFFFFF)) 
    \r[rxstatus][4]_i_17 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [10]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [1]),
        .I2(\m100.u0/ethc0/rxo[byte_count] [0]),
        .I3(\m100.u0/ethc0/rxo[byte_count] [5]),
        .I4(\m100.u0/ethc0/rxo[byte_count] [2]),
        .O(\r[rxstatus][4]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFD00)) 
    \r[rxstatus][4]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rxdstate] [0]),
        .I1(\m100.u0/ethc0/v[rmsto][write] ),
        .I2(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I3(\m100.u0/ethc0/p_1_in4_in ),
        .O(\m100.u0/ethc0/v[rxstatus] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFF2FFFFFFFFF)) 
    \r[rxstatus][4]_i_3 
       (.I0(\r[rxstatus][4]_i_8_n_0 ),
        .I1(\r[rxstatus][4]_i_9_n_0 ),
        .I2(\r[rxstatus][4]_i_5_n_0 ),
        .I3(\r[rxstatus][4]_i_10_n_0 ),
        .I4(\r[rxstatus][4]_i_11_n_0 ),
        .I5(\m100.u0/ethc0/v[rxstatus]1135_out ),
        .O(\r[rxstatus][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \r[rxstatus][4]_i_5 
       (.I0(\m100.u0/ethc0/rxo[status] [0]),
        .I1(\m100.u0/ethc0/rxo[status] [2]),
        .I2(\m100.u0/ethc0/rxo[status] [1]),
        .O(\r[rxstatus][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFBFFFFFFFF)) 
    \r[rxstatus][4]_i_6 
       (.I0(\m100.u0/ethc0/rxo[byte_count] [8]),
        .I1(\m100.u0/ethc0/rxo[byte_count] [4]),
        .I2(\r[rxstatus][4]_i_16_n_0 ),
        .I3(\r[rxstatus][4]_i_17_n_0 ),
        .I4(\m100.u0/ethc0/rxo[byte_count] [9]),
        .I5(\m100.u0/ethc0/rxo[byte_count] [3]),
        .O(\r[rxstatus][4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \r[rxstatus][4]_i_7 
       (.I0(\m100.u0/ethc0/rxo[lentype] [7]),
        .I1(\m100.u0/ethc0/rxo[lentype] [9]),
        .I2(\m100.u0/ethc0/rxo[lentype] [8]),
        .I3(\m100.u0/ethc0/rxo[lentype] [6]),
        .I4(\m100.u0/ethc0/rxo[lentype] [10]),
        .I5(\r[rxlength][10]_i_7_n_0 ),
        .O(\r[rxstatus][4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEAAAAA)) 
    \r[rxstatus][4]_i_8 
       (.I0(\m100.u0/ethc0/rxo[lentype] [4]),
        .I1(\m100.u0/ethc0/rxo[lentype] [1]),
        .I2(\m100.u0/ethc0/rxo[lentype] [0]),
        .I3(\m100.u0/ethc0/rxo[lentype] [2]),
        .I4(\m100.u0/ethc0/rxo[lentype] [3]),
        .O(\r[rxstatus][4]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \r[rxstatus][4]_i_9 
       (.I0(\m100.u0/ethc0/rxo[lentype] [8]),
        .I1(\m100.u0/ethc0/rxo[lentype] [6]),
        .I2(\m100.u0/ethc0/rxo[lentype] [7]),
        .I3(\m100.u0/ethc0/rxo[lentype] [5]),
        .I4(\m100.u0/ethc0/rxo[lentype] [10]),
        .O(\r[rxstatus][4]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[seq][0]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[nak_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .O(\m100.u0/ethc0/v[seq] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \r[seq][0]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[seq] [0]),
        .O(\r[seq][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F2F2F2)) 
    \r[status][invaddr]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[addrdone]__0 ),
        .I1(\m100.u0/ethc0/r_reg[addrok_n_0_] ),
        .I2(\m100.u0/ethc0/r_reg[ctrlpkt]__0 ),
        .I3(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I4(\m100.u0/ethc0/p_0_in153_in ),
        .I5(\m100.u0/ethc0/r_reg[edclactive_n_0_] ),
        .O(\r[status][invaddr]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \r[status][invaddr]_i_3 
       (.I0(\r[status][txahberr]_i_2_n_0 ),
        .I1(\apbi[pwdata] [7]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [5]),
        .O(\m100.u0/ethc0/v[status][invaddr]45_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    \r[status][rx_err]_i_2 
       (.I0(\m100.u0/ethc0/rmsti[ready] ),
        .I1(\m100.u0/ethc0/p_0_in153_in ),
        .I2(\m100.u0/ethc0/r_reg[rxstatus_n_0_][2] ),
        .I3(\m100.u0/ethc0/p_1_in4_in ),
        .I4(\m100.u0/ethc0/r_reg[rxstatus_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[rxstatus_n_0_][1] ),
        .O(\m100.u0/ethc0/v[status][rx_err]15_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \r[status][rx_err]_i_3 
       (.I0(\r[status][txahberr]_i_2_n_0 ),
        .I1(\apbi[pwdata] [0]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [5]),
        .O(\m100.u0/ethc0/v[status][rx_err]18_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \r[status][rx_int]_i_2 
       (.I0(\m100.u0/ethc0/p_0_in153_in ),
        .I1(\m100.u0/ethc0/r_reg[rxstatus_n_0_][2] ),
        .I2(\m100.u0/ethc0/p_1_in4_in ),
        .I3(\m100.u0/ethc0/r_reg[rxstatus_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[rxstatus_n_0_][1] ),
        .I5(\m100.u0/ethc0/rmsti[ready] ),
        .O(\r[status][rx_int]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \r[status][rx_int]_i_3 
       (.I0(\r[status][txahberr]_i_2_n_0 ),
        .I1(\apbi[pwdata] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [5]),
        .O(\m100.u0/ethc0/v[status][rx_int]26_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \r[status][rxahberr]_i_2 
       (.I0(\r[status][txahberr]_i_2_n_0 ),
        .I1(\apbi[pwdata] [4]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [5]),
        .O(\m100.u0/ethc0/v[status][rxahberr]32_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[status][toosmall]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][9] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][8] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .O(\r[status][toosmall]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    \r[status][toosmall]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][7] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][6] ),
        .O(\r[status][toosmall]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    \r[status][toosmall]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][4] ),
        .O(\r[status][toosmall]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    \r[status][toosmall]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .O(\r[status][toosmall]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    \r[status][toosmall]_i_14 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][0] ),
        .O(\r[status][toosmall]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[status][toosmall]_i_15 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][7] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][6] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][6] ),
        .O(\r[status][toosmall]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[status][toosmall]_i_16 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][4] ),
        .O(\r[status][toosmall]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[status][toosmall]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][2] ),
        .O(\r[status][toosmall]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[status][toosmall]_i_18 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[rxlength_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[rxcnt_n_0_][0] ),
        .O(\r[status][toosmall]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000002000)) 
    \r[status][toosmall]_i_2 
       (.I0(\r[status][toosmall]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[gotframe_n_0_] ),
        .I2(\m100.u0/ethc0/v[status][toosmall]2 ),
        .I3(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I4(\m100.u0/ethc0/r_reg[edclactive_n_0_] ),
        .I5(\m100.u0/ethc0/p_0_in153_in ),
        .O(\m100.u0/ethc0/v[status][toosmall]39_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \r[status][toosmall]_i_3 
       (.I0(\r[status][txahberr]_i_2_n_0 ),
        .I1(\apbi[pwdata] [6]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [5]),
        .O(\m100.u0/ethc0/v[status][toosmall]42_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h45)) 
    \r[status][toosmall]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[ctrlpkt]__0 ),
        .I1(\m100.u0/ethc0/r_reg[addrok_n_0_] ),
        .I2(\m100.u0/ethc0/r_reg[addrdone]__0 ),
        .O(\r[status][toosmall]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[status][toosmall]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][10] ),
        .O(\r[status][toosmall]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    \r[status][toosmall]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[rxcnt_n_0_][9] ),
        .I1(\m100.u0/ethc0/r_reg[rxlength_n_0_][9] ),
        .I2(\m100.u0/ethc0/r_reg[rxcnt_n_0_][8] ),
        .I3(\m100.u0/ethc0/r_reg[rxlength_n_0_][8] ),
        .O(\r[status][toosmall]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r[status][toosmall]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[rxlength_n_0_][10] ),
        .I1(\m100.u0/ethc0/r_reg[rxcnt_n_0_][10] ),
        .O(\r[status][toosmall]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \r[status][tx_int]_i_2 
       (.I0(\apbi[paddr] [5]),
        .I1(\apbi[paddr] [3]),
        .I2(\r[status][txahberr]_i_2_n_0 ),
        .O(\r[status][tx_int]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    \r[status][txahberr]_i_2 
       (.I0(\apbi[paddr] [4]),
        .I1(\apbi[pwrite] ),
        .I2(apbi[15]),
        .I3(\apbi[penable] ),
        .I4(\apbi[paddr] [2]),
        .O(\r[status][txahberr]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \r[tarp]_i_2 
       (.I0(\m100.u0/erdata [26]),
        .I1(\m100.u0/erdata [29]),
        .I2(\m100.u0/erdata [17]),
        .I3(\m100.u0/erdata [19]),
        .I4(\r[tarp]_i_4_n_0 ),
        .O(\r[tarp]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \r[tarp]_i_3 
       (.I0(\m100.u0/erdata [16]),
        .I1(\m100.u0/erdata [30]),
        .I2(\m100.u0/erdata [20]),
        .I3(\m100.u0/erdata [21]),
        .I4(\r[tarp]_i_5_n_0 ),
        .O(\r[tarp]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    \r[tarp]_i_4 
       (.I0(\m100.u0/erdata [28]),
        .I1(\m100.u0/erdata [25]),
        .I2(\m100.u0/erdata [27]),
        .I3(\m100.u0/erdata [23]),
        .O(\r[tarp]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFD)) 
    \r[tarp]_i_5 
       (.I0(\m100.u0/erdata [18]),
        .I1(\m100.u0/erdata [31]),
        .I2(\m100.u0/erdata [24]),
        .I3(\m100.u0/erdata [22]),
        .O(\r[tarp]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h34333434)) 
    \r[tcnt][0]_i_1 
       (.I0(\r[tcnt][6]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I2(\r[tcnt][4]_i_5_n_0 ),
        .I3(\r[tcnt][4]_i_3_n_0 ),
        .I4(\r[tcnt][4]_i_6_n_0 ),
        .O(\m100.u0/eraddress [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCFB8)) 
    \r[tcnt][1]_i_1 
       (.I0(\r[tcnt][6]_i_4_n_0 ),
        .I1(\r[tcnt][6]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .O(\m100.u0/eraddress [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABBAAAAAABBABABA)) 
    \r[tcnt][2]_i_1 
       (.I0(\r[tcnt][2]_i_2_n_0 ),
        .I1(\r[tcnt][4]_i_6_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I3(\r[tcnt][3]_i_2_n_0 ),
        .I4(\r[tcnt][4]_i_5_n_0 ),
        .I5(\r[tcnt][6]_i_4_n_0 ),
        .O(\m100.u0/eraddress [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0007070705050005)) 
    \r[tcnt][2]_i_2 
       (.I0(\r[tcnt][4]_i_3_n_0 ),
        .I1(\r[tcnt][6]_i_4_n_0 ),
        .I2(\r[tcnt][2]_i_3_n_0 ),
        .I3(\r[tcnt][4]_i_8_n_0 ),
        .I4(\r[tcnt][3]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .O(\r[tcnt][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8222A222FFFFFFFF)) 
    \r[tcnt][2]_i_3 
       (.I0(\r[tcnt][2]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .I4(\r[txdstate][2]_i_5_n_0 ),
        .I5(\r[tcnt][4]_i_6_n_0 ),
        .O(\r[tcnt][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4808)) 
    \r[tcnt][2]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[tcnt][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCC8888CFFFB888)) 
    \r[tcnt][3]_i_1 
       (.I0(\r[tcnt][6]_i_4_n_0 ),
        .I1(\r[tcnt][6]_i_2_n_0 ),
        .I2(\r[tcnt][3]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[tcnt_n_0_][3] ),
        .I5(\r[tcnt][3]_i_3_n_0 ),
        .O(\m100.u0/eraddress [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[tcnt][3]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .O(\r[tcnt][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000010400040)) 
    \r[tcnt][3]_i_3 
       (.I0(\r[tcnt][4]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\r[txdstate][2]_i_2_n_0 ),
        .O(\r[tcnt][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF555F5FFF111F111)) 
    \r[tcnt][4]_i_1 
       (.I0(\r[tcnt][4]_i_2_n_0 ),
        .I1(\r[tcnt][4]_i_3_n_0 ),
        .I2(\r[tcnt][4]_i_4_n_0 ),
        .I3(\r[tcnt][4]_i_5_n_0 ),
        .I4(\r[tcnt][4]_i_6_n_0 ),
        .I5(\r[tcnt][4]_i_7_n_0 ),
        .O(\m100.u0/eraddress [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3FFFFCFFBFFFFEF)) 
    \r[tcnt][4]_i_2 
       (.I0(\r[tcnt][4]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\r[tcnt][4]_i_4_n_0 ),
        .O(\r[tcnt][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010000000100010)) 
    \r[tcnt][4]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\r[txdstate][1]_i_6_n_0 ),
        .I5(\r[tedcl]_i_2_n_0 ),
        .O(\r[tcnt][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6AAAAAAA)) 
    \r[tcnt][4]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .O(\r[tcnt][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \r[tcnt][4]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\r[tcnt][4]_i_9_n_0 ),
        .O(\r[tcnt][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6004)) 
    \r[tcnt][4]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[tcnt][4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[tcnt][4]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][4] ),
        .I1(\r[tcnt][6]_i_4_n_0 ),
        .O(\r[tcnt][4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDF7DFFFFDF7DDF7D)) 
    \r[tcnt][4]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\r[txdstate][1]_i_6_n_0 ),
        .I5(\r[tedcl]_i_2_n_0 ),
        .O(\r[tcnt][4]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFBFFFFFF)) 
    \r[tcnt][4]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\ahbmi[hresp] [1]),
        .I3(\ahbmi[hready] ),
        .I4(\m100.u0/ethc0/ahb0/r_reg ),
        .O(\r[tcnt][4]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4370)) 
    \r[tcnt][5]_i_1 
       (.I0(\r[tcnt][6]_i_4_n_0 ),
        .I1(\r[tcnt][6]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][5] ),
        .I3(\r[tcnt][6]_i_3_n_0 ),
        .O(\m100.u0/eraddress [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00009AAA)) 
    \r[tcnt][6]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][6] ),
        .I1(\r[tcnt][6]_i_2_n_0 ),
        .I2(\r[tcnt][6]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][5] ),
        .I4(\r[tcnt][6]_i_4_n_0 ),
        .O(\m100.u0/eraddress [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAEBFFFFEF)) 
    \r[tcnt][6]_i_2 
       (.I0(\r[tcnt][4]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\r[tcnt][4]_i_5_n_0 ),
        .O(\r[tcnt][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \r[tcnt][6]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .O(\r[tcnt][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FE00000000)) 
    \r[tcnt][6]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[abufs_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg ),
        .I3(\m100.u0/ethc0/p_6_in [14]),
        .I4(\r[tfwpnt][6]_i_3_n_0 ),
        .I5(\r[tcnt][6]_i_5_n_0 ),
        .O(\r[tcnt][6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[tcnt][6]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\r[tcnt][6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000FEFF)) 
    \r[tedcl]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I2(\r[txcnt][10]_i_9_n_0 ),
        .I3(\r[txcnt][6]_i_8_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tarp]__0 ),
        .I5(\m100.u0/ethc0/r_reg[tnak]__0 ),
        .O(\r[tedcl]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44454440)) 
    \r[tfcnt][0]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\r_reg[tfcnt][3]_i_2_n_7 ),
        .I2(\r[tfcnt][7]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r_reg[tfcnt][3]_i_3_n_7 ),
        .O(\r[tfcnt][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44454440)) 
    \r[tfcnt][1]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\r_reg[tfcnt][3]_i_2_n_6 ),
        .I2(\r[tfcnt][7]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r_reg[tfcnt][3]_i_3_n_6 ),
        .O(\r[tfcnt][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44454440)) 
    \r[tfcnt][2]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\r_reg[tfcnt][3]_i_2_n_5 ),
        .I2(\r[tfcnt][7]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r_reg[tfcnt][3]_i_3_n_5 ),
        .O(\r[tfcnt][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44454440)) 
    \r[tfcnt][3]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\r_reg[tfcnt][3]_i_2_n_4 ),
        .I2(\r[tfcnt][7]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r_reg[tfcnt][3]_i_3_n_4 ),
        .O(\r[tfcnt][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9F60)) 
    \r[tfcnt][3]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[txread] ),
        .I1(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I2(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I3(\r[tfcnt][3]_i_20_n_0 ),
        .O(\r[tfcnt][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h96AA)) 
    \r[tfcnt][3]_i_11 
       (.I0(\r[tfcnt][3]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txread] ),
        .I2(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .O(\r[tfcnt][3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h82AA)) 
    \r[tfcnt][3]_i_12 
       (.I0(\r[tfcnt][3]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txread] ),
        .I2(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .O(\r[tfcnt][3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF60)) 
    \r[tfcnt][3]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[txread] ),
        .I1(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I2(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I3(\r[tfcnt][3]_i_7_n_0 ),
        .O(\r[tfcnt][3]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6955)) 
    \r[tfcnt][3]_i_14 
       (.I0(\r[tfcnt][3]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txread] ),
        .I2(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .O(\r[tfcnt][3]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r[tfcnt][3]_i_15 
       (.I0(\r[tfcnt][3]_i_4_n_0 ),
        .I1(\r[tfcnt][7]_i_7_n_0 ),
        .O(\r[tfcnt][3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h82AA7D55)) 
    \r[tfcnt][3]_i_16 
       (.I0(\r[tfcnt][3]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txread] ),
        .I2(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I4(\r[tfcnt][3]_i_4_n_0 ),
        .O(\r[tfcnt][3]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9F6000FF)) 
    \r[tfcnt][3]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[txread] ),
        .I1(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I2(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I3(\r[tfcnt][3]_i_20_n_0 ),
        .I4(\r[tfcnt][3]_i_7_n_0 ),
        .O(\r[tfcnt][3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h96AA)) 
    \r[tfcnt][3]_i_18 
       (.I0(\r[tfcnt][3]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txread] ),
        .I2(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .O(\r[tfcnt][3]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \r[tfcnt][3]_i_19 
       (.I0(\m100.u0/ethc0/r_reg[tfcnt_n_0_][0] ),
        .I1(\a9.x[0].r0_i_34__1_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[tfcnt_n_0_][1] ),
        .O(\r[tfcnt][3]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h74FF740003000300)) 
    \r[tfcnt][3]_i_20 
       (.I0(\r[tfcnt][7]_i_16_n_0 ),
        .I1(\r[tfcnt][7]_i_17_n_0 ),
        .I2(\r[tfcnt][3]_i_21_n_0 ),
        .I3(\r[tfcnt][7]_i_20_n_0 ),
        .I4(\r[tfcnt][7]_i_19_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[tfcnt_n_0_][1] ),
        .O(\r[tfcnt][3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r[tfcnt][3]_i_21 
       (.I0(\a9.x[0].r0_i_34__1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[tfcnt_n_0_][0] ),
        .O(\r[tfcnt][3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h74740303FF000000)) 
    \r[tfcnt][3]_i_4 
       (.I0(\r[tfcnt][7]_i_16_n_0 ),
        .I1(\r[tfcnt][7]_i_17_n_0 ),
        .I2(\r[tfcnt][3]_i_19_n_0 ),
        .I3(\r[tfcnt][7]_i_19_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tfcnt_n_0_][2] ),
        .I5(\r[tfcnt][7]_i_20_n_0 ),
        .O(\r[tfcnt][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h9F)) 
    \r[tfcnt][3]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txread] ),
        .I1(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I2(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .O(\r[tfcnt][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h28)) 
    \r[tfcnt][3]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I2(\m100.u0/ethc0/r_reg[txread] ),
        .O(\r[tfcnt][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4C43CCCC4C430000)) 
    \r[tfcnt][3]_i_7 
       (.I0(\r[tfcnt][7]_i_16_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[tfcnt_n_0_][0] ),
        .I2(\r[tfcnt][7]_i_17_n_0 ),
        .I3(\a9.x[0].r0_i_34__1_n_0 ),
        .I4(\r[tfcnt][7]_i_20_n_0 ),
        .I5(\r[tfcnt][7]_i_19_n_0 ),
        .O(\r[tfcnt][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r[tfcnt][3]_i_8 
       (.I0(\r[tfcnt][3]_i_4_n_0 ),
        .I1(\r[tfcnt][7]_i_7_n_0 ),
        .O(\r[tfcnt][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9F60)) 
    \r[tfcnt][3]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[txread] ),
        .I1(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I2(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I3(\r[tfcnt][3]_i_4_n_0 ),
        .O(\r[tfcnt][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44454440)) 
    \r[tfcnt][4]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\r_reg[tfcnt][7]_i_2_n_7 ),
        .I2(\r[tfcnt][7]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r_reg[tfcnt][7]_i_4_n_7 ),
        .O(\r[tfcnt][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44454440)) 
    \r[tfcnt][5]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\r_reg[tfcnt][7]_i_2_n_6 ),
        .I2(\r[tfcnt][7]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r_reg[tfcnt][7]_i_4_n_6 ),
        .O(\r[tfcnt][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44454440)) 
    \r[tfcnt][6]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\r_reg[tfcnt][7]_i_2_n_5 ),
        .I2(\r[tfcnt][7]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r_reg[tfcnt][7]_i_4_n_5 ),
        .O(\r[tfcnt][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44454440)) 
    \r[tfcnt][7]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\r_reg[tfcnt][7]_i_2_n_4 ),
        .I2(\r[tfcnt][7]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r_reg[tfcnt][7]_i_4_n_4 ),
        .O(\r[tfcnt][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r[tfcnt][7]_i_10 
       (.I0(\r[tfcnt][7]_i_6_n_0 ),
        .I1(\r[tfcnt][7]_i_5_n_0 ),
        .O(\r[tfcnt][7]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r[tfcnt][7]_i_11 
       (.I0(\r[tfcnt][7]_i_7_n_0 ),
        .I1(\r[tfcnt][7]_i_6_n_0 ),
        .O(\r[tfcnt][7]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA5656AAAAA656AA)) 
    \r[tfcnt][7]_i_12 
       (.I0(\r[tfcnt][7]_i_23_n_0 ),
        .I1(\r[tfcnt][7]_i_19_n_0 ),
        .I2(\r[tfcnt][7]_i_20_n_0 ),
        .I3(\r[tfcnt][7]_i_24_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tfcnt_n_0_][7] ),
        .I5(\r[tfcnt][7]_i_25_n_0 ),
        .O(\r[tfcnt][7]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[tfcnt][7]_i_13 
       (.I0(\r[tfcnt][7]_i_5_n_0 ),
        .I1(\r[tfcnt][7]_i_23_n_0 ),
        .O(\r[tfcnt][7]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r[tfcnt][7]_i_14 
       (.I0(\r[tfcnt][7]_i_6_n_0 ),
        .I1(\r[tfcnt][7]_i_5_n_0 ),
        .O(\r[tfcnt][7]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r[tfcnt][7]_i_15 
       (.I0(\r[tfcnt][7]_i_7_n_0 ),
        .I1(\r[tfcnt][7]_i_6_n_0 ),
        .O(\r[tfcnt][7]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6006)) 
    \r[tfcnt][7]_i_16 
       (.I0(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I1(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .O(\r[tfcnt][7]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1001)) 
    \r[tfcnt][7]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[tfcnt][7]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \r[tfcnt][7]_i_18 
       (.I0(\m100.u0/ethc0/r_reg[tfcnt_n_0_][1] ),
        .I1(\a9.x[0].r0_i_34__1_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[tfcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[tfcnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[tfcnt_n_0_][3] ),
        .I5(\m100.u0/ethc0/r_reg[tfcnt_n_0_][4] ),
        .O(\r[tfcnt][7]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFF9FF0FFFF09)) 
    \r[tfcnt][7]_i_19 
       (.I0(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .I1(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[tfcnt][7]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1004)) 
    \r[tfcnt][7]_i_20 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\r[tfcnt][7]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00800000)) 
    \r[tfcnt][7]_i_21 
       (.I0(\m100.u0/ethc0/r_reg[tfcnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[tfcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[tfcnt_n_0_][0] ),
        .I3(\a9.x[0].r0_i_34__1_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tfcnt_n_0_][1] ),
        .O(\r[tfcnt][7]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hDFFF)) 
    \r[tfcnt][7]_i_22 
       (.I0(\m100.u0/ethc0/r_reg[tfcnt_n_0_][1] ),
        .I1(\a9.x[0].r0_i_34__1_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[tfcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[tfcnt_n_0_][2] ),
        .O(\r[tfcnt][7]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555F7FF55FFF7FF)) 
    \r[tfcnt][7]_i_23 
       (.I0(\r[tfcnt][7]_i_26_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[tfcnt_n_0_][5] ),
        .I2(\r[tfcnt][7]_i_27_n_0 ),
        .I3(\r[tfcnt][7]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tfcnt_n_0_][6] ),
        .I5(\r[tfcnt][7]_i_19_n_0 ),
        .O(\r[tfcnt][7]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \r[tfcnt][7]_i_24 
       (.I0(\r[txburstav]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\a9.x[0].r0_i_34__1_n_0 ),
        .O(\r[tfcnt][7]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF6FFFFF6FFFFFFFF)) 
    \r[tfcnt][7]_i_25 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\r[tfwpnt][6]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .I4(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .I5(\r[tfwpnt][6]_i_5_n_0 ),
        .O(\r[tfcnt][7]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFF7FFFF)) 
    \r[tfcnt][7]_i_26 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\r[tfcnt][7]_i_16_n_0 ),
        .I5(\r[tfcnt][7]_i_24_n_0 ),
        .O(\r[tfcnt][7]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF7FFFFFFFFFFFFF)) 
    \r[tfcnt][7]_i_27 
       (.I0(\m100.u0/ethc0/r_reg[tfcnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[tfcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[tfcnt_n_0_][0] ),
        .I3(\r[tfcnt][7]_i_28_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tfcnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[tfcnt_n_0_][4] ),
        .O(\r[tfcnt][7]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF0009)) 
    \r[tfcnt][7]_i_28 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\a9.x[0].r0_i_34__1_n_0 ),
        .O(\r[tfcnt][7]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \r[tfcnt][7]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[tfcnt][7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47473030FF000000)) 
    \r[tfcnt][7]_i_5 
       (.I0(\r[tfcnt][7]_i_16_n_0 ),
        .I1(\r[tfcnt][7]_i_17_n_0 ),
        .I2(\r[tfcnt][7]_i_18_n_0 ),
        .I3(\r[tfcnt][7]_i_19_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tfcnt_n_0_][5] ),
        .I5(\r[tfcnt][7]_i_20_n_0 ),
        .O(\r[tfcnt][7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47473030FF000000)) 
    \r[tfcnt][7]_i_6 
       (.I0(\r[tfcnt][7]_i_16_n_0 ),
        .I1(\r[tfcnt][7]_i_17_n_0 ),
        .I2(\r[tfcnt][7]_i_21_n_0 ),
        .I3(\r[tfcnt][7]_i_19_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tfcnt_n_0_][4] ),
        .I5(\r[tfcnt][7]_i_20_n_0 ),
        .O(\r[tfcnt][7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h74740303FF000000)) 
    \r[tfcnt][7]_i_7 
       (.I0(\r[tfcnt][7]_i_16_n_0 ),
        .I1(\r[tfcnt][7]_i_17_n_0 ),
        .I2(\r[tfcnt][7]_i_22_n_0 ),
        .I3(\r[tfcnt][7]_i_19_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tfcnt_n_0_][3] ),
        .I5(\r[tfcnt][7]_i_20_n_0 ),
        .O(\r[tfcnt][7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA5656AAAAA656AA)) 
    \r[tfcnt][7]_i_8 
       (.I0(\r[tfcnt][7]_i_23_n_0 ),
        .I1(\r[tfcnt][7]_i_19_n_0 ),
        .I2(\r[tfcnt][7]_i_20_n_0 ),
        .I3(\r[tfcnt][7]_i_24_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tfcnt_n_0_][7] ),
        .I5(\r[tfcnt][7]_i_25_n_0 ),
        .O(\r[tfcnt][7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[tfcnt][7]_i_9 
       (.I0(\r[tfcnt][7]_i_5_n_0 ),
        .I1(\r[tfcnt][7]_i_23_n_0 ),
        .O(\r[tfcnt][7]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000440)) 
    \r[tfrpnt][0]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I2(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[txread] ),
        .I4(\m100.u0/txraddress [0]),
        .O(\r[tfrpnt][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000044004400000)) 
    \r[tfrpnt][1]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I2(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[txread] ),
        .I4(\m100.u0/txraddress [1]),
        .I5(\m100.u0/txraddress [0]),
        .O(\r[tfrpnt][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040404040000000)) 
    \r[tfrpnt][2]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I2(\m100.u0/ethc0/v[tfrpnt]1 ),
        .I3(\m100.u0/txraddress [0]),
        .I4(\m100.u0/txraddress [1]),
        .I5(\m100.u0/txraddress [2]),
        .O(\r[tfrpnt][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    \r[tfrpnt][3]_i_1 
       (.I0(\r[tfrpnt][4]_i_2_n_0 ),
        .I1(\m100.u0/txraddress [1]),
        .I2(\m100.u0/txraddress [0]),
        .I3(\m100.u0/txraddress [2]),
        .I4(\m100.u0/txraddress [3]),
        .O(\r[tfrpnt][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2AAAAAAA80000000)) 
    \r[tfrpnt][4]_i_1 
       (.I0(\r[tfrpnt][4]_i_2_n_0 ),
        .I1(\m100.u0/txraddress [2]),
        .I2(\m100.u0/txraddress [0]),
        .I3(\m100.u0/txraddress [1]),
        .I4(\m100.u0/txraddress [3]),
        .I5(\m100.u0/txraddress [4]),
        .O(\r[tfrpnt][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0060)) 
    \r[tfrpnt][4]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txread] ),
        .I1(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I2(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I3(\r[abufs][2]_i_6_n_0 ),
        .O(\r[tfrpnt][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000044004400000)) 
    \r[tfrpnt][5]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I2(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[txread] ),
        .I4(\r[tfrpnt][5]_i_2_n_0 ),
        .I5(\m100.u0/txraddress [5]),
        .O(\r[tfrpnt][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \r[tfrpnt][5]_i_2 
       (.I0(\m100.u0/txraddress [3]),
        .I1(\m100.u0/txraddress [1]),
        .I2(\m100.u0/txraddress [0]),
        .I3(\m100.u0/txraddress [2]),
        .I4(\m100.u0/txraddress [4]),
        .O(\r[tfrpnt][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFBEAA)) 
    \r[tfrpnt][6]_i_1 
       (.I0(\r[tfrpnt][6]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txread] ),
        .I2(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I4(\m100.u0/ethc0/rin[status][txahberr] ),
        .I5(\r[abufs][2]_i_6_n_0 ),
        .O(\r[tfrpnt][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000006600000)) 
    \r[tfrpnt][6]_i_2 
       (.I0(\m100.u0/txraddress [6]),
        .I1(\r[tfrpnt][6]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txread] ),
        .I3(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .I4(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I5(\r[abufs][2]_i_6_n_0 ),
        .O(\r[tfrpnt][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000D05555D0)) 
    \r[tfrpnt][6]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\r[tfwpnt][6]_i_5_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .I4(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .I5(\r[tfwpnt][6]_i_3_n_0 ),
        .O(\r[tfrpnt][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \r[tfrpnt][6]_i_4 
       (.I0(\m100.u0/txraddress [4]),
        .I1(\m100.u0/txraddress [2]),
        .I2(\m100.u0/txraddress [0]),
        .I3(\m100.u0/txraddress [1]),
        .I4(\m100.u0/txraddress [3]),
        .I5(\m100.u0/txraddress [5]),
        .O(\r[tfrpnt][6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \r[tfwpnt][0]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/txwaddress [0]),
        .O(\m100.u0/ethc0/v[tfwpnt] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT4 #(
    .INIT(16'h0220)) 
    \r[tfwpnt][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/txwaddress [1]),
        .I3(\m100.u0/txwaddress [0]),
        .O(\m100.u0/ethc0/v[tfwpnt] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT5 #(
    .INIT(32'h04404040)) 
    \r[tfwpnt][2]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/txwaddress [2]),
        .I3(\m100.u0/txwaddress [1]),
        .I4(\m100.u0/txwaddress [0]),
        .O(\r[tfwpnt][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0440404040404040)) 
    \r[tfwpnt][3]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/txwaddress [3]),
        .I3(\m100.u0/txwaddress [2]),
        .I4(\m100.u0/txwaddress [0]),
        .I5(\m100.u0/txwaddress [1]),
        .O(\r[tfwpnt][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2888888888888888)) 
    \r[tfwpnt][4]_i_1 
       (.I0(\r[tfwpnt][4]_i_2_n_0 ),
        .I1(\m100.u0/txwaddress [4]),
        .I2(\m100.u0/txwaddress [2]),
        .I3(\m100.u0/txwaddress [0]),
        .I4(\m100.u0/txwaddress [1]),
        .I5(\m100.u0/txwaddress [3]),
        .O(\m100.u0/ethc0/v[tfwpnt] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[tfwpnt][4]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[tfwpnt][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT4 #(
    .INIT(16'h0220)) 
    \r[tfwpnt][5]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/txwaddress [5]),
        .I3(\r[tfwpnt][6]_i_7_n_0 ),
        .O(\m100.u0/ethc0/v[tfwpnt] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF10005454)) 
    \r[tfwpnt][6]_i_1 
       (.I0(\r[tfwpnt][6]_i_3_n_0 ),
        .I1(\r[tfwpnt][6]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\r[tfwpnt][6]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\r[tfwpnt][6]_i_6_n_0 ),
        .O(\r[tfwpnt][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT5 #(
    .INIT(32'h14440000)) 
    \r[tfwpnt][6]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/txwaddress [6]),
        .I2(\m100.u0/txwaddress [5]),
        .I3(\r[tfwpnt][6]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[tfwpnt][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r[tfwpnt][6]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[tfwpnt][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[tfwpnt][6]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .I1(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .O(\r[tfwpnt][6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[tfwpnt][6]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I1(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .O(\r[tfwpnt][6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h03C000C030103010)) 
    \r[tfwpnt][6]_i_6 
       (.I0(\a9.x[0].r0_i_34__1_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r[tfwpnt][6]_i_5_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[tfwpnt][6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \r[tfwpnt][6]_i_7 
       (.I0(\m100.u0/txwaddress [3]),
        .I1(\m100.u0/txwaddress [1]),
        .I2(\m100.u0/txwaddress [0]),
        .I3(\m100.u0/txwaddress [2]),
        .I4(\m100.u0/txwaddress [4]),
        .O(\r[tfwpnt][6]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][13]_i_10 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [12]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][13]_i_14_n_6 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [4]),
        .O(\r[tmsto][addr][13]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][13]_i_11 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][13]_i_14_n_6 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdesc]__0 [4]),
        .I5(\r[tmsto][addr][13]_i_17_n_0 ),
        .O(\r[tmsto][addr][13]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][13]_i_12 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [11]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][13]_i_14_n_7 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [3]),
        .O(\r[tmsto][addr][13]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][13]_i_13 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][13]_i_14_n_7 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdesc]__0 [3]),
        .I5(\r[tmsto][addr][13]_i_18_n_0 ),
        .O(\r[tmsto][addr][13]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][13]_i_15 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [14]),
        .O(\r[tmsto][addr][13]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][13]_i_16 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdesc]__0 [5]),
        .I2(\r_reg[tmsto][addr][13]_i_14_n_5 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][13]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][13]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [12]),
        .O(\r[tmsto][addr][13]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][13]_i_18 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [11]),
        .O(\r[tmsto][addr][13]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][13]_i_2 
       (.I0(\r[tmsto][addr][13]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][13]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [16]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][13]_i_3 
       (.I0(\r[tmsto][addr][13]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][13]_i_9_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [15]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][13]_i_4 
       (.I0(\r[tmsto][addr][13]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][13]_i_11_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [14]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][13]_i_5 
       (.I0(\r[tmsto][addr][13]_i_12_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][13]_i_13_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [13]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][13]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][13]_i_6 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [14]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][13]_i_14_n_4 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [6]),
        .O(\r[tmsto][addr][13]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][13]_i_7 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][13]_i_14_n_4 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdesc]__0 [6]),
        .I5(\r[tmsto][addr][13]_i_15_n_0 ),
        .O(\r[tmsto][addr][13]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][13]_i_8 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [13]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][13]_i_14_n_5 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [5]),
        .O(\r[tmsto][addr][13]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF8080F000)) 
    \r[tmsto][addr][13]_i_9 
       (.I0(\m100.u0/ethc0/tmsti ),
        .I1(\r_reg[tmsto][addr][13]_i_14_n_5 ),
        .I2(\r[tmsto][addr][1]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txaddr]__0 [13]),
        .I4(\r[tmsto][data][31]_i_5_n_0 ),
        .I5(\r[tmsto][addr][13]_i_16_n_0 ),
        .O(\r[tmsto][addr][13]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][17]_i_10 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [16]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][17]_i_14_n_6 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [8]),
        .O(\r[tmsto][addr][17]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][17]_i_11 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][17]_i_14_n_6 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdesc]__0 [8]),
        .I5(\r[tmsto][addr][17]_i_17_n_0 ),
        .O(\r[tmsto][addr][17]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][17]_i_12 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [15]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][17]_i_14_n_7 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [7]),
        .O(\r[tmsto][addr][17]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][17]_i_13 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][17]_i_14_n_7 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdesc]__0 [7]),
        .I5(\r[tmsto][addr][17]_i_18_n_0 ),
        .O(\r[tmsto][addr][17]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][17]_i_15 
       (.I0(\r[tmsto][addr][1]_i_27_n_0 ),
        .I1(\r_reg[tmsto][addr][17]_i_14_n_4 ),
        .I2(\m100.u0/ethc0/r_reg[txdesc]__0 [10]),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][17]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][17]_i_16 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [17]),
        .O(\r[tmsto][addr][17]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][17]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [16]),
        .O(\r[tmsto][addr][17]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][17]_i_18 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [15]),
        .O(\r[tmsto][addr][17]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][17]_i_2 
       (.I0(\r[tmsto][addr][17]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][17]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [20]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][17]_i_3 
       (.I0(\r[tmsto][addr][17]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][17]_i_9_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [19]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][17]_i_4 
       (.I0(\r[tmsto][addr][17]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][17]_i_11_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [18]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][17]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][17]_i_5 
       (.I0(\r[tmsto][addr][17]_i_12_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][17]_i_13_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [17]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][17]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][17]_i_6 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [18]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][17]_i_14_n_4 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [10]),
        .O(\r[tmsto][addr][17]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF80AA8000)) 
    \r[tmsto][addr][17]_i_7 
       (.I0(\r[tmsto][addr][1]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/tmsti ),
        .I2(\r_reg[tmsto][addr][17]_i_14_n_4 ),
        .I3(\r[tmsto][data][31]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [18]),
        .I5(\r[tmsto][addr][17]_i_15_n_0 ),
        .O(\r[tmsto][addr][17]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][17]_i_8 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [17]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][17]_i_14_n_5 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [9]),
        .O(\r[tmsto][addr][17]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][17]_i_9 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][17]_i_14_n_5 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdesc]__0 [9]),
        .I5(\r[tmsto][addr][17]_i_16_n_0 ),
        .O(\r[tmsto][addr][17]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFEEEE)) 
    \r[tmsto][addr][1]_i_1 
       (.I0(\r[tmsto][addr][1]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/tmsti[retry] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/tmsti ),
        .I4(\r[tmsto][addr][1]_i_5_n_0 ),
        .I5(\r[tmsto][addr][1]_i_6_n_0 ),
        .O(\r[tmsto][addr][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF044)) 
    \r[tmsto][addr][1]_i_10 
       (.I0(\r[tmsto][addr][1]_i_18_n_0 ),
        .I1(\r_reg[tmsto][addr][1]_i_17_n_7 ),
        .I2(\m100.u0/ethc0/r_reg[tmsto][addr] [1]),
        .I3(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FEFFFF)) 
    \r[tmsto][addr][1]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[abufs_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg ),
        .I3(\m100.u0/ethc0/p_6_in [14]),
        .I4(\m100.u0/ethc0/p_6_in [0]),
        .O(\r[tmsto][addr][1]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][1]_i_12 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [2]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][1]_i_17_n_4 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdsel_n_0_][4] ),
        .O(\r[tmsto][addr][1]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][1]_i_13 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][1]_i_17_n_4 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdsel_n_0_][4] ),
        .I5(\r[tmsto][addr][1]_i_21_n_0 ),
        .O(\r[tmsto][addr][1]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][1]_i_14 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [1]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][1]_i_17_n_5 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdsel_n_0_][3] ),
        .O(\r[tmsto][addr][1]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF80AA8000)) 
    \r[tmsto][addr][1]_i_15 
       (.I0(\r[tmsto][addr][1]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/tmsti ),
        .I2(\r_reg[tmsto][addr][1]_i_17_n_5 ),
        .I3(\r[tmsto][data][31]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [1]),
        .I5(\r[tmsto][addr][1]_i_22_n_0 ),
        .O(\r[tmsto][addr][1]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFDFFFF5FFDF)) 
    \r[tmsto][addr][1]_i_16 
       (.I0(\m100.u0/ethc0/r_reg[txaddr]__0 [0]),
        .I1(\r_reg[tmsto][write]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\r[tmsto][addr][1]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFDFFF00F)) 
    \r[tmsto][addr][1]_i_18 
       (.I0(\m100.u0/ethc0/tmsti ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[tmsto][addr][1]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF7CCFF)) 
    \r[tmsto][addr][1]_i_19 
       (.I0(\m100.u0/ethc0/tmsti ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[tmsto][addr][1]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFBFF)) 
    \r[tmsto][addr][1]_i_20 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[tmsto][addr][1]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][1]_i_21 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [2]),
        .O(\r[tmsto][addr][1]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][1]_i_22 
       (.I0(\r[tmsto][addr][1]_i_27_n_0 ),
        .I1(\r_reg[tmsto][addr][1]_i_17_n_5 ),
        .I2(\m100.u0/ethc0/r_reg[txdsel_n_0_][3] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][1]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \r[tmsto][addr][1]_i_25 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [2]),
        .O(\r[tmsto][addr][1]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \r[tmsto][addr][1]_i_27 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[tmsto][addr][1]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3033301130003011)) 
    \r[tmsto][addr][1]_i_3 
       (.I0(\r[tmsto][addr][1]_i_11_n_0 ),
        .I1(\r[txcnt][10]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/tmsti ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[txden]__0 ),
        .O(\r[tmsto][addr][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0080008000000080)) 
    \r[tmsto][addr][1]_i_4 
       (.I0(\ahbmi[hready] ),
        .I1(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I2(\m100.u0/ethc0/ahb0/r_reg[bg]__0 ),
        .I3(\m100.u0/ethc0/ahb0/r_reg[retry]__0 ),
        .I4(\m100.u0/ethc0/r_reg[rmsto][req_n_0_] ),
        .I5(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\m100.u0/ethc0/tmsti ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \r[tmsto][addr][1]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[tmsto][addr][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000B800)) 
    \r[tmsto][addr][1]_i_6 
       (.I0(\r[tfwpnt][6]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/tmsti ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[tmsto][addr][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][1]_i_7 
       (.I0(\r[tmsto][addr][1]_i_12_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][1]_i_13_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [4]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][1]_i_8 
       (.I0(\r[tmsto][addr][1]_i_14_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][1]_i_15_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [3]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FF5D5D)) 
    \r[tmsto][addr][1]_i_9 
       (.I0(\r[tmsto][addr][1]_i_16_n_0 ),
        .I1(\r_reg[tmsto][addr][1]_i_17_n_6 ),
        .I2(\r[tmsto][addr][1]_i_18_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[tmsto][addr] [2]),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][21]_i_10 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [20]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][21]_i_14_n_6 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [12]),
        .O(\r[tmsto][addr][21]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][21]_i_11 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][21]_i_14_n_6 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdesc]__0 [12]),
        .I5(\r[tmsto][addr][21]_i_17_n_0 ),
        .O(\r[tmsto][addr][21]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][21]_i_12 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [19]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][21]_i_14_n_7 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [11]),
        .O(\r[tmsto][addr][21]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF8080F000)) 
    \r[tmsto][addr][21]_i_13 
       (.I0(\m100.u0/ethc0/tmsti ),
        .I1(\r_reg[tmsto][addr][21]_i_14_n_7 ),
        .I2(\r[tmsto][addr][1]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txaddr]__0 [19]),
        .I4(\r[tmsto][data][31]_i_5_n_0 ),
        .I5(\r[tmsto][addr][21]_i_18_n_0 ),
        .O(\r[tmsto][addr][21]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][21]_i_15 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdesc]__0 [14]),
        .I2(\r_reg[tmsto][addr][21]_i_14_n_4 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][21]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][21]_i_16 
       (.I0(\r[tmsto][addr][1]_i_27_n_0 ),
        .I1(\r_reg[tmsto][addr][21]_i_14_n_5 ),
        .I2(\m100.u0/ethc0/r_reg[txdesc]__0 [13]),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][21]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][21]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [20]),
        .O(\r[tmsto][addr][21]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][21]_i_18 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdesc]__0 [11]),
        .I2(\r_reg[tmsto][addr][21]_i_14_n_7 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][21]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][21]_i_2 
       (.I0(\r[tmsto][addr][21]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][21]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [24]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][21]_i_3 
       (.I0(\r[tmsto][addr][21]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][21]_i_9_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [23]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][21]_i_4 
       (.I0(\r[tmsto][addr][21]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][21]_i_11_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [22]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][21]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][21]_i_5 
       (.I0(\r[tmsto][addr][21]_i_12_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][21]_i_13_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [21]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][21]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][21]_i_6 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [22]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][21]_i_14_n_4 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [14]),
        .O(\r[tmsto][addr][21]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF80AA8000)) 
    \r[tmsto][addr][21]_i_7 
       (.I0(\r[tmsto][addr][1]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/tmsti ),
        .I2(\r_reg[tmsto][addr][21]_i_14_n_4 ),
        .I3(\r[tmsto][data][31]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [22]),
        .I5(\r[tmsto][addr][21]_i_15_n_0 ),
        .O(\r[tmsto][addr][21]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][21]_i_8 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [21]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][21]_i_14_n_5 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [13]),
        .O(\r[tmsto][addr][21]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF80AA8000)) 
    \r[tmsto][addr][21]_i_9 
       (.I0(\r[tmsto][addr][1]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/tmsti ),
        .I2(\r_reg[tmsto][addr][21]_i_14_n_5 ),
        .I3(\r[tmsto][data][31]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [21]),
        .I5(\r[tmsto][addr][21]_i_16_n_0 ),
        .O(\r[tmsto][addr][21]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][25]_i_10 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [24]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][25]_i_14_n_6 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [16]),
        .O(\r[tmsto][addr][25]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][25]_i_11 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][25]_i_14_n_6 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdesc]__0 [16]),
        .I5(\r[tmsto][addr][25]_i_17_n_0 ),
        .O(\r[tmsto][addr][25]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][25]_i_12 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [23]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][25]_i_14_n_7 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [15]),
        .O(\r[tmsto][addr][25]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF80AA8000)) 
    \r[tmsto][addr][25]_i_13 
       (.I0(\r[tmsto][addr][1]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/tmsti ),
        .I2(\r_reg[tmsto][addr][25]_i_14_n_7 ),
        .I3(\r[tmsto][data][31]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [23]),
        .I5(\r[tmsto][addr][25]_i_18_n_0 ),
        .O(\r[tmsto][addr][25]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][25]_i_15 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [26]),
        .O(\r[tmsto][addr][25]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][25]_i_16 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdesc]__0 [17]),
        .I2(\r_reg[tmsto][addr][25]_i_14_n_5 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][25]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][25]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [24]),
        .O(\r[tmsto][addr][25]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][25]_i_18 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdesc]__0 [15]),
        .I2(\r_reg[tmsto][addr][25]_i_14_n_7 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][25]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][25]_i_2 
       (.I0(\r[tmsto][addr][25]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][25]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [28]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][25]_i_3 
       (.I0(\r[tmsto][addr][25]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][25]_i_9_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [27]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][25]_i_4 
       (.I0(\r[tmsto][addr][25]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][25]_i_11_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [26]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][25]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][25]_i_5 
       (.I0(\r[tmsto][addr][25]_i_12_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][25]_i_13_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [25]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][25]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][25]_i_6 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [26]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][25]_i_14_n_4 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [18]),
        .O(\r[tmsto][addr][25]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][25]_i_7 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][25]_i_14_n_4 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdesc]__0 [18]),
        .I5(\r[tmsto][addr][25]_i_15_n_0 ),
        .O(\r[tmsto][addr][25]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][25]_i_8 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [25]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][25]_i_14_n_5 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [17]),
        .O(\r[tmsto][addr][25]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF8080F000)) 
    \r[tmsto][addr][25]_i_9 
       (.I0(\m100.u0/ethc0/tmsti ),
        .I1(\r_reg[tmsto][addr][25]_i_14_n_5 ),
        .I2(\r[tmsto][addr][1]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txaddr]__0 [25]),
        .I4(\r[tmsto][data][31]_i_5_n_0 ),
        .I5(\r[tmsto][addr][25]_i_16_n_0 ),
        .O(\r[tmsto][addr][25]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][29]_i_10 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][29]_i_11_n_7 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdesc]__0 [19]),
        .I5(\r[tmsto][addr][29]_i_14_n_0 ),
        .O(\r[tmsto][addr][29]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][29]_i_12 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdesc]__0 [21]),
        .I2(\r_reg[tmsto][addr][29]_i_11_n_5 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][29]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][29]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [28]),
        .O(\r[tmsto][addr][29]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][29]_i_14 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [27]),
        .O(\r[tmsto][addr][29]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7070707770707070)) 
    \r[tmsto][addr][29]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][addr] [31]),
        .I1(\m100.u0/ethc0/tmsti[retry] ),
        .I2(\r[tmsto][addr][29]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\r[tmsto][addr][29]_i_6_n_0 ),
        .O(\r[tmsto][addr][29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][29]_i_3 
       (.I0(\r[tmsto][addr][29]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][29]_i_8_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [30]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][29]_i_4 
       (.I0(\r[tmsto][addr][29]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][29]_i_10_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [29]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][29]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF8080F000)) 
    \r[tmsto][addr][29]_i_5 
       (.I0(\m100.u0/ethc0/tmsti ),
        .I1(\r_reg[tmsto][addr][29]_i_11_n_5 ),
        .I2(\r[tmsto][addr][1]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txaddr]__0 [29]),
        .I4(\r[tmsto][data][31]_i_5_n_0 ),
        .I5(\r[tmsto][addr][29]_i_12_n_0 ),
        .O(\r[tmsto][addr][29]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][29]_i_6 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [29]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][29]_i_11_n_5 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [21]),
        .O(\r[tmsto][addr][29]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][29]_i_7 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [28]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][29]_i_11_n_6 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [20]),
        .O(\r[tmsto][addr][29]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][29]_i_8 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][29]_i_11_n_6 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdesc]__0 [20]),
        .I5(\r[tmsto][addr][29]_i_13_n_0 ),
        .O(\r[tmsto][addr][29]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][29]_i_9 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [27]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][29]_i_11_n_7 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [19]),
        .O(\r[tmsto][addr][29]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][5]_i_10 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [4]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][5]_i_14_n_6 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdsel_n_0_][6] ),
        .O(\r[tmsto][addr][5]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF80AA8000)) 
    \r[tmsto][addr][5]_i_11 
       (.I0(\r[tmsto][addr][1]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/tmsti ),
        .I2(\r_reg[tmsto][addr][5]_i_14_n_6 ),
        .I3(\r[tmsto][data][31]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [4]),
        .I5(\r[tmsto][addr][5]_i_17_n_0 ),
        .O(\r[tmsto][addr][5]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][5]_i_12 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [3]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][5]_i_14_n_7 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdsel_n_0_][5] ),
        .O(\r[tmsto][addr][5]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF80AA8000)) 
    \r[tmsto][addr][5]_i_13 
       (.I0(\r[tmsto][addr][1]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/tmsti ),
        .I2(\r_reg[tmsto][addr][5]_i_14_n_7 ),
        .I3(\r[tmsto][data][31]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [3]),
        .I5(\r[tmsto][addr][5]_i_18_n_0 ),
        .O(\r[tmsto][addr][5]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[tmsto][addr][5]_i_15 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [6]),
        .O(\r[tmsto][addr][5]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][5]_i_16 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdsel_n_0_][7] ),
        .I2(\r_reg[tmsto][addr][5]_i_14_n_5 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][5]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][5]_i_17 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdsel_n_0_][6] ),
        .I2(\r_reg[tmsto][addr][5]_i_14_n_6 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][5]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][5]_i_18 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdsel_n_0_][5] ),
        .I2(\r_reg[tmsto][addr][5]_i_14_n_7 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][5]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][5]_i_2 
       (.I0(\r[tmsto][addr][5]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][5]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [8]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][5]_i_3 
       (.I0(\r[tmsto][addr][5]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][5]_i_9_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [7]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][5]_i_4 
       (.I0(\r[tmsto][addr][5]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][5]_i_11_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [6]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][5]_i_5 
       (.I0(\r[tmsto][addr][5]_i_12_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][5]_i_13_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [5]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][5]_i_6 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [6]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][5]_i_14_n_4 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdsel_n_0_][8] ),
        .O(\r[tmsto][addr][5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF4FFF4F4)) 
    \r[tmsto][addr][5]_i_7 
       (.I0(\r[tmsto][addr][1]_i_19_n_0 ),
        .I1(\r_reg[tmsto][addr][5]_i_14_n_4 ),
        .I2(\m100.u0/ethc0/tmsti[retry] ),
        .I3(\r[tmsto][addr][1]_i_20_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdsel_n_0_][8] ),
        .I5(\r[tmsto][addr][5]_i_15_n_0 ),
        .O(\r[tmsto][addr][5]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][5]_i_8 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [5]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][5]_i_14_n_5 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdsel_n_0_][7] ),
        .O(\r[tmsto][addr][5]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF8080F000)) 
    \r[tmsto][addr][5]_i_9 
       (.I0(\m100.u0/ethc0/tmsti ),
        .I1(\r_reg[tmsto][addr][5]_i_14_n_5 ),
        .I2(\r[tmsto][addr][1]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txaddr]__0 [5]),
        .I4(\r[tmsto][data][31]_i_5_n_0 ),
        .I5(\r[tmsto][addr][5]_i_16_n_0 ),
        .O(\r[tmsto][addr][5]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][9]_i_10 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [8]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][9]_i_14_n_6 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [0]),
        .O(\r[tmsto][addr][9]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF80AA8000)) 
    \r[tmsto][addr][9]_i_11 
       (.I0(\r[tmsto][addr][1]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/tmsti ),
        .I2(\r_reg[tmsto][addr][9]_i_14_n_6 ),
        .I3(\r[tmsto][data][31]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [8]),
        .I5(\r[tmsto][addr][9]_i_17_n_0 ),
        .O(\r[tmsto][addr][9]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][9]_i_12 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [7]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][9]_i_14_n_7 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdsel_n_0_][9] ),
        .O(\r[tmsto][addr][9]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF80AA8000)) 
    \r[tmsto][addr][9]_i_13 
       (.I0(\r[tmsto][addr][1]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/tmsti ),
        .I2(\r_reg[tmsto][addr][9]_i_14_n_7 ),
        .I3(\r[tmsto][data][31]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txaddr]__0 [7]),
        .I5(\r[tmsto][addr][9]_i_18_n_0 ),
        .O(\r[tmsto][addr][9]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][9]_i_15 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdesc]__0 [2]),
        .I2(\r_reg[tmsto][addr][9]_i_14_n_4 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][9]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][9]_i_16 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdesc]__0 [1]),
        .I2(\r_reg[tmsto][addr][9]_i_14_n_5 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][9]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][9]_i_17 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdesc]__0 [0]),
        .I2(\r_reg[tmsto][addr][9]_i_14_n_6 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][9]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF44F4)) 
    \r[tmsto][addr][9]_i_18 
       (.I0(\r[tmsto][addr][1]_i_20_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdsel_n_0_][9] ),
        .I2(\r_reg[tmsto][addr][9]_i_14_n_7 ),
        .I3(\r[tmsto][addr][1]_i_27_n_0 ),
        .I4(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][9]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][9]_i_2 
       (.I0(\r[tmsto][addr][9]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][9]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [12]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][9]_i_3 
       (.I0(\r[tmsto][addr][9]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][9]_i_9_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [11]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][9]_i_4 
       (.I0(\r[tmsto][addr][9]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][9]_i_11_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [10]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FDFFFFFF02FF02)) 
    \r[tmsto][addr][9]_i_5 
       (.I0(\r[tmsto][addr][9]_i_12_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[tmsto][addr][9]_i_13_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][addr] [9]),
        .I5(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][addr][9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][9]_i_6 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [10]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][9]_i_14_n_4 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [2]),
        .O(\r[tmsto][addr][9]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF8080F000)) 
    \r[tmsto][addr][9]_i_7 
       (.I0(\m100.u0/ethc0/tmsti ),
        .I1(\r_reg[tmsto][addr][9]_i_14_n_4 ),
        .I2(\r[tmsto][addr][1]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txaddr]__0 [10]),
        .I4(\r[tmsto][data][31]_i_5_n_0 ),
        .I5(\r[tmsto][addr][9]_i_15_n_0 ),
        .O(\r[tmsto][addr][9]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEF4F404040)) 
    \r[tmsto][addr][9]_i_8 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txaddr]__0 [9]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r_reg[tmsto][addr][9]_i_14_n_5 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdesc]__0 [1]),
        .O(\r[tmsto][addr][9]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF8080F000)) 
    \r[tmsto][addr][9]_i_9 
       (.I0(\m100.u0/ethc0/tmsti ),
        .I1(\r_reg[tmsto][addr][9]_i_14_n_5 ),
        .I2(\r[tmsto][addr][1]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txaddr]__0 [9]),
        .I4(\r[tmsto][data][31]_i_5_n_0 ),
        .I5(\r[tmsto][addr][9]_i_16_n_0 ),
        .O(\r[tmsto][addr][9]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F44FFFF4F440000)) 
    \r[tmsto][data][14]_i_1 
       (.I0(\r[tmsto][data][14]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\r[tmsto][data][31]_i_3_n_0 ),
        .I3(\m100.u0/erdata [14]),
        .I4(\m100.u0/ethc0/v[tmsto][data] ),
        .I5(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][14] ),
        .O(\r[tmsto][data][14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h14D7)) 
    \r[tmsto][data][14]_i_2 
       (.I0(\m100.u0/ethc0/txo[status] [0]),
        .I1(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[txstatus_n_0_][0] ),
        .O(\r[tmsto][data][14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F44FFFF4F440000)) 
    \r[tmsto][data][15]_i_1 
       (.I0(\r[tmsto][data][15]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\r[tmsto][data][31]_i_3_n_0 ),
        .I3(\m100.u0/erdata [15]),
        .I4(\m100.u0/ethc0/v[tmsto][data] ),
        .I5(\m100.u0/ethc0/r_reg[tmsto][data_n_0_][15] ),
        .O(\r[tmsto][data][15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h14D7)) 
    \r[tmsto][data][15]_i_2 
       (.I0(\m100.u0/ethc0/txo[status] [1]),
        .I1(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[txstatus_n_0_][1] ),
        .O(\r[tmsto][data][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[tmsto][data][31]_i_1 
       (.I0(\r[tmsto][data][31]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/v[tmsto][data] ),
        .O(\r[tmsto][data][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0024FFFF)) 
    \r[tmsto][data][31]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\r[tmsto][data][31]_i_4_n_0 ),
        .I4(\r[tmsto][data][31]_i_3_n_0 ),
        .O(\m100.u0/ethc0/v[tmsto][data] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hD8DDFFFF)) 
    \r[tmsto][data][31]_i_3 
       (.I0(\r[tmsto][data][31]_i_5_n_0 ),
        .I1(\r[tmsto][data][31]_i_6_n_0 ),
        .I2(\r[txdstate][1]_i_6_n_0 ),
        .I3(\r[tedcl]_i_2_n_0 ),
        .I4(\r[tmsto][addr][1]_i_5_n_0 ),
        .O(\r[tmsto][data][31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF99990FFF)) 
    \r[tmsto][data][31]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I1(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[txden]__0 ),
        .I3(\r_reg[tmsto][write]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[tmsto][data][31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBA)) 
    \r[tmsto][data][31]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\r[tmsto][data][31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF7FF)) 
    \r[tmsto][data][31]_i_6 
       (.I0(\m100.u0/ethc0/ahb0/r_reg ),
        .I1(\ahbmi[hready] ),
        .I2(\ahbmi[hresp] [1]),
        .I3(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .O(\r[tmsto][data][31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFECCCE)) 
    \r[tmsto][req]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I1(\m100.u0/ethc0/tmsti[retry] ),
        .I2(\r[tmsto][req]_i_2_n_0 ),
        .I3(\r[tmsto][req]_i_3_n_0 ),
        .I4(\r[tmsto][req]_i_4_n_0 ),
        .I5(\m100.u0/ethc0/rin[tmsto][req] ),
        .O(\r[tmsto][req]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFDDDFFFFF)) 
    \r[tmsto][req]_i_10 
       (.I0(\r[tmsto][req]_i_16_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I3(\m100.u0/ethc0/r_reg[txburstav]__0 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[tmsto][req]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF200)) 
    \r[tmsto][req]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/tmsti[retry] ),
        .O(\r[tmsto][req]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF2FF)) 
    \r[tmsto][req]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\r[tedcl]_i_2_n_0 ),
        .O(\r[tmsto][req]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF0F0F0F0F8F0F8)) 
    \r[tmsto][req]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\r_reg[tmsto][write]_i_2_n_0 ),
        .I2(\r[tmsto][req]_i_17_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\r[tfwpnt][6]_i_5_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[tmsto][req]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r[tmsto][req]_i_14 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[tmsto][req]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFB2220FFFFFFFF)) 
    \r[tmsto][req]_i_15 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/tmsti[ready] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I5(\r[txcnt][6]_i_8_n_0 ),
        .O(\r[tmsto][req]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h90000090)) 
    \r[tmsto][req]_i_16 
       (.I0(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I1(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .I4(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .O(\r[tmsto][req]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE000E00FE000E000)) 
    \r[tmsto][req]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[txburstav]__0 ),
        .I1(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\m100.u0/ethc0/p_6_in [0]),
        .O(\r[tmsto][req]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555544454445444)) 
    \r[tmsto][req]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\r[tmsto][req]_i_5_n_0 ),
        .I2(\r[tmsto][req]_i_6_n_0 ),
        .I3(\m100.u0/ethc0/p_6_in [0]),
        .I4(\m100.u0/ethc0/tmsti ),
        .I5(\r[tmsto][req]_i_7_n_0 ),
        .O(\r[tmsto][req]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF5454FF54)) 
    \r[tmsto][req]_i_3 
       (.I0(\r[tmsto][req]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/tmsti[retry] ),
        .I2(\r[tmsto][req]_i_9_n_0 ),
        .I3(\r[txstart_sync]_i_3_n_0 ),
        .I4(\r[tmsto][req]_i_10_n_0 ),
        .I5(\r[tmsto][write]_i_4_n_0 ),
        .O(\r[tmsto][req]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF3FFFFFF000F050)) 
    \r[tmsto][req]_i_4 
       (.I0(\r[txdstate][1]_i_6_n_0 ),
        .I1(\r[tmsto][req]_i_9_n_0 ),
        .I2(\r[tmsto][addr][1]_i_5_n_0 ),
        .I3(\r[tmsto][req]_i_11_n_0 ),
        .I4(\r[tmsto][req]_i_12_n_0 ),
        .I5(\r[tmsto][req]_i_13_n_0 ),
        .O(\r[tmsto][req]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00280000)) 
    \r[tmsto][req]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\r[tmsto][req]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111100000001)) 
    \r[tmsto][req]_i_6 
       (.I0(\r[tmsto][req]_i_14_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[abufs_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[abufs_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg ),
        .I5(\m100.u0/ethc0/p_6_in [14]),
        .O(\r[tmsto][req]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000F0000F070F050)) 
    \r[tmsto][req]_i_7 
       (.I0(\r[tmsto][req]_i_15_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txburstcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txburstcnt_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\r[tmsto][req]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFF08FFFFFFFF)) 
    \r[tmsto][req]_i_8 
       (.I0(\r[tedcl]_i_2_n_0 ),
        .I1(\r[txdstate][1]_i_6_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[tmsto][req]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4444FF4F)) 
    \r[tmsto][req]_i_9 
       (.I0(\r[tmsto][req]_i_15_n_0 ),
        .I1(\m100.u0/ethc0/tmsti ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[tmsto][req]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88808080)) 
    \r[tmsto][write]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txlength_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txlength_n_0_][1] ),
        .O(\r[tmsto][write]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBB0B0BBB)) 
    \r[tmsto][write]_i_3 
       (.I0(\r[txdstate][1]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I4(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .O(\r[tmsto][write]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \r[tmsto][write]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\r_reg[tmsto][write]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txden]__0 ),
        .O(\r[tmsto][write]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000112210001133)) 
    \r[tmsto][write]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\r[tfwpnt][6]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\r[tmsto][addr][1]_i_11_n_0 ),
        .O(\r[tmsto][write]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \r[tmsto][write]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txlength_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[txlength_n_0_][4] ),
        .I5(\r[tmsto][write]_i_8_n_0 ),
        .O(\r[tmsto][write]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEAAAAAAA)) 
    \r[tmsto][write]_i_7 
       (.I0(\r[tmsto][write]_i_9_n_0 ),
        .I1(\r[tmsto][write]_i_10_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][8] ),
        .I3(\m100.u0/ethc0/r_reg[txlength_n_0_][6] ),
        .I4(\m100.u0/ethc0/r_reg[txlength_n_0_][5] ),
        .O(\r[tmsto][write]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \r[tmsto][write]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][6] ),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][7] ),
        .I3(\m100.u0/ethc0/r_reg[txlength_n_0_][9] ),
        .I4(\m100.u0/ethc0/r_reg[txlength_n_0_][8] ),
        .O(\r[tmsto][write]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAAAAAAAAAAAAAAA)) 
    \r[tmsto][write]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][9] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[txlength_n_0_][6] ),
        .I4(\m100.u0/ethc0/r_reg[txlength_n_0_][7] ),
        .I5(\m100.u0/ethc0/r_reg[txlength_n_0_][8] ),
        .O(\r[tmsto][write]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT4 #(
    .INIT(16'h15EA)) 
    \r[tpnt][0]_i_1 
       (.I0(\r[abufs][2]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/rin[status][txahberr] ),
        .I2(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I3(\m100.u0/eraddress [7]),
        .O(\r[tpnt][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT5 #(
    .INIT(32'h557FAA80)) 
    \r[tpnt][1]_i_1 
       (.I0(\m100.u0/eraddress [7]),
        .I1(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I2(\m100.u0/ethc0/rin[status][txahberr] ),
        .I3(\r[abufs][2]_i_6_n_0 ),
        .I4(\m100.u0/eraddress [8]),
        .O(\r[tpnt][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r[tpnt][1]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\m100.u0/ethc0/rin[status][txahberr] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][10]_i_1 
       (.I0(\m100.u0/erdata [10]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [10]),
        .O(\r[txaddr][10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][11]_i_1 
       (.I0(\m100.u0/erdata [11]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [11]),
        .O(\r[txaddr][11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][12]_i_1 
       (.I0(\m100.u0/erdata [12]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [12]),
        .O(\r[txaddr][12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][13]_i_1 
       (.I0(\m100.u0/erdata [13]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [13]),
        .O(\r[txaddr][13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][14]_i_1 
       (.I0(\m100.u0/erdata [14]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [14]),
        .O(\r[txaddr][14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][15]_i_1 
       (.I0(\m100.u0/erdata [15]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [15]),
        .O(\r[txaddr][15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][16]_i_1 
       (.I0(\m100.u0/erdata [16]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [16]),
        .O(\r[txaddr][16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][17]_i_1 
       (.I0(\m100.u0/erdata [17]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [17]),
        .O(\r[txaddr][17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][18]_i_1 
       (.I0(\m100.u0/erdata [18]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [18]),
        .O(\r[txaddr][18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][19]_i_1 
       (.I0(\m100.u0/erdata [19]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [19]),
        .O(\r[txaddr][19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][20]_i_1 
       (.I0(\m100.u0/erdata [20]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [20]),
        .O(\r[txaddr][20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][21]_i_1 
       (.I0(\m100.u0/erdata [21]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [21]),
        .O(\r[txaddr][21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][22]_i_1 
       (.I0(\m100.u0/erdata [22]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [22]),
        .O(\r[txaddr][22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][23]_i_1 
       (.I0(\m100.u0/erdata [23]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [23]),
        .O(\r[txaddr][23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][24]_i_1 
       (.I0(\m100.u0/erdata [24]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [24]),
        .O(\r[txaddr][24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][25]_i_1 
       (.I0(\m100.u0/erdata [25]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [25]),
        .O(\r[txaddr][25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][26]_i_1 
       (.I0(\m100.u0/erdata [26]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [26]),
        .O(\r[txaddr][26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][27]_i_1 
       (.I0(\m100.u0/erdata [27]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [27]),
        .O(\r[txaddr][27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][28]_i_1 
       (.I0(\m100.u0/erdata [28]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [28]),
        .O(\r[txaddr][28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][29]_i_1 
       (.I0(\m100.u0/erdata [29]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [29]),
        .O(\r[txaddr][29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][2]_i_1 
       (.I0(\m100.u0/erdata [2]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [2]),
        .O(\r[txaddr][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][30]_i_1 
       (.I0(\m100.u0/erdata [30]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [30]),
        .O(\r[txaddr][30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF2000)) 
    \r[txaddr][31]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/tmsti[ready] ),
        .I3(\r[txstatus][1]_i_2_n_0 ),
        .I4(\r[txaddr][31]_i_4_n_0 ),
        .O(\r[txaddr][31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][31]_i_2 
       (.I0(\m100.u0/erdata [31]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [31]),
        .O(\r[txaddr][31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h04000000)) 
    \r[txaddr][31]_i_3 
       (.I0(\ahbmi[hresp] [0]),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\ahbmi[hresp] [1]),
        .I3(\ahbmi[hready] ),
        .I4(\m100.u0/ethc0/ahb0/r_reg ),
        .O(\m100.u0/ethc0/tmsti[ready] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00100000)) 
    \r[txaddr][31]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I3(\r[txdstate][2]_i_5_n_0 ),
        .I4(\r[txlength][10]_i_10_n_0 ),
        .O(\r[txaddr][31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][3]_i_1 
       (.I0(\m100.u0/erdata [3]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [3]),
        .O(\r[txaddr][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][4]_i_1 
       (.I0(\m100.u0/erdata [4]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [4]),
        .O(\r[txaddr][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][5]_i_1 
       (.I0(\m100.u0/erdata [5]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [5]),
        .O(\r[txaddr][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][6]_i_1 
       (.I0(\m100.u0/erdata [6]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [6]),
        .O(\r[txaddr][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][7]_i_1 
       (.I0(\m100.u0/erdata [7]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [7]),
        .O(\r[txaddr][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][8]_i_1 
       (.I0(\m100.u0/erdata [8]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [8]),
        .O(\r[txaddr][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[txaddr][9]_i_1 
       (.I0(\m100.u0/erdata [9]),
        .I1(\r[txaddr][31]_i_4_n_0 ),
        .I2(\ahbmi[hrdata] [9]),
        .O(\r[txaddr][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000D5FF)) 
    \r[txburstav]_i_1 
       (.I0(\r[txdstate][0]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\r[txburstav]_i_2_n_0 ),
        .O(\r[txburstav]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02FF0200)) 
    \r[txburstav]_i_2 
       (.I0(\r[txdataav]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[tfcnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[tfcnt_n_0_][6] ),
        .I3(\m100.u0/ethc0/r_reg[tfcnt_n_0_][7] ),
        .I4(\r[txburstav]_i_3_n_0 ),
        .O(\r[txburstav]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \r[txburstav]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[tfcnt_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[tfcnt_n_0_][6] ),
        .I2(\m100.u0/ethc0/r_reg[tfcnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[tfcnt_n_0_][4] ),
        .I4(\m100.u0/ethc0/r_reg[tfcnt_n_0_][5] ),
        .I5(\r[txburstav]_i_4_n_0 ),
        .O(\r[txburstav]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \r[txburstav]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[tfcnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[tfcnt_n_0_][0] ),
        .O(\r[txburstav]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FFFFAFAE0000)) 
    \r[txburstcnt][0]_i_1 
       (.I0(\m100.u0/ethc0/tmsti[retry] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\r[txburstcnt][1]_i_5_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txburstcnt_n_0_][0] ),
        .O(\r[txburstcnt][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9998FFFF66640000)) 
    \r[txburstcnt][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txburstcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/tmsti[retry] ),
        .I2(\r[txburstcnt][1]_i_3_n_0 ),
        .I3(\r[txburstcnt][1]_i_4_n_0 ),
        .I4(\r[txburstcnt][1]_i_5_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txburstcnt_n_0_][1] ),
        .O(\r[txburstcnt][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \r[txburstcnt][1]_i_2 
       (.I0(\ahbmi[hresp] [1]),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\m100.u0/ethc0/ahb0/r_reg ),
        .I3(\ahbmi[hready] ),
        .O(\m100.u0/ethc0/tmsti[retry] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[txburstcnt][1]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txburstcnt][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[txburstcnt][1]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txburstcnt][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAABBBABBFB)) 
    \r[txburstcnt][1]_i_5 
       (.I0(\m100.u0/ethc0/tmsti[retry] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/tmsti ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[txburstcnt][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFE0FFE0FFFFFFE0)) 
    \r[txcnt][0]_i_1 
       (.I0(\r[tcnt][4]_i_5_n_0 ),
        .I1(\r[txcnt][7]_i_5_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I3(\r[txcnt][0]_i_2_n_0 ),
        .I4(\m100.u0/erdata [0]),
        .I5(\r[txlength][10]_i_5_n_0 ),
        .O(\r[txcnt][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000F040400000404)) 
    \r[txcnt][0]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[txlength_n_0_][0] ),
        .O(\r[txcnt][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFF01FFFF)) 
    \r[txcnt][10]_i_1 
       (.I0(\r[txcnt][10]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\r[txcnt][10]_i_4_n_0 ),
        .I3(\r[tcnt][4]_i_5_n_0 ),
        .I4(\r[txlength][10]_i_5_n_0 ),
        .I5(\r[txcnt][10]_i_5_n_0 ),
        .O(\r[txcnt][10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF1F1F11F11111111)) 
    \r[txcnt][10]_i_2 
       (.I0(\r[txcnt][10]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][10] ),
        .I3(\r[txcnt][10]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][9] ),
        .I5(\r[tcnt][4]_i_5_n_0 ),
        .O(\r[txcnt][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r[txcnt][10]_i_3 
       (.I0(\r_reg[tmsto][write]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txden]__0 ),
        .O(\r[txcnt][10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r[txcnt][10]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[txcnt][10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0005010500010101)) 
    \r[txcnt][10]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\a9.x[0].r0_i_34__1_n_0 ),
        .I5(\m100.u0/ethc0/tmsti[ready] ),
        .O(\r[txcnt][10]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFF4BFF)) 
    \r[txcnt][10]_i_6 
       (.I0(\r[txcnt][9]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][9] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][10] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\r[txcnt][10]_i_8_n_0 ),
        .O(\r[txcnt][10]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r[txcnt][10]_i_7 
       (.I0(\r[txcnt][10]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][6] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][8] ),
        .I5(\m100.u0/ethc0/r_reg[txcnt_n_0_][7] ),
        .O(\r[txcnt][10]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E0FF0000E00000)) 
    \r[txcnt][10]_i_8 
       (.I0(\r[txcnt][10]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][9] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][10] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[txlength_n_0_][10] ),
        .O(\r[txcnt][10]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r[txcnt][10]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .O(\r[txcnt][10]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFF0C0D0C)) 
    \r[txcnt][1]_i_1 
       (.I0(\r[txcnt][6]_i_4_n_0 ),
        .I1(\r[txcnt][1]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .I4(\r[tcnt][4]_i_5_n_0 ),
        .I5(\r[txcnt][1]_i_3_n_0 ),
        .O(\r[txcnt][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0028FF2800280028)) 
    \r[txcnt][1]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[txlength_n_0_][1] ),
        .O(\r[txcnt][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \r[txcnt][1]_i_3 
       (.I0(\r[txlength][7]_i_4_n_0 ),
        .I1(\m100.u0/erdata [1]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r[txcnt][5]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I5(\r[txcnt][1]_i_4_n_0 ),
        .O(\r[txcnt][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    \r[txcnt][1]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][4] ),
        .I4(\m100.u0/ethc0/r_reg[tcnt_n_0_][5] ),
        .I5(\m100.u0/ethc0/r_reg[tcnt_n_0_][6] ),
        .O(\r[txcnt][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h22FF22222F2F2F2F)) 
    \r[txcnt][2]_i_1 
       (.I0(\r[txcnt][7]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I2(\r[txcnt][2]_i_2_n_0 ),
        .I3(\r[txcnt][2]_i_3_n_0 ),
        .I4(\r[txcnt][5]_i_4_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[txcnt][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB0BFBFB0BFBFBFBF)) 
    \r[txcnt][2]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r[txcnt][7]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\r[txcnt][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0EEEEEEE)) 
    \r[txcnt][2]_i_3 
       (.I0(\r[tcnt][4]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/erdata [2]),
        .I4(\r[txlength][10]_i_12_n_0 ),
        .O(\r[txcnt][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h03005555)) 
    \r[txcnt][3]_i_1 
       (.I0(\r[txcnt][3]_i_2_n_0 ),
        .I1(\r[txcnt][3]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[txcnt][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F6F6F6)) 
    \r[txcnt][3]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I2(\r[txcnt][6]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txlength_n_0_][3] ),
        .I4(\r[txcnt][6]_i_5_n_0 ),
        .I5(\r[txcnt][3]_i_4_n_0 ),
        .O(\r[txcnt][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00F6F6F6F6F6F6F6)) 
    \r[txcnt][3]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I2(\r[tcnt][4]_i_9_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/erdata [3]),
        .I5(\r[txlength][10]_i_12_n_0 ),
        .O(\r[txcnt][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000078F00000)) 
    \r[txcnt][3]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txcnt][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF0000F1F1F1F1)) 
    \r[txcnt][4]_i_1 
       (.I0(\r[txcnt][4]_i_2_n_0 ),
        .I1(\r[txcnt][6]_i_4_n_0 ),
        .I2(\r[txcnt][4]_i_3_n_0 ),
        .I3(\r[txcnt][4]_i_4_n_0 ),
        .I4(\r[txcnt][5]_i_4_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[txcnt][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h56)) 
    \r[txcnt][4]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .O(\r[txcnt][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F20202020202F20)) 
    \r[txcnt][4]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\r[txcnt][9]_i_4_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .O(\r[txcnt][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00F6F6F6F6F6F6F6)) 
    \r[txcnt][4]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .I1(\r[txcnt][10]_i_9_n_0 ),
        .I2(\r[tcnt][4]_i_9_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/erdata [4]),
        .I5(\r[txlength][10]_i_12_n_0 ),
        .O(\r[txcnt][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0C5D0C5DFF5D0C5D)) 
    \r[txcnt][5]_i_1 
       (.I0(\r[txcnt][5]_i_2_n_0 ),
        .I1(\r[txcnt][7]_i_5_n_0 ),
        .I2(\r[txcnt][5]_i_3_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r[txcnt][5]_i_4_n_0 ),
        .I5(\r[txcnt][5]_i_5_n_0 ),
        .O(\r[txcnt][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB0BFBFB0BFBFBFBF)) 
    \r[txcnt][5]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\r[txcnt][5]_i_6_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\r[txcnt][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5556)) 
    \r[txcnt][5]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .O(\r[txcnt][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[txcnt][5]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[txcnt][5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0EEEEEEE)) 
    \r[txcnt][5]_i_5 
       (.I0(\r[txcnt][5]_i_3_n_0 ),
        .I1(\r[tcnt][4]_i_9_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/erdata [5]),
        .I4(\r[txlength][10]_i_12_n_0 ),
        .O(\r[txcnt][5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \r[txcnt][5]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .O(\r[txcnt][5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFAFAAABAAABAAAB)) 
    \r[txcnt][6]_i_1 
       (.I0(\r[txcnt][6]_i_2_n_0 ),
        .I1(\r[txcnt][6]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[txcnt][6]_i_4_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txlength_n_0_][6] ),
        .I5(\r[txcnt][6]_i_5_n_0 ),
        .O(\r[txcnt][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h888A88888888888A)) 
    \r[txcnt][6]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\r[txcnt][6]_i_6_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\r[txcnt][6]_i_7_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txcnt_n_0_][6] ),
        .O(\r[txcnt][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55555556)) 
    \r[txcnt][6]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][6] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .O(\r[txcnt][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBBBFB)) 
    \r[txcnt][6]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\r[txcnt][6]_i_8_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .O(\r[txcnt][6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[txcnt][6]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[txcnt][6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8080000080FF0000)) 
    \r[txcnt][6]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/erdata [6]),
        .I2(\r[txlength][10]_i_12_n_0 ),
        .I3(\r[tcnt][4]_i_9_n_0 ),
        .I4(\r[txdstate][0]_i_2_n_0 ),
        .I5(\r[txcnt][6]_i_3_n_0 ),
        .O(\r[txcnt][6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \r[txcnt][6]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .O(\r[txcnt][6]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \r[txcnt][6]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][10] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][9] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][7] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][8] ),
        .I4(\r[txcnt][6]_i_9_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txcnt_n_0_][6] ),
        .O(\r[txcnt][6]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r[txcnt][6]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .O(\r[txcnt][6]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF4F4F4F1F1FFF1)) 
    \r[txcnt][7]_i_1 
       (.I0(\r[txcnt][7]_i_2_n_0 ),
        .I1(\r[txcnt][7]_i_3_n_0 ),
        .I2(\r[txcnt][7]_i_4_n_0 ),
        .I3(\r[txcnt][7]_i_5_n_0 ),
        .I4(\r[txcnt][7]_i_6_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txcnt_n_0_][7] ),
        .O(\r[txcnt][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \r[txcnt][7]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\r[txcnt][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF7FFFFFFFFFFFFF)) 
    \r[txcnt][7]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I3(\r[txcnt][7]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .I5(\m100.u0/ethc0/r_reg[txcnt_n_0_][6] ),
        .O(\r[txcnt][7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \r[txcnt][7]_i_4 
       (.I0(\r[txlength][10]_i_5_n_0 ),
        .I1(\m100.u0/erdata [7]),
        .I2(\r[tcnt][4]_i_5_n_0 ),
        .I3(\r[txcnt][7]_i_8_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txlength_n_0_][7] ),
        .I5(\r[txcnt][9]_i_5_n_0 ),
        .O(\r[txcnt][7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[txcnt][7]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\r[txcnt][6]_i_4_n_0 ),
        .O(\r[txcnt][7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \r[txcnt][7]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][6] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .O(\r[txcnt][7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \r[txcnt][7]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .O(\r[txcnt][7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555555555555556)) 
    \r[txcnt][7]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][6] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .I5(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .O(\r[txcnt][7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF02000002)) 
    \r[txcnt][8]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][8] ),
        .I4(\r[txcnt][8]_i_2_n_0 ),
        .I5(\r[txcnt][8]_i_3_n_0 ),
        .O(\r[txcnt][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF7FFFFFF)) 
    \r[txcnt][8]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][6] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .I2(\r[txcnt][9]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][7] ),
        .O(\r[txcnt][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFECCCCCCCCFE)) 
    \r[txcnt][8]_i_3 
       (.I0(\r[tcnt][4]_i_5_n_0 ),
        .I1(\r[txcnt][8]_i_4_n_0 ),
        .I2(\r[txcnt][7]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][7] ),
        .I4(\r[txcnt][7]_i_6_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txcnt_n_0_][8] ),
        .O(\r[txcnt][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h808F808080808080)) 
    \r[txcnt][8]_i_4 
       (.I0(\m100.u0/erdata [8]),
        .I1(\r[txlength][10]_i_6_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[txlength_n_0_][8] ),
        .O(\r[txcnt][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF02000002)) 
    \r[txcnt][9]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][9] ),
        .I4(\r[txcnt][9]_i_2_n_0 ),
        .I5(\r[txcnt][9]_i_3_n_0 ),
        .O(\r[txcnt][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF7FFFFFFFFFFFFFF)) 
    \r[txcnt][9]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .I2(\r[txcnt][9]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][6] ),
        .I5(\m100.u0/ethc0/r_reg[txcnt_n_0_][8] ),
        .O(\r[txcnt][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF30FF30FFFFFFBA)) 
    \r[txcnt][9]_i_3 
       (.I0(\r[txcnt][7]_i_5_n_0 ),
        .I1(\r[txcnt][9]_i_5_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][9] ),
        .I3(\r[txcnt][9]_i_6_n_0 ),
        .I4(\r[tcnt][4]_i_5_n_0 ),
        .I5(\r[txcnt][9]_i_7_n_0 ),
        .O(\r[txcnt][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \r[txcnt][9]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .O(\r[txcnt][9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \r[txcnt][9]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txcnt][9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    \r[txcnt][9]_i_6 
       (.I0(\r[txlength][10]_i_12_n_0 ),
        .I1(\m100.u0/erdata [9]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txcnt][9]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5556)) 
    \r[txcnt][9]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][9] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][7] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][8] ),
        .I3(\r[txcnt][7]_i_6_n_0 ),
        .O(\r[txcnt][9]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[txdata][31]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txread] ),
        .I1(\m100.u0/ethc0/r_reg[txreadack]__0 ),
        .O(\m100.u0/ethc0/v[tfrpnt]1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFFFFFFFEFEFEFEF)) 
    \r[txdataav]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[tfcnt_n_0_][7] ),
        .I1(\m100.u0/ethc0/r_reg[tfcnt_n_0_][6] ),
        .I2(\r[txdataav]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdataav_n_0_] ),
        .I4(\m100.u0/ethc0/v[tfrpnt]1 ),
        .I5(\m100.u0/ethc0/r_reg[tfcnt_n_0_][0] ),
        .O(\m100.u0/txrenable ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \r[txdataav]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[tfcnt_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[tfcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[tfcnt_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[tfcnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[tfcnt_n_0_][3] ),
        .O(\r[txdataav]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \r[txdesc][31]_i_1 
       (.I0(\apbo[prdata][14]_INST_0_i_5_n_0 ),
        .I1(\apbi[pwrite] ),
        .I2(apbi[15]),
        .I3(\apbi[penable] ),
        .I4(\apbi[paddr] [2]),
        .I5(\apbi[paddr] [3]),
        .O(\m100.u0/ethc0/v[txdsel] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r[txdone][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I1(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I2(\r[txdone][1]_i_2_n_0 ),
        .O(\r[txdone][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF0FFDFFFFF0FFF)) 
    \r[txdone][1]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txstart]__0 ),
        .I1(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[txdone][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1F10)) 
    \r[txdsel][3]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txwrap_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[txdsel_n_0_][3] ),
        .I2(\r[txdsel][9]_i_3_n_0 ),
        .I3(\apbi[pwdata] [3]),
        .O(\r[txdsel][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h06FF0600)) 
    \r[txdsel][4]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdsel_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[txdsel_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txwrap_n_0_] ),
        .I3(\r[txdsel][9]_i_3_n_0 ),
        .I4(\apbi[pwdata] [4]),
        .O(\r[txdsel][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1540FFFF15400000)) 
    \r[txdsel][5]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txwrap_n_0_] ),
        .I1(\m100.u0/ethc0/r_reg[txdsel_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdsel_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[txdsel_n_0_][5] ),
        .I4(\r[txdsel][9]_i_3_n_0 ),
        .I5(\apbi[pwdata] [5]),
        .O(\r[txdsel][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h14FF1400)) 
    \r[txdsel][6]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txwrap_n_0_] ),
        .I1(\r[txdsel][6]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdsel_n_0_][6] ),
        .I3(\r[txdsel][9]_i_3_n_0 ),
        .I4(\apbi[pwdata] [6]),
        .O(\r[txdsel][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \r[txdsel][6]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdsel_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[txdsel_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdsel_n_0_][5] ),
        .O(\r[txdsel][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h14FF1400)) 
    \r[txdsel][7]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txwrap_n_0_] ),
        .I1(\r[txdsel][7]_i_2_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdsel_n_0_][7] ),
        .I3(\r[txdsel][9]_i_3_n_0 ),
        .I4(\apbi[pwdata] [7]),
        .O(\r[txdsel][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \r[txdsel][7]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdsel_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[txdsel_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdsel_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[txdsel_n_0_][6] ),
        .O(\r[txdsel][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h14FF1400)) 
    \r[txdsel][8]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txwrap_n_0_] ),
        .I1(\r[txdsel][9]_i_4_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdsel_n_0_][8] ),
        .I3(\r[txdsel][9]_i_3_n_0 ),
        .I4(\apbi[pwdata] [8]),
        .O(\r[txdsel][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r[txdsel][9]_i_1 
       (.I0(\m100.u0/ethc0/v[txdsel] ),
        .I1(\r[txdsel][9]_i_3_n_0 ),
        .O(\r[txdsel][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0078FFFF00780000)) 
    \r[txdsel][9]_i_2 
       (.I0(\r[txdsel][9]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdsel_n_0_][8] ),
        .I2(\m100.u0/ethc0/r_reg[txdsel_n_0_][9] ),
        .I3(\m100.u0/ethc0/r_reg[txwrap_n_0_] ),
        .I4(\r[txdsel][9]_i_3_n_0 ),
        .I5(\apbi[pwdata] [9]),
        .O(\r[txdsel][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00080000)) 
    \r[txdsel][9]_i_3 
       (.I0(\m100.u0/ethc0/tmsti[ready] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txdsel][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \r[txdsel][9]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txdsel_n_0_][6] ),
        .I1(\m100.u0/ethc0/r_reg[txdsel_n_0_][4] ),
        .I2(\m100.u0/ethc0/r_reg[txdsel_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdsel_n_0_][5] ),
        .I4(\m100.u0/ethc0/r_reg[txdsel_n_0_][7] ),
        .O(\r[txdsel][9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEEE22E2)) 
    \r[txdstate][0]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\r[txdstate][3]_i_5_n_0 ),
        .I2(\r[txdstate][0]_i_2_n_0 ),
        .I3(\r[txdstate][0]_i_3_n_0 ),
        .I4(\r[txdstate][0]_i_4_n_0 ),
        .I5(\m100.u0/ethc0/rin[tmsto][req] ),
        .O(\r[txdstate][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[txdstate][0]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[txdstate][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FFFFFFFFFDFD)) 
    \r[txdstate][0]_i_3 
       (.I0(\r[tedcl]_i_2_n_0 ),
        .I1(\r[tfwpnt][6]_i_5_n_0 ),
        .I2(\r[tfwpnt][6]_i_4_n_0 ),
        .I3(\r[txdstate][2]_i_2_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\r[txdstate][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0101010101054145)) 
    \r[txdstate][0]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\r[txcnt][10]_i_3_n_0 ),
        .I4(\r[txdstate][0]_i_5_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[txdstate][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF6F6F6F6FFF6FFFF)) 
    \r[txdstate][0]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .I1(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I3(\r[txdstate][0]_i_6_n_0 ),
        .I4(\r[txdstate][0]_i_7_n_0 ),
        .I5(\r[tfwpnt][6]_i_5_n_0 ),
        .O(\r[txdstate][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF4FFF4FFFFFFF4)) 
    \r[txdstate][0]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][8] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][6] ),
        .I5(\m100.u0/ethc0/r_reg[txcnt_n_0_][7] ),
        .O(\r[txdstate][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \r[txdstate][0]_i_7 
       (.I0(\r[txdstate][0]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][4] ),
        .I5(\m100.u0/ethc0/r_reg[txcnt_n_0_][5] ),
        .O(\r[txdstate][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \r[txdstate][0]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][8] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][7] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][9] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][10] ),
        .O(\r[txdstate][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000002E2E2E22)) 
    \r[txdstate][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\r[txdstate][3]_i_5_n_0 ),
        .I2(\r[txdstate][1]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r[txdstate][1]_i_3_n_0 ),
        .I5(\m100.u0/ethc0/rin[tmsto][req] ),
        .O(\r[txdstate][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000099000000000F)) 
    \r[txdstate][1]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I1(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I2(\m100.u0/ethc0/v[tmsto][req]1149_out ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[txdstate][1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h10F010F0FFFF10F0)) 
    \r[txdstate][1]_i_2 
       (.I0(\r[txdstate][1]_i_5_n_0 ),
        .I1(\r[txdstate][1]_i_6_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\r[txdstate][1]_i_7_n_0 ),
        .I4(\r[txdstate][1]_i_8_n_0 ),
        .I5(\r[txdstate][1]_i_9_n_0 ),
        .O(\r[txdstate][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFFF4F)) 
    \r[txdstate][1]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txden]__0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\r[txdstate][3]_i_10_n_0 ),
        .I5(\r[txdstate][1]_i_10_n_0 ),
        .O(\r[txdstate][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \r[txdstate][1]_i_4 
       (.I0(\m100.u0/ethc0/v[tmsto][req]0139_out ),
        .I1(\m100.u0/ethc0/p_6_in [6]),
        .I2(rst),
        .O(\m100.u0/ethc0/rin[tmsto][req] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFBEFFFFFFFF)) 
    \r[txdstate][1]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .I3(\r[tfwpnt][6]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\r[tedcl]_i_2_n_0 ),
        .O(\r[txdstate][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \r[txdstate][1]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[write_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[write_n_0_][2] ),
        .I2(\m100.u0/eraddress [8]),
        .I3(\m100.u0/ethc0/r_reg[write_n_0_][1] ),
        .I4(\m100.u0/eraddress [7]),
        .I5(\m100.u0/ethc0/r_reg[write_n_0_][0] ),
        .O(\r[txdstate][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F00010F010F)) 
    \r[txdstate][1]_i_7 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I1(\r[tmsto][data][31]_i_6_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\r[txdstate][2]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txdstate][1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[txdstate][1]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txdstate][1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h28AAAA28)) 
    \r[txdstate][1]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I4(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .O(\r[txdstate][1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF1FFFFFFF100)) 
    \r[txdstate][2]_i_1 
       (.I0(\r[txdstate][2]_i_2_n_0 ),
        .I1(\r[txdstate][2]_i_3_n_0 ),
        .I2(\r[txdstate][2]_i_4_n_0 ),
        .I3(\r[txdstate][3]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/v[tmsto][req]0139_out ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[txdstate][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFBFF)) 
    \r[txdstate][2]_i_2 
       (.I0(\r[txdstate][2]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .O(\r[txdstate][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBFFF)) 
    \r[txdstate][2]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txdstate][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040000011401100)) 
    \r[txdstate][2]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\r[tfwpnt][6]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\r[txdstate][2]_i_6_n_0 ),
        .O(\r[txdstate][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFEFF)) 
    \r[txdstate][2]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][6] ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][5] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][4] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][3] ),
        .O(\r[txdstate][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE0EEEFEEEFEEEFEE)) 
    \r[txdstate][2]_i_6 
       (.I0(\r[tfwpnt][6]_i_4_n_0 ),
        .I1(\r[txdstate][3]_i_15_n_0 ),
        .I2(\r[txcnt][5]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txden]__0 ),
        .I5(\r_reg[tmsto][write]_i_2_n_0 ),
        .O(\r[txdstate][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF2FFFFFFF200)) 
    \r[txdstate][3]_i_1 
       (.I0(\r[txdstate][3]_i_2_n_0 ),
        .I1(\r[txdstate][3]_i_3_n_0 ),
        .I2(\r[txdstate][3]_i_4_n_0 ),
        .I3(\r[txdstate][3]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/v[tmsto][req]0139_out ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[txdstate][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h20AA0000000020AA)) 
    \r[txdstate][3]_i_10 
       (.I0(\r[txdstate][3]_i_15_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .I5(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .O(\r[txdstate][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h41FF41FF41FF4100)) 
    \r[txdstate][3]_i_11 
       (.I0(\r[tfwpnt][6]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .I2(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I5(\a9.x[0].r0_i_34__1_n_0 ),
        .O(\r[txdstate][3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4FFF4F0F4FFF4FF)) 
    \r[txdstate][3]_i_12 
       (.I0(\r[txdstate][3]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\r[txdstate][3]_i_16_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\r[txdstate][3]_i_17_n_0 ),
        .I5(\r[txstart_sync]_i_3_n_0 ),
        .O(\r[txdstate][3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FF1D001D)) 
    \r[txdstate][3]_i_13 
       (.I0(\m100.u0/ethc0/p_6_in [0]),
        .I1(\m100.u0/ethc0/v[tmsto][req]1149_out ),
        .I2(\m100.u0/erenable ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\r[txdstate][3]_i_18_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txdstate][3]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0808080808880808)) 
    \r[txdstate][3]_i_14 
       (.I0(\r[txdstate][3]_i_19_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\r[txdstate][3]_i_20_n_0 ),
        .I3(\r[tfwpnt][6]_i_5_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txstart]__0 ),
        .I5(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .O(\r[txdstate][3]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6F006600)) 
    \r[txdstate][3]_i_15 
       (.I0(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I1(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I2(\r[txdstate][0]_i_6_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I4(\r[txdstate][0]_i_7_n_0 ),
        .O(\r[txdstate][3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h08FF)) 
    \r[txdstate][3]_i_16 
       (.I0(\m100.u0/ethc0/tmsti[ready] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txdstate][3]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFEFFFF)) 
    \r[txdstate][3]_i_17 
       (.I0(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I1(\m100.u0/ethc0/r_reg[txburstav]__0 ),
        .I2(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\r[tfwpnt][6]_i_5_n_0 ),
        .O(\r[txdstate][3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \r[txdstate][3]_i_18 
       (.I0(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/tmsti[ready] ),
        .O(\r[txdstate][3]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hECFCECCCEFFCEFCC)) 
    \r[txdstate][3]_i_19 
       (.I0(\r[txdstate][2]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\r[txstart_sync]_i_5_n_0 ),
        .I5(\r[txdstate][3]_i_21_n_0 ),
        .O(\r[txdstate][3]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8F)) 
    \r[txdstate][3]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[txdstate][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \r[txdstate][3]_i_20 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txdstate][3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h04000000)) 
    \r[txdstate][3]_i_21 
       (.I0(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .I1(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I2(\ahbmi[hresp] [1]),
        .I3(\ahbmi[hready] ),
        .I4(\m100.u0/ethc0/ahb0/r_reg ),
        .O(\r[txdstate][3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBFFFB0FFBFFFBFF)) 
    \r[txdstate][3]_i_3 
       (.I0(\r[txdstate][3]_i_7_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\r[txdstate][3]_i_8_n_0 ),
        .I5(\r[txdstate][3]_i_9_n_0 ),
        .O(\r[txdstate][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABAAAAAA)) 
    \r[txdstate][3]_i_4 
       (.I0(\r[tcnt][6]_i_4_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\r[txdstate][3]_i_10_n_0 ),
        .O(\r[txdstate][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000BABABFBA)) 
    \r[txdstate][3]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\r[txdstate][3]_i_11_n_0 ),
        .I2(\r[txburstcnt][1]_i_4_n_0 ),
        .I3(\r[txdstate][3]_i_12_n_0 ),
        .I4(\r[txdstate][3]_i_13_n_0 ),
        .I5(\r[txdstate][3]_i_14_n_0 ),
        .O(\r[txdstate][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000008000000)) 
    \r[txdstate][3]_i_6 
       (.I0(\m100.u0/ethc0/ahb0/r_reg ),
        .I1(\ahbmi[hready] ),
        .I2(\ahbmi[hresp] [1]),
        .I3(\m100.u0/ethc0/ahb0/r_reg[bo]__0 ),
        .I4(\ahbmi[hresp] [0]),
        .I5(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .O(\m100.u0/ethc0/v[tmsto][req]0139_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAA2AAAAA8AA)) 
    \r[txdstate][3]_i_7 
       (.I0(\r[txstart_sync]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I4(\r[txdstate][2]_i_5_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[tarp]__0 ),
        .O(\r[txdstate][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA8)) 
    \r[txdstate][3]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\r[tmsto][data][31]_i_6_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .O(\r[txdstate][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF6FFFFFFFFFFFF)) 
    \r[txdstate][3]_i_9 
       (.I0(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .I1(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .I2(\r[tfwpnt][6]_i_5_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\r[tedcl]_i_2_n_0 ),
        .I5(\r[txdstate][1]_i_6_n_0 ),
        .O(\r[txdstate][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000002F22FFFF)) 
    \r[txlength][0]_i_1 
       (.I0(\m100.u0/erdata [0]),
        .I1(\r[txlength][6]_i_2_n_0 ),
        .I2(\r[txlength][8]_i_2_n_0 ),
        .I3(\ahbmi[hrdata] [0]),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I5(\r[txlength][0]_i_2_n_0 ),
        .O(\r[txlength][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00007707)) 
    \r[txlength][0]_i_2 
       (.I0(\r[txlength][10]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][0] ),
        .I2(\ahbmi[hrdata] [0]),
        .I3(\r[txlength][10]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[txlength][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \r[txlength][10]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[tarp]0 ),
        .I1(\m100.u0/ethc0/v[txirq] ),
        .I2(\r[txlength][10]_i_5_n_0 ),
        .O(\r[txlength][10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4000)) 
    \r[txlength][10]_i_10 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[txlength][10]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \r[txlength][10]_i_11 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .O(\r[txlength][10]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0100)) 
    \r[txlength][10]_i_12 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I1(\r[txdstate][2]_i_5_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .O(\r[txlength][10]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFBFFFF)) 
    \r[txlength][10]_i_13 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][6] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\r[txlength][10]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0015FFFF)) 
    \r[txlength][10]_i_14 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txlength_n_0_][5] ),
        .I4(\m100.u0/ethc0/r_reg[txlength_n_0_][6] ),
        .O(\r[txlength][10]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    \r[txlength][10]_i_15 
       (.I0(\m100.u0/erdata [16]),
        .I1(\m100.u0/erdata [18]),
        .I2(\m100.u0/erdata [26]),
        .I3(\m100.u0/erdata [19]),
        .I4(\r[txlength][10]_i_17_n_0 ),
        .O(\r[txlength][10]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \r[txlength][10]_i_16 
       (.I0(\m100.u0/erdata [28]),
        .I1(\m100.u0/erdata [30]),
        .I2(\m100.u0/erdata [29]),
        .I3(\m100.u0/erdata [31]),
        .I4(\m100.u0/erdata [25]),
        .O(\r[txlength][10]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r[txlength][10]_i_17 
       (.I0(\m100.u0/erdata [21]),
        .I1(\m100.u0/erdata [20]),
        .I2(\m100.u0/erdata [23]),
        .I3(\m100.u0/erdata [22]),
        .O(\r[txlength][10]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4700773347004700)) 
    \r[txlength][10]_i_2 
       (.I0(\r[txlength][10]_i_6_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\r[txlength][10]_i_7_n_0 ),
        .I3(\ahbmi[hrdata] [10]),
        .I4(\r[txlength][10]_i_8_n_0 ),
        .I5(\r[txlength][10]_i_9_n_0 ),
        .O(\r[txlength][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \r[txlength][10]_i_3 
       (.I0(\r[txlength][10]_i_10_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][6] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][5] ),
        .I4(\m100.u0/ethc0/r_reg[tcnt_n_0_][4] ),
        .I5(\r[txlength][10]_i_11_n_0 ),
        .O(\m100.u0/ethc0/r_reg[tarp]0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \r[txlength][10]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\r[txcnt][5]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .I5(\m100.u0/ethc0/tmsti[ready] ),
        .O(\m100.u0/ethc0/v[txirq] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF7FFFFF)) 
    \r[txlength][10]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I4(\r[txlength][10]_i_12_n_0 ),
        .O(\r[txlength][10]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \r[txlength][10]_i_6 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][5] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][3] ),
        .I4(\m100.u0/ethc0/r_reg[tcnt_n_0_][4] ),
        .I5(\r[txlength][10]_i_13_n_0 ),
        .O(\r[txlength][10]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \r[txlength][10]_i_7 
       (.I0(\r[txlength][10]_i_11_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][6] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][5] ),
        .I4(\m100.u0/ethc0/r_reg[tcnt_n_0_][4] ),
        .I5(\r[tfcnt][7]_i_3_n_0 ),
        .O(\r[txlength][10]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h59555555)) 
    \r[txlength][10]_i_8 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][10] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][9] ),
        .I2(\r[txlength][10]_i_14_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txlength_n_0_][8] ),
        .I4(\m100.u0/ethc0/r_reg[txlength_n_0_][7] ),
        .O(\r[txlength][10]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA8AAAAAAAAAAA)) 
    \r[txlength][10]_i_9 
       (.I0(\r[txlength][10]_i_7_n_0 ),
        .I1(\r[txlength][10]_i_15_n_0 ),
        .I2(\r[txlength][10]_i_16_n_0 ),
        .I3(\m100.u0/erdata [17]),
        .I4(\m100.u0/erdata [24]),
        .I5(\m100.u0/erdata [27]),
        .O(\r[txlength][10]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F44FFFF4F440000)) 
    \r[txlength][1]_i_1 
       (.I0(\r[txlength][8]_i_2_n_0 ),
        .I1(\ahbmi[hrdata] [1]),
        .I2(\r[txlength][6]_i_2_n_0 ),
        .I3(\m100.u0/erdata [1]),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I5(\r[txlength][1]_i_2_n_0 ),
        .O(\r[txlength][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hDDD0)) 
    \r[txlength][1]_i_2 
       (.I0(\r[txlength][10]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][1] ),
        .I2(\r[txlength][10]_i_7_n_0 ),
        .I3(\ahbmi[hrdata] [1]),
        .O(\r[txlength][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000002F22FFFF)) 
    \r[txlength][2]_i_1 
       (.I0(\m100.u0/erdata [2]),
        .I1(\r[txlength][6]_i_2_n_0 ),
        .I2(\r[txlength][8]_i_2_n_0 ),
        .I3(\ahbmi[hrdata] [2]),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I5(\r[txlength][2]_i_2_n_0 ),
        .O(\r[txlength][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000DD0D)) 
    \r[txlength][2]_i_2 
       (.I0(\r[txlength][10]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][2] ),
        .I2(\ahbmi[hrdata] [2]),
        .I3(\r[txlength][10]_i_7_n_0 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[txlength][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F44FFFF4F440000)) 
    \r[txlength][3]_i_1 
       (.I0(\r[txlength][8]_i_2_n_0 ),
        .I1(\ahbmi[hrdata] [3]),
        .I2(\r[txlength][6]_i_2_n_0 ),
        .I3(\m100.u0/erdata [3]),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I5(\r[txlength][3]_i_2_n_0 ),
        .O(\r[txlength][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7D7D7D00)) 
    \r[txlength][3]_i_2 
       (.I0(\r[txlength][10]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][3] ),
        .I3(\r[txlength][10]_i_7_n_0 ),
        .I4(\ahbmi[hrdata] [3]),
        .O(\r[txlength][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000002F22FFFF)) 
    \r[txlength][4]_i_1 
       (.I0(\m100.u0/erdata [4]),
        .I1(\r[txlength][6]_i_2_n_0 ),
        .I2(\r[txlength][8]_i_2_n_0 ),
        .I3(\ahbmi[hrdata] [4]),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I5(\r[txlength][4]_i_2_n_0 ),
        .O(\r[txlength][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000007D7D007D)) 
    \r[txlength][4]_i_2 
       (.I0(\r[txlength][10]_i_9_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][4] ),
        .I2(\r[txlength][4]_i_3_n_0 ),
        .I3(\ahbmi[hrdata] [4]),
        .I4(\r[txlength][10]_i_7_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[txlength][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[txlength][4]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][3] ),
        .O(\r[txlength][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F44FFFF4F440000)) 
    \r[txlength][5]_i_1 
       (.I0(\r[txlength][8]_i_2_n_0 ),
        .I1(\ahbmi[hrdata] [5]),
        .I2(\r[txlength][6]_i_2_n_0 ),
        .I3(\m100.u0/erdata [5]),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I5(\r[txlength][5]_i_2_n_0 ),
        .O(\r[txlength][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hE00EEEEE)) 
    \r[txlength][5]_i_2 
       (.I0(\r[txlength][10]_i_7_n_0 ),
        .I1(\ahbmi[hrdata] [5]),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][5] ),
        .I3(\r[txlength][5]_i_3_n_0 ),
        .I4(\r[txlength][10]_i_9_n_0 ),
        .O(\r[txlength][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \r[txlength][5]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][4] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][2] ),
        .O(\r[txlength][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000002F22FFFF)) 
    \r[txlength][6]_i_1 
       (.I0(\m100.u0/erdata [6]),
        .I1(\r[txlength][6]_i_2_n_0 ),
        .I2(\r[txlength][8]_i_2_n_0 ),
        .I3(\ahbmi[hrdata] [6]),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I5(\r[txlength][6]_i_3_n_0 ),
        .O(\r[txlength][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFEA)) 
    \r[txlength][6]_i_2 
       (.I0(\r[txlength][8]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .O(\r[txlength][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000006F6F006F)) 
    \r[txlength][6]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][6] ),
        .I1(\r[txlength][6]_i_4_n_0 ),
        .I2(\r[txlength][10]_i_9_n_0 ),
        .I3(\ahbmi[hrdata] [6]),
        .I4(\r[txlength][10]_i_7_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .O(\r[txlength][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0015)) 
    \r[txlength][6]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][5] ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txlength_n_0_][4] ),
        .O(\r[txlength][6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h90FF9090)) 
    \r[txlength][7]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txlength_n_0_][7] ),
        .I1(\r[txlength][10]_i_14_n_0 ),
        .I2(\r[txlength][10]_i_9_n_0 ),
        .I3(\r[txlength][10]_i_7_n_0 ),
        .I4(\ahbmi[hrdata] [7]),
        .O(\r[txlength][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4F444444)) 
    \r[txlength][7]_i_3 
       (.I0(\r[txlength][8]_i_2_n_0 ),
        .I1(\ahbmi[hrdata] [7]),
        .I2(\r[txlength][8]_i_5_n_0 ),
        .I3(\m100.u0/erdata [7]),
        .I4(\r[txlength][7]_i_4_n_0 ),
        .O(\r[txlength][7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h15)) 
    \r[txlength][7]_i_4 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .O(\r[txlength][7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDF0DDFFCCF0CCF0)) 
    \r[txlength][8]_i_1 
       (.I0(\r[txlength][8]_i_2_n_0 ),
        .I1(\r[txlength][8]_i_3_n_0 ),
        .I2(\r[txlength][8]_i_4_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I4(\r[txlength][10]_i_7_n_0 ),
        .I5(\ahbmi[hrdata] [8]),
        .O(\r[txlength][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0800)) 
    \r[txlength][8]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\r[txlength][10]_i_12_n_0 ),
        .O(\r[txlength][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00001500)) 
    \r[txlength][8]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I3(\m100.u0/erdata [8]),
        .I4(\r[txlength][8]_i_5_n_0 ),
        .O(\r[txlength][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h82A0)) 
    \r[txlength][8]_i_4 
       (.I0(\r[txlength][10]_i_9_n_0 ),
        .I1(\r[txlength][10]_i_14_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][8] ),
        .I3(\m100.u0/ethc0/r_reg[txlength_n_0_][7] ),
        .O(\r[txlength][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFDFFFFFF)) 
    \r[txlength][8]_i_5 
       (.I0(\r[txdstate][1]_i_6_n_0 ),
        .I1(\m100.u0/erdata [10]),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I5(\r[txcnt][1]_i_4_n_0 ),
        .O(\r[txlength][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF44F4444)) 
    \r[txlength][9]_i_2 
       (.I0(\r[txlength][10]_i_7_n_0 ),
        .I1(\ahbmi[hrdata] [9]),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][9] ),
        .I3(\r[txlength][9]_i_4_n_0 ),
        .I4(\r[txlength][10]_i_9_n_0 ),
        .O(\r[txlength][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8A8A8A8ABA8A8A8)) 
    \r[txlength][9]_i_3 
       (.I0(\ahbmi[hrdata] [9]),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][0] ),
        .I2(\r[txlength][9]_i_5_n_0 ),
        .I3(\m100.u0/erdata [9]),
        .I4(\r[txdstate][1]_i_6_n_0 ),
        .I5(\m100.u0/erdata [10]),
        .O(\r[txlength][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r[txlength][9]_i_4 
       (.I0(\r[txlength][10]_i_14_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txlength_n_0_][8] ),
        .I2(\m100.u0/ethc0/r_reg[txlength_n_0_][7] ),
        .O(\r[txlength][9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    \r[txlength][9]_i_5 
       (.I0(\r[txdstate][2]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[tcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[tcnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .O(\r[txlength][9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF0001FFFE0000)) 
    \r[txrestart][1]_i_1 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .I5(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .O(\r[txrestart][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3F3C3C3DFF3DFC3)) 
    \r[txstart]_i_2 
       (.I0(\r[tfwpnt][6]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I4(\r[txstart]_i_3_n_0 ),
        .I5(\r[tfwpnt][6]_i_4_n_0 ),
        .O(\r[txstart]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r[txstart]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[txstart]__0 ),
        .I1(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I2(\a9.x[0].r0_i_34__1_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[tmsto][req_n_0_] ),
        .O(\r[txstart]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \r[txstart_sync]_i_2 
       (.I0(\r[txstart_sync]_i_5_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[tedcl]__0 ),
        .I4(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I5(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .O(\r[txstart_sync]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFD)) 
    \r[txstart_sync]_i_3 
       (.I0(\r[txcnt][6]_i_8_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txcnt_n_0_][2] ),
        .I2(\m100.u0/ethc0/r_reg[txcnt_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txcnt_n_0_][0] ),
        .I4(\m100.u0/ethc0/r_reg[txcnt_n_0_][1] ),
        .O(\r[txstart_sync]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFE3E3E3)) 
    \r[txstart_sync]_i_4 
       (.I0(\r[txstart]_i_3_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I3(\r[tedcl]_i_2_n_0 ),
        .I4(\r[txdstate][1]_i_6_n_0 ),
        .O(\r[txstart_sync]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r[txstart_sync]_i_5 
       (.I0(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I1(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I2(\m100.u0/ethc0/r_reg[txrestart]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[txrestart]__0 [0]),
        .O(\r[txstart_sync]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45544004)) 
    \r[txstatus][0]_i_1 
       (.I0(\r[txstatus][1]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txstatus_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I4(\m100.u0/ethc0/txo[status] [0]),
        .O(\r[txstatus][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45544004)) 
    \r[txstatus][1]_i_1 
       (.I0(\r[txstatus][1]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/r_reg[txstatus_n_0_][1] ),
        .I2(\m100.u0/ethc0/r_reg[txdone]__0 [1]),
        .I3(\m100.u0/ethc0/r_reg[txdone]__0 [0]),
        .I4(\m100.u0/ethc0/txo[status] [1]),
        .O(\r[txstatus][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \r[txstatus][1]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[txdstate_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[txdstate_n_0_][0] ),
        .I2(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ),
        .I3(\m100.u0/ethc0/r_reg[txdstate_n_0_][1] ),
        .O(\r[txstatus][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \r[udpsrc][15]_i_1 
       (.I0(\r[udpsrc][15]_i_2_n_0 ),
        .I1(\m100.u0/ethc0/v[writeok]1 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][1] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I4(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I5(\m100.u0/ethc0/r_reg[ecnt_n_0_][0] ),
        .O(\m100.u0/ethc0/v[udpsrc] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1000)) 
    \r[udpsrc][15]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[edclrstate] [1]),
        .I1(\m100.u0/ethc0/r_reg[edclrstate] [3]),
        .I2(\m100.u0/ethc0/r_reg[edclrstate] [0]),
        .I3(\m100.u0/ethc0/r_reg[edclrstate] [2]),
        .O(\r[udpsrc][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r[udpsrc][15]_i_3 
       (.I0(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I1(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .O(\m100.u0/ethc0/v[writeok]1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBF80)) 
    \r[write][0]_i_1 
       (.I0(\m100.u0/rxwdata [17]),
        .I1(\r[udpsrc][15]_i_2_n_0 ),
        .I2(\r[write][0]_i_2_n_0 ),
        .I3(\m100.u0/ethc0/r_reg[write_n_0_][0] ),
        .O(\r[write][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \r[write][0]_i_2 
       (.I0(\m100.u0/ethc0/v[writeok]1 ),
        .I1(\r[ecnt][3]_i_3_n_0 ),
        .I2(\m100.u0/ethc0/r_reg[ecnt_n_0_][2] ),
        .I3(\m100.u0/ethc0/r_reg[ecnt_n_0_][3] ),
        .I4(\m100.u0/ewaddressm [7]),
        .I5(\m100.u0/ewaddressm [8]),
        .O(\r[write][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBFFFFFF08000000)) 
    \r[write][1]_i_1 
       (.I0(\m100.u0/rxwdata [17]),
        .I1(\r[udpsrc][15]_i_2_n_0 ),
        .I2(\m100.u0/ewaddressm [8]),
        .I3(\m100.u0/ewaddressm [7]),
        .I4(\r[ewr]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[write_n_0_][1] ),
        .O(\r[write][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBFFFFFF08000000)) 
    \r[write][2]_i_1 
       (.I0(\m100.u0/rxwdata [17]),
        .I1(\r[udpsrc][15]_i_2_n_0 ),
        .I2(\m100.u0/ewaddressm [7]),
        .I3(\m100.u0/ewaddressm [8]),
        .I4(\r[ewr]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[write_n_0_][2] ),
        .O(\r[write][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFFFFFF80000000)) 
    \r[write][3]_i_1 
       (.I0(\m100.u0/rxwdata [17]),
        .I1(\r[udpsrc][15]_i_2_n_0 ),
        .I2(\m100.u0/ewaddressm [7]),
        .I3(\m100.u0/ewaddressm [8]),
        .I4(\r[ewr]_i_2_n_0 ),
        .I5(\m100.u0/ethc0/r_reg[write_n_0_][3] ),
        .O(\r[write][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD7D7D71414141414)) 
    \r[writeok]_i_2 
       (.I0(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .I1(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I2(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I3(\m100.u0/ethc0/r_reg[rxdstate] [2]),
        .I4(\m100.u0/ethc0/r_reg[rxdoneold]__1 ),
        .I5(\m100.u0/ethc0/p_0_in153_in ),
        .O(\r[writeok]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[addrok]_i_4 
       (.CI(\r_reg[addrok]_i_5_n_0 ),
        .CO(r_reg),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .S({etho,etho,\r[addrok]_i_6_n_0 ,\r[addrok]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[addrok]_i_5 
       (.CI(etho),
        .CO({\r_reg[addrok]_i_5_n_0 ,\r_reg[addrok]_i_5_n_1 ,\r_reg[addrok]_i_5_n_2 ,\r_reg[addrok]_i_5_n_3 }),
        .CYINIT(apbo),
        .DI({etho,etho,etho,etho}),
        .S({\r[addrok]_i_8_n_0 ,\r[addrok]_i_9_n_0 ,\r[addrok]_i_10_n_0 ,\r[addrok]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[edclactive]_i_6 
       (.CI(\r_reg[edclactive]_i_7_n_0 ),
        .CO({\r_reg[edclactive]_i_6_n_0 ,\r_reg[edclactive]_i_6_n_1 ,\r_reg[edclactive]_i_6_n_2 ,\r_reg[edclactive]_i_6_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,apbo,apbo}),
        .S({etho,etho,\r[edclactive]_i_8_n_0 ,\r[edclactive]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[edclactive]_i_7 
       (.CI(etho),
        .CO({\r_reg[edclactive]_i_7_n_0 ,\r_reg[edclactive]_i_7_n_1 ,\r_reg[edclactive]_i_7_n_2 ,\r_reg[edclactive]_i_7_n_3 }),
        .CYINIT(etho),
        .DI({apbo,apbo,apbo,apbo}),
        .S({\r[edclactive]_i_10_n_0 ,\r[edclactive]_i_11_n_0 ,\r[edclactive]_i_12_n_0 ,\r[edclactive]_i_13_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[ipcrc][11]_i_2 
       (.CI(\r_reg[ipcrc][7]_i_2_n_0 ),
        .CO({\r_reg[ipcrc][11]_i_2_n_0 ,\r_reg[ipcrc][11]_i_2_n_1 ,\r_reg[ipcrc][11]_i_2_n_2 ,\r_reg[ipcrc][11]_i_2_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O(\m100.u0/ethc0/crcadder [11:8]),
        .S({\m100.u0/ethc0/r_reg[ipcrc_n_0_][11] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][10] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][9] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][8] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[ipcrc][11]_i_3 
       (.CI(\r_reg[ipcrc][7]_i_3_n_0 ),
        .CO({\r_reg[ipcrc][11]_i_3_n_0 ,\r_reg[ipcrc][11]_i_3_n_1 ,\r_reg[ipcrc][11]_i_3_n_2 ,\r_reg[ipcrc][11]_i_3_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/r_reg[ipcrc_n_0_][11] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][10] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][9] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][8] }),
        .O(\m100.u0/ethc0/p_1_in [11:8]),
        .S({\r[ipcrc][11]_i_8_n_0 ,\r[ipcrc][11]_i_9_n_0 ,\r[ipcrc][11]_i_10_n_0 ,\r[ipcrc][11]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[ipcrc][15]_i_2 
       (.CI(\r_reg[ipcrc][11]_i_2_n_0 ),
        .CO({\r_reg[ipcrc][15]_i_2_n_0 ,\r_reg[ipcrc][15]_i_2_n_1 ,\r_reg[ipcrc][15]_i_2_n_2 ,\r_reg[ipcrc][15]_i_2_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O(\m100.u0/ethc0/crcadder [15:12]),
        .S({\m100.u0/ethc0/r_reg[ipcrc_n_0_][15] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][14] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][13] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][12] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[ipcrc][15]_i_3 
       (.CI(\r_reg[ipcrc][11]_i_3_n_0 ),
        .CO({\r_reg[ipcrc][15]_i_3_n_0 ,\r_reg[ipcrc][15]_i_3_n_1 ,\r_reg[ipcrc][15]_i_3_n_2 ,\r_reg[ipcrc][15]_i_3_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/r_reg[ipcrc_n_0_][15] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][14] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][13] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][12] }),
        .O(\m100.u0/ethc0/p_1_in [15:12]),
        .S({\r[ipcrc][15]_i_8_n_0 ,\r[ipcrc][15]_i_9_n_0 ,\r[ipcrc][15]_i_10_n_0 ,\r[ipcrc][15]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[ipcrc][16]_i_2 
       (.CI(\r_reg[ipcrc][15]_i_2_n_0 ),
        .CO({\r_reg[ipcrc][16]_i_2_n_0 ,\r_reg[ipcrc][16]_i_2_n_1 ,\r_reg[ipcrc][16]_i_2_n_2 ,\m100.u0/ethc0/crcadder [16]}),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .S({etho,etho,etho,apbo}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[ipcrc][17]_i_4 
       (.CI(\r_reg[ipcrc][15]_i_3_n_0 ),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[ipcrc][17]_i_4_n_4 ,\r_reg[ipcrc][17]_i_4_n_5 ,\m100.u0/ethc0/p_1_in [17:16]}),
        .S({etho,etho,\m100.u0/ethc0/a }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[ipcrc][3]_i_2 
       (.CI(etho),
        .CO({\r_reg[ipcrc][3]_i_2_n_0 ,\r_reg[ipcrc][3]_i_2_n_1 ,\r_reg[ipcrc][3]_i_2_n_2 ,\r_reg[ipcrc][3]_i_2_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,\m100.u0/ethc0/a }),
        .O(\m100.u0/ethc0/crcadder [3:0]),
        .S({\m100.u0/ethc0/r_reg[ipcrc_n_0_][3] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][2] ,\r[ipcrc][3]_i_6_n_0 ,\r[ipcrc][3]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[ipcrc][3]_i_3 
       (.CI(etho),
        .CO({\r_reg[ipcrc][3]_i_3_n_0 ,\r_reg[ipcrc][3]_i_3_n_1 ,\r_reg[ipcrc][3]_i_3_n_2 ,\r_reg[ipcrc][3]_i_3_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/r_reg[ipcrc_n_0_][3] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][2] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][1] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][0] }),
        .O(\m100.u0/ethc0/p_1_in [3:0]),
        .S({\r[ipcrc][3]_i_8_n_0 ,\r[ipcrc][3]_i_9_n_0 ,\r[ipcrc][3]_i_10_n_0 ,\r[ipcrc][3]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[ipcrc][7]_i_2 
       (.CI(\r_reg[ipcrc][3]_i_2_n_0 ),
        .CO({\r_reg[ipcrc][7]_i_2_n_0 ,\r_reg[ipcrc][7]_i_2_n_1 ,\r_reg[ipcrc][7]_i_2_n_2 ,\r_reg[ipcrc][7]_i_2_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O(\m100.u0/ethc0/crcadder [7:4]),
        .S({\m100.u0/ethc0/r_reg[ipcrc_n_0_][7] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][6] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][5] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][4] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[ipcrc][7]_i_3 
       (.CI(\r_reg[ipcrc][3]_i_3_n_0 ),
        .CO({\r_reg[ipcrc][7]_i_3_n_0 ,\r_reg[ipcrc][7]_i_3_n_1 ,\r_reg[ipcrc][7]_i_3_n_2 ,\r_reg[ipcrc][7]_i_3_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/r_reg[ipcrc_n_0_][7] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][6] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][5] ,\m100.u0/ethc0/r_reg[ipcrc_n_0_][4] }),
        .O(\m100.u0/ethc0/p_1_in [7:4]),
        .S({\r[ipcrc][7]_i_8_n_0 ,\r[ipcrc][7]_i_9_n_0 ,\r[ipcrc][7]_i_10_n_0 ,\r[ipcrc][7]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_reg[mdio_ctrl][write]_i_2 
       (.I0(\r[mdio_ctrl][write]_i_6_n_0 ),
        .I1(\r[mdio_ctrl][write]_i_7_n_0 ),
        .O(\r_reg[mdio_ctrl][write]_i_2_n_0 ),
        .S(\m100.u0/ethc0/r_reg[mdio_state] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_reg[mdioo]_i_5 
       (.I0(\r[mdioo]_i_13_n_0 ),
        .I1(\r[mdioo]_i_14_n_0 ),
        .O(\r_reg[mdioo]_i_5_n_0 ),
        .S(\m100.u0/ethc0/r_reg[mdio_state] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[msbgood]_i_10 
       (.CI(etho),
        .CO({\r_reg[msbgood]_i_10_n_0 ,\r_reg[msbgood]_i_10_n_1 ,\r_reg[msbgood]_i_10_n_2 ,\r_reg[msbgood]_i_10_n_3 }),
        .CYINIT(apbo),
        .DI({etho,etho,etho,etho}),
        .S({\r[msbgood]_i_15_n_0 ,\r[msbgood]_i_16_n_0 ,\r[msbgood]_i_17_n_0 ,\r[msbgood]_i_18_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[msbgood]_i_3 
       (.CI(\r_reg[msbgood]_i_5_n_0 ),
        .CO({\r_reg[msbgood]_i_3_n_0 ,\r_reg[msbgood]_i_3_n_1 ,\r_reg[msbgood]_i_3_n_2 ,\r_reg[msbgood]_i_3_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .S({etho,\r[msbgood]_i_6_n_0 ,\r[msbgood]_i_7_n_0 ,\r[msbgood]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[msbgood]_i_5 
       (.CI(\r_reg[msbgood]_i_10_n_0 ),
        .CO({\r_reg[msbgood]_i_5_n_0 ,\r_reg[msbgood]_i_5_n_1 ,\r_reg[msbgood]_i_5_n_2 ,\r_reg[msbgood]_i_5_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .S({\r[msbgood]_i_11_n_0 ,\r[msbgood]_i_12_n_0 ,\r[msbgood]_i_13_n_0 ,\r[msbgood]_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[nak]_i_2 
       (.CI(\r_reg[nak]_i_3_n_0 ),
        .CO({\r_reg[nak]_i_2_n_0 ,\r_reg[nak]_i_2_n_1 ,\r_reg[nak]_i_2_n_2 ,\m100.u0/ethc0/v[nak]1 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .S({etho,etho,etho,\r[nak]_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[nak]_i_3 
       (.CI(etho),
        .CO({\r_reg[nak]_i_3_n_0 ,\r_reg[nak]_i_3_n_1 ,\r_reg[nak]_i_3_n_2 ,\r_reg[nak]_i_3_n_3 }),
        .CYINIT(apbo),
        .DI({etho,etho,etho,etho}),
        .S({\r[nak]_i_5_n_0 ,\r[nak]_i_6_n_0 ,\r[nak]_i_7_n_0 ,\r[nak]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_reg[rfrpnt][0]_i_1 
       (.I0(\r[rfrpnt][0]_i_2_n_0 ),
        .I1(\r[rfrpnt][0]_i_3_n_0 ),
        .O(\m100.u0/rxraddress [0]),
        .S(\m100.u0/ethc0/r_reg[rxdstate] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][13]_i_1 
       (.CI(\r_reg[rmsto][addr][9]_i_1_n_0 ),
        .CO({\r_reg[rmsto][addr][13]_i_1_n_0 ,\r_reg[rmsto][addr][13]_i_1_n_1 ,\r_reg[rmsto][addr][13]_i_1_n_2 ,\r_reg[rmsto][addr][13]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] }),
        .O({\r_reg[rmsto][addr][13]_i_1_n_4 ,\r_reg[rmsto][addr][13]_i_1_n_5 ,\r_reg[rmsto][addr][13]_i_1_n_6 ,\r_reg[rmsto][addr][13]_i_1_n_7 }),
        .S({\r[rmsto][addr][13]_i_2_n_0 ,\r[rmsto][addr][13]_i_3_n_0 ,\r[rmsto][addr][13]_i_4_n_0 ,\r[rmsto][addr][13]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][13]_i_10 
       (.CI(\r_reg[rmsto][addr][9]_i_10_n_0 ),
        .CO({\r_reg[rmsto][addr][13]_i_10_n_0 ,\r_reg[rmsto][addr][13]_i_10_n_1 ,\r_reg[rmsto][addr][13]_i_10_n_2 ,\r_reg[rmsto][addr][13]_i_10_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[rmsto][addr][13]_i_10_n_4 ,\r_reg[rmsto][addr][13]_i_10_n_5 ,\r_reg[rmsto][addr][13]_i_10_n_6 ,\r_reg[rmsto][addr][13]_i_10_n_7 }),
        .S(\m100.u0/ethc0/r_reg[rmsto][addr] [16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][17]_i_1 
       (.CI(\r_reg[rmsto][addr][13]_i_1_n_0 ),
        .CO({\r_reg[rmsto][addr][17]_i_1_n_0 ,\r_reg[rmsto][addr][17]_i_1_n_1 ,\r_reg[rmsto][addr][17]_i_1_n_2 ,\r_reg[rmsto][addr][17]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] }),
        .O({\r_reg[rmsto][addr][17]_i_1_n_4 ,\r_reg[rmsto][addr][17]_i_1_n_5 ,\r_reg[rmsto][addr][17]_i_1_n_6 ,\r_reg[rmsto][addr][17]_i_1_n_7 }),
        .S({\r[rmsto][addr][17]_i_2_n_0 ,\r[rmsto][addr][17]_i_3_n_0 ,\r[rmsto][addr][17]_i_4_n_0 ,\r[rmsto][addr][17]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][17]_i_10 
       (.CI(\r_reg[rmsto][addr][13]_i_10_n_0 ),
        .CO({\r_reg[rmsto][addr][17]_i_10_n_0 ,\r_reg[rmsto][addr][17]_i_10_n_1 ,\r_reg[rmsto][addr][17]_i_10_n_2 ,\r_reg[rmsto][addr][17]_i_10_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[rmsto][addr][17]_i_10_n_4 ,\r_reg[rmsto][addr][17]_i_10_n_5 ,\r_reg[rmsto][addr][17]_i_10_n_6 ,\r_reg[rmsto][addr][17]_i_10_n_7 }),
        .S(\m100.u0/ethc0/r_reg[rmsto][addr] [20:17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][1]_i_10 
       (.CI(etho),
        .CO({\r_reg[rmsto][addr][1]_i_10_n_0 ,\r_reg[rmsto][addr][1]_i_10_n_1 ,\r_reg[rmsto][addr][1]_i_10_n_2 ,\r_reg[rmsto][addr][1]_i_10_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,\m100.u0/ethc0/r_reg[rmsto][addr] [2],etho}),
        .O({\r_reg[rmsto][addr][1]_i_10_n_4 ,\r_reg[rmsto][addr][1]_i_10_n_5 ,\r_reg[rmsto][addr][1]_i_10_n_6 ,\r_reg[rmsto][addr][1]_i_10_n_7 }),
        .S({\m100.u0/ethc0/r_reg[rmsto][addr] [4:3],\r[rmsto][addr][1]_i_13_n_0 ,\m100.u0/ethc0/r_reg[rmsto][addr] [1]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][1]_i_2 
       (.CI(etho),
        .CO({\r_reg[rmsto][addr][1]_i_2_n_0 ,\r_reg[rmsto][addr][1]_i_2_n_1 ,\r_reg[rmsto][addr][1]_i_2_n_2 ,\r_reg[rmsto][addr][1]_i_2_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,etho}),
        .O({\r_reg[rmsto][addr][1]_i_2_n_4 ,\r_reg[rmsto][addr][1]_i_2_n_5 ,\r_reg[rmsto][addr][1]_i_2_n_6 ,\r_reg[rmsto][addr][1]_i_2_n_7 }),
        .S({\r[rmsto][addr][1]_i_3_n_0 ,\r[rmsto][addr][1]_i_4_n_0 ,\r[rmsto][addr][1]_i_5_n_0 ,\r[rmsto][addr][1]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][21]_i_1 
       (.CI(\r_reg[rmsto][addr][17]_i_1_n_0 ),
        .CO({\r_reg[rmsto][addr][21]_i_1_n_0 ,\r_reg[rmsto][addr][21]_i_1_n_1 ,\r_reg[rmsto][addr][21]_i_1_n_2 ,\r_reg[rmsto][addr][21]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] }),
        .O({\r_reg[rmsto][addr][21]_i_1_n_4 ,\r_reg[rmsto][addr][21]_i_1_n_5 ,\r_reg[rmsto][addr][21]_i_1_n_6 ,\r_reg[rmsto][addr][21]_i_1_n_7 }),
        .S({\r[rmsto][addr][21]_i_2_n_0 ,\r[rmsto][addr][21]_i_3_n_0 ,\r[rmsto][addr][21]_i_4_n_0 ,\r[rmsto][addr][21]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][21]_i_10 
       (.CI(\r_reg[rmsto][addr][17]_i_10_n_0 ),
        .CO({\r_reg[rmsto][addr][21]_i_10_n_0 ,\r_reg[rmsto][addr][21]_i_10_n_1 ,\r_reg[rmsto][addr][21]_i_10_n_2 ,\r_reg[rmsto][addr][21]_i_10_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[rmsto][addr][21]_i_10_n_4 ,\r_reg[rmsto][addr][21]_i_10_n_5 ,\r_reg[rmsto][addr][21]_i_10_n_6 ,\r_reg[rmsto][addr][21]_i_10_n_7 }),
        .S(\m100.u0/ethc0/r_reg[rmsto][addr] [24:21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][25]_i_1 
       (.CI(\r_reg[rmsto][addr][21]_i_1_n_0 ),
        .CO({\r_reg[rmsto][addr][25]_i_1_n_0 ,\r_reg[rmsto][addr][25]_i_1_n_1 ,\r_reg[rmsto][addr][25]_i_1_n_2 ,\r_reg[rmsto][addr][25]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] }),
        .O({\r_reg[rmsto][addr][25]_i_1_n_4 ,\r_reg[rmsto][addr][25]_i_1_n_5 ,\r_reg[rmsto][addr][25]_i_1_n_6 ,\r_reg[rmsto][addr][25]_i_1_n_7 }),
        .S({\r[rmsto][addr][25]_i_2_n_0 ,\r[rmsto][addr][25]_i_3_n_0 ,\r[rmsto][addr][25]_i_4_n_0 ,\r[rmsto][addr][25]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][25]_i_10 
       (.CI(\r_reg[rmsto][addr][21]_i_10_n_0 ),
        .CO({\r_reg[rmsto][addr][25]_i_10_n_0 ,\r_reg[rmsto][addr][25]_i_10_n_1 ,\r_reg[rmsto][addr][25]_i_10_n_2 ,\r_reg[rmsto][addr][25]_i_10_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[rmsto][addr][25]_i_10_n_4 ,\r_reg[rmsto][addr][25]_i_10_n_5 ,\r_reg[rmsto][addr][25]_i_10_n_6 ,\r_reg[rmsto][addr][25]_i_10_n_7 }),
        .S(\m100.u0/ethc0/r_reg[rmsto][addr] [28:25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][29]_i_1 
       (.CI(\r_reg[rmsto][addr][25]_i_1_n_0 ),
        .CYINIT(etho),
        .DI({etho,etho,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] }),
        .O({\r_reg[rmsto][addr][29]_i_1_n_4 ,\r_reg[rmsto][addr][29]_i_1_n_5 ,\r_reg[rmsto][addr][29]_i_1_n_6 ,\r_reg[rmsto][addr][29]_i_1_n_7 }),
        .S({etho,\r[rmsto][addr][29]_i_2_n_0 ,\r[rmsto][addr][29]_i_3_n_0 ,\r[rmsto][addr][29]_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][29]_i_8 
       (.CI(\r_reg[rmsto][addr][25]_i_10_n_0 ),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[rmsto][addr][29]_i_8_n_4 ,\r_reg[rmsto][addr][29]_i_8_n_5 ,\r_reg[rmsto][addr][29]_i_8_n_6 ,\r_reg[rmsto][addr][29]_i_8_n_7 }),
        .S({etho,\m100.u0/ethc0/r_reg[rmsto][addr] [31:29]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][5]_i_1 
       (.CI(\r_reg[rmsto][addr][1]_i_2_n_0 ),
        .CO({\r_reg[rmsto][addr][5]_i_1_n_0 ,\r_reg[rmsto][addr][5]_i_1_n_1 ,\r_reg[rmsto][addr][5]_i_1_n_2 ,\r_reg[rmsto][addr][5]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] }),
        .O({\r_reg[rmsto][addr][5]_i_1_n_4 ,\r_reg[rmsto][addr][5]_i_1_n_5 ,\r_reg[rmsto][addr][5]_i_1_n_6 ,\r_reg[rmsto][addr][5]_i_1_n_7 }),
        .S({\r[rmsto][addr][5]_i_2_n_0 ,\r[rmsto][addr][5]_i_3_n_0 ,\r[rmsto][addr][5]_i_4_n_0 ,\r[rmsto][addr][5]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][5]_i_10 
       (.CI(\r_reg[rmsto][addr][1]_i_10_n_0 ),
        .CO({\r_reg[rmsto][addr][5]_i_10_n_0 ,\r_reg[rmsto][addr][5]_i_10_n_1 ,\r_reg[rmsto][addr][5]_i_10_n_2 ,\r_reg[rmsto][addr][5]_i_10_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[rmsto][addr][5]_i_10_n_4 ,\r_reg[rmsto][addr][5]_i_10_n_5 ,\r_reg[rmsto][addr][5]_i_10_n_6 ,\r_reg[rmsto][addr][5]_i_10_n_7 }),
        .S(\m100.u0/ethc0/r_reg[rmsto][addr] [8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][9]_i_1 
       (.CI(\r_reg[rmsto][addr][5]_i_1_n_0 ),
        .CO({\r_reg[rmsto][addr][9]_i_1_n_0 ,\r_reg[rmsto][addr][9]_i_1_n_1 ,\r_reg[rmsto][addr][9]_i_1_n_2 ,\r_reg[rmsto][addr][9]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] ,\m100.u0/ethc0/rmsti[retry] }),
        .O({\r_reg[rmsto][addr][9]_i_1_n_4 ,\r_reg[rmsto][addr][9]_i_1_n_5 ,\r_reg[rmsto][addr][9]_i_1_n_6 ,\r_reg[rmsto][addr][9]_i_1_n_7 }),
        .S({\r[rmsto][addr][9]_i_2_n_0 ,\r[rmsto][addr][9]_i_3_n_0 ,\r[rmsto][addr][9]_i_4_n_0 ,\r[rmsto][addr][9]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][addr][9]_i_10 
       (.CI(\r_reg[rmsto][addr][5]_i_10_n_0 ),
        .CO({\r_reg[rmsto][addr][9]_i_10_n_0 ,\r_reg[rmsto][addr][9]_i_10_n_1 ,\r_reg[rmsto][addr][9]_i_10_n_2 ,\r_reg[rmsto][addr][9]_i_10_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[rmsto][addr][9]_i_10_n_4 ,\r_reg[rmsto][addr][9]_i_10_n_5 ,\r_reg[rmsto][addr][9]_i_10_n_6 ,\r_reg[rmsto][addr][9]_i_10_n_7 }),
        .S(\m100.u0/ethc0/r_reg[rmsto][addr] [12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][req]_i_10 
       (.CI(etho),
        .CO({\r_reg[rmsto][req]_i_10_n_0 ,\r_reg[rmsto][req]_i_10_n_1 ,\r_reg[rmsto][req]_i_10_n_2 ,\r_reg[rmsto][req]_i_10_n_3 }),
        .CYINIT(apbo),
        .DI({\r[rmsto][req]_i_20_n_0 ,\r[rmsto][req]_i_21_n_0 ,\r[rmsto][req]_i_22_n_0 ,\r[rmsto][req]_i_23_n_0 }),
        .S({\r[rmsto][req]_i_24_n_0 ,\r[rmsto][req]_i_25_n_0 ,\r[rmsto][req]_i_26_n_0 ,\r[rmsto][req]_i_27_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][req]_i_15 
       (.CI(etho),
        .CO({\r_reg[rmsto][req]_i_15_n_0 ,\r_reg[rmsto][req]_i_15_n_1 ,\r_reg[rmsto][req]_i_15_n_2 ,\r_reg[rmsto][req]_i_15_n_3 }),
        .CYINIT(apbo),
        .DI({\r[rmsto][req]_i_30_n_0 ,\r[rmsto][req]_i_31_n_0 ,\r[rmsto][req]_i_32_n_0 ,\r[rmsto][req]_i_33_n_0 }),
        .S({\r[rmsto][req]_i_34_n_0 ,\r[rmsto][req]_i_35_n_0 ,\r[rmsto][req]_i_36_n_0 ,\r[rmsto][req]_i_37_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][req]_i_8 
       (.CI(\r_reg[rmsto][req]_i_10_n_0 ),
        .CO({\r_reg[rmsto][req]_i_8_n_0 ,\r_reg[rmsto][req]_i_8_n_1 ,\m100.u0/ethc0/v[rmsto][req]2136_in ,\r_reg[rmsto][req]_i_8_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,\r[rmsto][req]_i_11_n_0 ,\r[rmsto][req]_i_12_n_0 }),
        .S({etho,etho,\r[rmsto][req]_i_13_n_0 ,\r[rmsto][req]_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rmsto][req]_i_9 
       (.CI(\r_reg[rmsto][req]_i_15_n_0 ),
        .CO({\r_reg[rmsto][req]_i_9_n_0 ,\r_reg[rmsto][req]_i_9_n_1 ,\m100.u0/ethc0/v[rmsto][req]2137_in ,\r_reg[rmsto][req]_i_9_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,\r[rmsto][req]_i_16_n_0 ,\r[rmsto][req]_i_17_n_0 }),
        .S({etho,etho,\r[rmsto][req]_i_18_n_0 ,\r[rmsto][req]_i_19_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rxcnt][10]_i_8 
       (.CI(\r_reg[rxcnt][10]_i_9_n_0 ),
        .CO({\r_reg[rxcnt][10]_i_8_n_0 ,\r_reg[rxcnt][10]_i_8_n_1 ,\r_reg[rxcnt][10]_i_8_n_2 ,\r_reg[rxcnt][10]_i_8_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,\r[rxcnt][10]_i_10_n_0 ,\r[rxcnt][10]_i_11_n_0 }),
        .S({etho,etho,\r[rxcnt][10]_i_12_n_0 ,\r[rxcnt][10]_i_13_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[rxcnt][10]_i_9 
       (.CI(etho),
        .CO({\r_reg[rxcnt][10]_i_9_n_0 ,\r_reg[rxcnt][10]_i_9_n_1 ,\r_reg[rxcnt][10]_i_9_n_2 ,\r_reg[rxcnt][10]_i_9_n_3 }),
        .CYINIT(etho),
        .DI({\r[rxcnt][10]_i_14_n_0 ,\r[rxcnt][10]_i_15_n_0 ,\r[rxcnt][10]_i_16_n_0 ,\r[rxcnt][10]_i_17_n_0 }),
        .S({\r[rxcnt][10]_i_18_n_0 ,\r[rxcnt][10]_i_19_n_0 ,\r[rxcnt][10]_i_20_n_0 ,\r[rxcnt][10]_i_21_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[rxstatus][4]_i_4 
       (.CI(etho),
        .CO({\m100.u0/ethc0/v[rxstatus]2130_in ,\r_reg[rxstatus][4]_i_4_n_1 ,\r_reg[rxstatus][4]_i_4_n_2 ,\r_reg[rxstatus][4]_i_4_n_3 }),
        .CYINIT(etho),
        .DI({apbo,apbo,apbo,apbo}),
        .S({\r[rxstatus][4]_i_12_n_0 ,\r[rxstatus][4]_i_13_n_0 ,\r[rxstatus][4]_i_14_n_0 ,\r[rxstatus][4]_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[seq][0]_i_2 
       (.CI(etho),
        .CO({\r_reg[seq][0]_i_2_n_0 ,\r_reg[seq][0]_i_2_n_1 ,\r_reg[seq][0]_i_2_n_2 ,\r_reg[seq][0]_i_2_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,apbo}),
        .O({\r_reg[seq][0]_i_2_n_4 ,\r_reg[seq][0]_i_2_n_5 ,\r_reg[seq][0]_i_2_n_6 ,\r_reg[seq][0]_i_2_n_7 }),
        .S({\m100.u0/ethc0/r_reg[seq] [3:1],\r[seq][0]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[seq][12]_i_1 
       (.CI(\r_reg[seq][8]_i_1_n_0 ),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[seq][12]_i_1_n_4 ,\r_reg[seq][12]_i_1_n_5 ,\r_reg[seq][12]_i_1_n_6 ,\r_reg[seq][12]_i_1_n_7 }),
        .S({etho,etho,\m100.u0/ethc0/r_reg[seq] [13:12]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[seq][4]_i_1 
       (.CI(\r_reg[seq][0]_i_2_n_0 ),
        .CO({\r_reg[seq][4]_i_1_n_0 ,\r_reg[seq][4]_i_1_n_1 ,\r_reg[seq][4]_i_1_n_2 ,\r_reg[seq][4]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[seq][4]_i_1_n_4 ,\r_reg[seq][4]_i_1_n_5 ,\r_reg[seq][4]_i_1_n_6 ,\r_reg[seq][4]_i_1_n_7 }),
        .S(\m100.u0/ethc0/r_reg[seq] [7:4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[seq][8]_i_1 
       (.CI(\r_reg[seq][4]_i_1_n_0 ),
        .CO({\r_reg[seq][8]_i_1_n_0 ,\r_reg[seq][8]_i_1_n_1 ,\r_reg[seq][8]_i_1_n_2 ,\r_reg[seq][8]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[seq][8]_i_1_n_4 ,\r_reg[seq][8]_i_1_n_5 ,\r_reg[seq][8]_i_1_n_6 ,\r_reg[seq][8]_i_1_n_7 }),
        .S(\m100.u0/ethc0/r_reg[seq] [11:8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[status][toosmall]_i_5 
       (.CI(\r_reg[status][toosmall]_i_6_n_0 ),
        .CO({\r_reg[status][toosmall]_i_5_n_0 ,\r_reg[status][toosmall]_i_5_n_1 ,\m100.u0/ethc0/v[status][toosmall]2 ,\r_reg[status][toosmall]_i_5_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,\r[status][toosmall]_i_7_n_0 ,\r[status][toosmall]_i_8_n_0 }),
        .S({etho,etho,\r[status][toosmall]_i_9_n_0 ,\r[status][toosmall]_i_10_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[status][toosmall]_i_6 
       (.CI(etho),
        .CO({\r_reg[status][toosmall]_i_6_n_0 ,\r_reg[status][toosmall]_i_6_n_1 ,\r_reg[status][toosmall]_i_6_n_2 ,\r_reg[status][toosmall]_i_6_n_3 }),
        .CYINIT(apbo),
        .DI({\r[status][toosmall]_i_11_n_0 ,\r[status][toosmall]_i_12_n_0 ,\r[status][toosmall]_i_13_n_0 ,\r[status][toosmall]_i_14_n_0 }),
        .S({\r[status][toosmall]_i_15_n_0 ,\r[status][toosmall]_i_16_n_0 ,\r[status][toosmall]_i_17_n_0 ,\r[status][toosmall]_i_18_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tfcnt][3]_i_2 
       (.CI(etho),
        .CO({\r_reg[tfcnt][3]_i_2_n_0 ,\r_reg[tfcnt][3]_i_2_n_1 ,\r_reg[tfcnt][3]_i_2_n_2 ,\r_reg[tfcnt][3]_i_2_n_3 }),
        .CYINIT(etho),
        .DI({\r[tfcnt][3]_i_4_n_0 ,\r[tfcnt][3]_i_5_n_0 ,\r[tfcnt][3]_i_6_n_0 ,\r[tfcnt][3]_i_7_n_0 }),
        .O({\r_reg[tfcnt][3]_i_2_n_4 ,\r_reg[tfcnt][3]_i_2_n_5 ,\r_reg[tfcnt][3]_i_2_n_6 ,\r_reg[tfcnt][3]_i_2_n_7 }),
        .S({\r[tfcnt][3]_i_8_n_0 ,\r[tfcnt][3]_i_9_n_0 ,\r[tfcnt][3]_i_10_n_0 ,\r[tfcnt][3]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tfcnt][3]_i_3 
       (.CI(etho),
        .CO({\r_reg[tfcnt][3]_i_3_n_0 ,\r_reg[tfcnt][3]_i_3_n_1 ,\r_reg[tfcnt][3]_i_3_n_2 ,\r_reg[tfcnt][3]_i_3_n_3 }),
        .CYINIT(apbo),
        .DI({\r[tfcnt][3]_i_4_n_0 ,\r[tfcnt][3]_i_12_n_0 ,\r[tfcnt][3]_i_13_n_0 ,\r[tfcnt][3]_i_14_n_0 }),
        .O({\r_reg[tfcnt][3]_i_3_n_4 ,\r_reg[tfcnt][3]_i_3_n_5 ,\r_reg[tfcnt][3]_i_3_n_6 ,\r_reg[tfcnt][3]_i_3_n_7 }),
        .S({\r[tfcnt][3]_i_15_n_0 ,\r[tfcnt][3]_i_16_n_0 ,\r[tfcnt][3]_i_17_n_0 ,\r[tfcnt][3]_i_18_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tfcnt][7]_i_2 
       (.CI(\r_reg[tfcnt][3]_i_2_n_0 ),
        .CYINIT(etho),
        .DI({etho,\r[tfcnt][7]_i_5_n_0 ,\r[tfcnt][7]_i_6_n_0 ,\r[tfcnt][7]_i_7_n_0 }),
        .O({\r_reg[tfcnt][7]_i_2_n_4 ,\r_reg[tfcnt][7]_i_2_n_5 ,\r_reg[tfcnt][7]_i_2_n_6 ,\r_reg[tfcnt][7]_i_2_n_7 }),
        .S({\r[tfcnt][7]_i_8_n_0 ,\r[tfcnt][7]_i_9_n_0 ,\r[tfcnt][7]_i_10_n_0 ,\r[tfcnt][7]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tfcnt][7]_i_4 
       (.CI(\r_reg[tfcnt][3]_i_3_n_0 ),
        .CYINIT(etho),
        .DI({etho,\r[tfcnt][7]_i_5_n_0 ,\r[tfcnt][7]_i_6_n_0 ,\r[tfcnt][7]_i_7_n_0 }),
        .O({\r_reg[tfcnt][7]_i_4_n_4 ,\r_reg[tfcnt][7]_i_4_n_5 ,\r_reg[tfcnt][7]_i_4_n_6 ,\r_reg[tfcnt][7]_i_4_n_7 }),
        .S({\r[tfcnt][7]_i_12_n_0 ,\r[tfcnt][7]_i_13_n_0 ,\r[tfcnt][7]_i_14_n_0 ,\r[tfcnt][7]_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][13]_i_1 
       (.CI(\r_reg[tmsto][addr][9]_i_1_n_0 ),
        .CO({\r_reg[tmsto][addr][13]_i_1_n_0 ,\r_reg[tmsto][addr][13]_i_1_n_1 ,\r_reg[tmsto][addr][13]_i_1_n_2 ,\r_reg[tmsto][addr][13]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] }),
        .O({\r_reg[tmsto][addr][13]_i_1_n_4 ,\r_reg[tmsto][addr][13]_i_1_n_5 ,\r_reg[tmsto][addr][13]_i_1_n_6 ,\r_reg[tmsto][addr][13]_i_1_n_7 }),
        .S({\r[tmsto][addr][13]_i_2_n_0 ,\r[tmsto][addr][13]_i_3_n_0 ,\r[tmsto][addr][13]_i_4_n_0 ,\r[tmsto][addr][13]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][13]_i_14 
       (.CI(\r_reg[tmsto][addr][9]_i_14_n_0 ),
        .CO({\r_reg[tmsto][addr][13]_i_14_n_0 ,\r_reg[tmsto][addr][13]_i_14_n_1 ,\r_reg[tmsto][addr][13]_i_14_n_2 ,\r_reg[tmsto][addr][13]_i_14_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[tmsto][addr][13]_i_14_n_4 ,\r_reg[tmsto][addr][13]_i_14_n_5 ,\r_reg[tmsto][addr][13]_i_14_n_6 ,\r_reg[tmsto][addr][13]_i_14_n_7 }),
        .S(\m100.u0/ethc0/r_reg[tmsto][addr] [16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][17]_i_1 
       (.CI(\r_reg[tmsto][addr][13]_i_1_n_0 ),
        .CO({\r_reg[tmsto][addr][17]_i_1_n_0 ,\r_reg[tmsto][addr][17]_i_1_n_1 ,\r_reg[tmsto][addr][17]_i_1_n_2 ,\r_reg[tmsto][addr][17]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] }),
        .O({\r_reg[tmsto][addr][17]_i_1_n_4 ,\r_reg[tmsto][addr][17]_i_1_n_5 ,\r_reg[tmsto][addr][17]_i_1_n_6 ,\r_reg[tmsto][addr][17]_i_1_n_7 }),
        .S({\r[tmsto][addr][17]_i_2_n_0 ,\r[tmsto][addr][17]_i_3_n_0 ,\r[tmsto][addr][17]_i_4_n_0 ,\r[tmsto][addr][17]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][17]_i_14 
       (.CI(\r_reg[tmsto][addr][13]_i_14_n_0 ),
        .CO({\r_reg[tmsto][addr][17]_i_14_n_0 ,\r_reg[tmsto][addr][17]_i_14_n_1 ,\r_reg[tmsto][addr][17]_i_14_n_2 ,\r_reg[tmsto][addr][17]_i_14_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[tmsto][addr][17]_i_14_n_4 ,\r_reg[tmsto][addr][17]_i_14_n_5 ,\r_reg[tmsto][addr][17]_i_14_n_6 ,\r_reg[tmsto][addr][17]_i_14_n_7 }),
        .S(\m100.u0/ethc0/r_reg[tmsto][addr] [20:17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][1]_i_17 
       (.CI(etho),
        .CO({\r_reg[tmsto][addr][1]_i_17_n_0 ,\r_reg[tmsto][addr][1]_i_17_n_1 ,\r_reg[tmsto][addr][1]_i_17_n_2 ,\r_reg[tmsto][addr][1]_i_17_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,\m100.u0/ethc0/r_reg[tmsto][addr] [2],etho}),
        .O({\r_reg[tmsto][addr][1]_i_17_n_4 ,\r_reg[tmsto][addr][1]_i_17_n_5 ,\r_reg[tmsto][addr][1]_i_17_n_6 ,\r_reg[tmsto][addr][1]_i_17_n_7 }),
        .S({\m100.u0/ethc0/r_reg[tmsto][addr] [4:3],\r[tmsto][addr][1]_i_25_n_0 ,\m100.u0/ethc0/r_reg[tmsto][addr] [1]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][1]_i_2 
       (.CI(etho),
        .CO({\r_reg[tmsto][addr][1]_i_2_n_0 ,\r_reg[tmsto][addr][1]_i_2_n_1 ,\r_reg[tmsto][addr][1]_i_2_n_2 ,\r_reg[tmsto][addr][1]_i_2_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,etho}),
        .O({\r_reg[tmsto][addr][1]_i_2_n_4 ,\r_reg[tmsto][addr][1]_i_2_n_5 ,\r_reg[tmsto][addr][1]_i_2_n_6 ,\r_reg[tmsto][addr][1]_i_2_n_7 }),
        .S({\r[tmsto][addr][1]_i_7_n_0 ,\r[tmsto][addr][1]_i_8_n_0 ,\r[tmsto][addr][1]_i_9_n_0 ,\r[tmsto][addr][1]_i_10_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][21]_i_1 
       (.CI(\r_reg[tmsto][addr][17]_i_1_n_0 ),
        .CO({\r_reg[tmsto][addr][21]_i_1_n_0 ,\r_reg[tmsto][addr][21]_i_1_n_1 ,\r_reg[tmsto][addr][21]_i_1_n_2 ,\r_reg[tmsto][addr][21]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] }),
        .O({\r_reg[tmsto][addr][21]_i_1_n_4 ,\r_reg[tmsto][addr][21]_i_1_n_5 ,\r_reg[tmsto][addr][21]_i_1_n_6 ,\r_reg[tmsto][addr][21]_i_1_n_7 }),
        .S({\r[tmsto][addr][21]_i_2_n_0 ,\r[tmsto][addr][21]_i_3_n_0 ,\r[tmsto][addr][21]_i_4_n_0 ,\r[tmsto][addr][21]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][21]_i_14 
       (.CI(\r_reg[tmsto][addr][17]_i_14_n_0 ),
        .CO({\r_reg[tmsto][addr][21]_i_14_n_0 ,\r_reg[tmsto][addr][21]_i_14_n_1 ,\r_reg[tmsto][addr][21]_i_14_n_2 ,\r_reg[tmsto][addr][21]_i_14_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[tmsto][addr][21]_i_14_n_4 ,\r_reg[tmsto][addr][21]_i_14_n_5 ,\r_reg[tmsto][addr][21]_i_14_n_6 ,\r_reg[tmsto][addr][21]_i_14_n_7 }),
        .S(\m100.u0/ethc0/r_reg[tmsto][addr] [24:21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][25]_i_1 
       (.CI(\r_reg[tmsto][addr][21]_i_1_n_0 ),
        .CO({\r_reg[tmsto][addr][25]_i_1_n_0 ,\r_reg[tmsto][addr][25]_i_1_n_1 ,\r_reg[tmsto][addr][25]_i_1_n_2 ,\r_reg[tmsto][addr][25]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] }),
        .O({\r_reg[tmsto][addr][25]_i_1_n_4 ,\r_reg[tmsto][addr][25]_i_1_n_5 ,\r_reg[tmsto][addr][25]_i_1_n_6 ,\r_reg[tmsto][addr][25]_i_1_n_7 }),
        .S({\r[tmsto][addr][25]_i_2_n_0 ,\r[tmsto][addr][25]_i_3_n_0 ,\r[tmsto][addr][25]_i_4_n_0 ,\r[tmsto][addr][25]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][25]_i_14 
       (.CI(\r_reg[tmsto][addr][21]_i_14_n_0 ),
        .CO({\r_reg[tmsto][addr][25]_i_14_n_0 ,\r_reg[tmsto][addr][25]_i_14_n_1 ,\r_reg[tmsto][addr][25]_i_14_n_2 ,\r_reg[tmsto][addr][25]_i_14_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[tmsto][addr][25]_i_14_n_4 ,\r_reg[tmsto][addr][25]_i_14_n_5 ,\r_reg[tmsto][addr][25]_i_14_n_6 ,\r_reg[tmsto][addr][25]_i_14_n_7 }),
        .S(\m100.u0/ethc0/r_reg[tmsto][addr] [28:25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][29]_i_1 
       (.CI(\r_reg[tmsto][addr][25]_i_1_n_0 ),
        .CYINIT(etho),
        .DI({etho,etho,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] }),
        .O({\r_reg[tmsto][addr][29]_i_1_n_4 ,\r_reg[tmsto][addr][29]_i_1_n_5 ,\r_reg[tmsto][addr][29]_i_1_n_6 ,\r_reg[tmsto][addr][29]_i_1_n_7 }),
        .S({etho,\r[tmsto][addr][29]_i_2_n_0 ,\r[tmsto][addr][29]_i_3_n_0 ,\r[tmsto][addr][29]_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][29]_i_11 
       (.CI(\r_reg[tmsto][addr][25]_i_14_n_0 ),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[tmsto][addr][29]_i_11_n_4 ,\r_reg[tmsto][addr][29]_i_11_n_5 ,\r_reg[tmsto][addr][29]_i_11_n_6 ,\r_reg[tmsto][addr][29]_i_11_n_7 }),
        .S({etho,\m100.u0/ethc0/r_reg[tmsto][addr] [31:29]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][5]_i_1 
       (.CI(\r_reg[tmsto][addr][1]_i_2_n_0 ),
        .CO({\r_reg[tmsto][addr][5]_i_1_n_0 ,\r_reg[tmsto][addr][5]_i_1_n_1 ,\r_reg[tmsto][addr][5]_i_1_n_2 ,\r_reg[tmsto][addr][5]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] }),
        .O({\r_reg[tmsto][addr][5]_i_1_n_4 ,\r_reg[tmsto][addr][5]_i_1_n_5 ,\r_reg[tmsto][addr][5]_i_1_n_6 ,\r_reg[tmsto][addr][5]_i_1_n_7 }),
        .S({\r[tmsto][addr][5]_i_2_n_0 ,\r[tmsto][addr][5]_i_3_n_0 ,\r[tmsto][addr][5]_i_4_n_0 ,\r[tmsto][addr][5]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][5]_i_14 
       (.CI(\r_reg[tmsto][addr][1]_i_17_n_0 ),
        .CO({\r_reg[tmsto][addr][5]_i_14_n_0 ,\r_reg[tmsto][addr][5]_i_14_n_1 ,\r_reg[tmsto][addr][5]_i_14_n_2 ,\r_reg[tmsto][addr][5]_i_14_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[tmsto][addr][5]_i_14_n_4 ,\r_reg[tmsto][addr][5]_i_14_n_5 ,\r_reg[tmsto][addr][5]_i_14_n_6 ,\r_reg[tmsto][addr][5]_i_14_n_7 }),
        .S(\m100.u0/ethc0/r_reg[tmsto][addr] [8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][9]_i_1 
       (.CI(\r_reg[tmsto][addr][5]_i_1_n_0 ),
        .CO({\r_reg[tmsto][addr][9]_i_1_n_0 ,\r_reg[tmsto][addr][9]_i_1_n_1 ,\r_reg[tmsto][addr][9]_i_1_n_2 ,\r_reg[tmsto][addr][9]_i_1_n_3 }),
        .CYINIT(etho),
        .DI({\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] ,\m100.u0/ethc0/tmsti[retry] }),
        .O({\r_reg[tmsto][addr][9]_i_1_n_4 ,\r_reg[tmsto][addr][9]_i_1_n_5 ,\r_reg[tmsto][addr][9]_i_1_n_6 ,\r_reg[tmsto][addr][9]_i_1_n_7 }),
        .S({\r[tmsto][addr][9]_i_2_n_0 ,\r[tmsto][addr][9]_i_3_n_0 ,\r[tmsto][addr][9]_i_4_n_0 ,\r[tmsto][addr][9]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_reg[tmsto][addr][9]_i_14 
       (.CI(\r_reg[tmsto][addr][5]_i_14_n_0 ),
        .CO({\r_reg[tmsto][addr][9]_i_14_n_0 ,\r_reg[tmsto][addr][9]_i_14_n_1 ,\r_reg[tmsto][addr][9]_i_14_n_2 ,\r_reg[tmsto][addr][9]_i_14_n_3 }),
        .CYINIT(etho),
        .DI({etho,etho,etho,etho}),
        .O({\r_reg[tmsto][addr][9]_i_14_n_4 ,\r_reg[tmsto][addr][9]_i_14_n_5 ,\r_reg[tmsto][addr][9]_i_14_n_6 ,\r_reg[tmsto][addr][9]_i_14_n_7 }),
        .S(\m100.u0/ethc0/r_reg[tmsto][addr] [12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_reg[tmsto][write]_i_2 
       (.I0(\r[tmsto][write]_i_6_n_0 ),
        .I1(\r[tmsto][write]_i_7_n_0 ),
        .O(\r_reg[tmsto][write]_i_2_n_0 ),
        .S(\m100.u0/ethc0/r_reg[txlength_n_0_][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_reg[txlength][7]_i_1 
       (.I0(\r[txlength][7]_i_2_n_0 ),
        .I1(\r[txlength][7]_i_3_n_0 ),
        .O(\r_reg[txlength][7]_i_1_n_0 ),
        .S(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_reg[txlength][9]_i_1 
       (.I0(\r[txlength][9]_i_2_n_0 ),
        .I1(\r[txlength][9]_i_3_n_0 ),
        .O(\r_reg[txlength][9]_i_1_n_0 ),
        .S(\m100.u0/ethc0/r_reg[txdstate_n_0_][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h06)) 
    rfd_reg_0_3_0_5_i_1
       (.I0(\m100.u0/ethc0/r_reg[rxwriteack]__0 ),
        .I1(\m100.u0/ethc0/r_reg[rxwrite] ),
        .I2(\m100.u0/ethc0/r_reg[rfcnt_n_0_][2] ),
        .O(\m100.u0/rxwrite ));
endmodule
