module fm_3d_core
   (clk_i,
    rst_i,
    int_o,
    s_wb_stb_i,
    s_wb_we_i,
    s_wb_adr_i,
    s_wb_ack_o,
    s_wb_sel_i,
    s_wb_dat_i,
    s_wb_dat_o,
    m_wb_stb_o,
    m_wb_we_o,
    m_wb_adr_o,
    m_wb_ack_i,
    m_wb_sel_o,
    m_wb_dat_o,
    backdoor,
    m_wb_dat_i);
  output backdoor;
  input clk_i;
  input rst_i;
  output int_o;
  input s_wb_stb_i;
  input s_wb_we_i;
  input [7:2]s_wb_adr_i;
  output s_wb_ack_o;
  input [3:0]s_wb_sel_i;
  input [31:0]s_wb_dat_i;
  output [31:0]s_wb_dat_o;
  output m_wb_stb_o;
  output m_wb_we_o;
  output [31:2]m_wb_adr_o;
  input m_wb_ack_i;
  output [3:0]m_wb_sel_o;
  output [31:0]m_wb_dat_o;
  input [31:0]m_wb_dat_i;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire FSM_onehot_r_state;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[2]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[3]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[4]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[5]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[5]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[5]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[5]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[5]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[5]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[5]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[5]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[6]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[6]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[6]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]FSM_onehot_r_state_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state_reg[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state_reg[5]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_onehot_r_state_reg[5]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire FSM_sequential_r_state;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_state[0]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_state[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_state[1]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_state[1]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_state[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_state[2]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_state[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_state[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_state[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_r_state[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire FSM_sequential_r_state_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire GND_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire VCC_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__0_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__0_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__0_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__0_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__0_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__0_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__0_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__0_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__0_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__0_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__1_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__1_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__1_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__1_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__1_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__1_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__1_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__1_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry__1_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_10__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_10__10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_10__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_10__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_10__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_10__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_10__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_10__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_10__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_10__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_10__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_11__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_11__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_12__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_12__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_13__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_13__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_14__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_15__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_16__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_3__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_3__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_3__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_3__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_3__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_3__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_3__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_3__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_3__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_4__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_4__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_4__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_4__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_4__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_4__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_4__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_4__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_4__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_5__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_5__10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_5__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_5__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_5__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_5__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_5__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_5__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_5__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_5__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_5__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_6__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_6__10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_6__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_6__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_6__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_6__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_6__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_6__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_6__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_6__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_6__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_7__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_7__10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_7__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_7__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_7__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_7__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_7__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_7__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_7__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_7__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_7__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_8__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_8__10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_8__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_8__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_8__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_8__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_8__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_8__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_8__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_8__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_8__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_9__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_9__10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_9__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_9__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_9__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_9__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_9__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_9__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_9__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_9__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_9__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__1_carry_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__0_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__0_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__0_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__0_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__0_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__0_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__1_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__1_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__1_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__1_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__1_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry__1_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__5_carry_i_9_n_0_repN;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__0_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__0_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__0_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__0_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__0_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__0_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__1_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__1_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__1_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry__1_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire _inferred__8__0_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk_i;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire f_multi_return_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g1_b6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire int_o;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire m_wb_ack_i;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:2]m_wb_adr_o;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[13]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[13]_INST_0_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[13]_INST_0_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[13]_INST_0_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[17]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[17]_INST_0_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[17]_INST_0_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[17]_INST_0_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[21]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[21]_INST_0_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[21]_INST_0_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[21]_INST_0_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[25]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[25]_INST_0_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[25]_INST_0_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[25]_INST_0_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[29]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[29]_INST_0_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[29]_INST_0_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[29]_INST_0_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[31]_INST_0_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[31]_INST_0_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[5]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[5]_INST_0_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[5]_INST_0_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[5]_INST_0_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[9]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[9]_INST_0_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[9]_INST_0_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \m_wb_adr_o[9]_INST_0_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]m_wb_dat_i;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:24]\^m_wb_dat_o ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]m_wb_sel_o;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire m_wb_stb_o;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire m_wb_we_o;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_adrs_m_reg_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_bc;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_bc[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_bc[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_bc[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_bc[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_bc[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_c;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_3__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_3__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_3__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_3__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_3__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_3__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_3__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_3__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_3__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_3__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_3__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_3__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_3__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_3__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_3__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_10__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_10__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_10__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_10__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_10__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_10__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_10__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_10__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_11__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_11__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_11__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_11__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_11__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_11__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_11__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_11__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_12__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_12__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_12__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_12__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_12__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_12__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_12__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_12__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_3__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_3__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_3__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_3__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_3__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_4__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_4__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_4__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_4__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_4__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_4__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_5__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_5__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_5__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_5__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_5__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_5__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_6__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_6__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_6__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_6__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_6__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_6__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_6__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_6__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_7__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_7__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_7__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_7__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_7__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_7__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_7__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_7__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_7__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_8__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_8__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_8__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_8__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_8__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_8__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_8__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_8__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_8__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_9__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_9__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_9__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_9__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_9__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_9__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_9__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_9__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[14]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[17]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[17]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[17]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[17]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[17]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[17]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[17]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[18]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[18]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_3__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_3__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_3__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_3__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_4__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_4__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_4__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_4__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_4__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_5__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_5__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_5__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_5__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_5__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_6__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_6__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_6__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_6__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_6__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_6__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_6__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_2__9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_3__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_3__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_3__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_3__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_3__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_3__9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[20]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[21]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[21]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[21]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[21]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[21]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[21]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[21]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[31]_inv_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_3__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_3__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_3__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_3__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_3__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_3__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_3__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_3__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_3__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_3__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_c[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_ccw_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_ce_tmp;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_ce_tmp_1z;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[0]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[0]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[0]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[0]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[0]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_4__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ce_tmp_1z[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_dma_size;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_dma_size[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_dma_size[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_dma_start_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_dma_start_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_dma_top_address;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_dma_top_address[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_dma_top_address[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_dma_top_address[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_dma_top_address[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_e2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_en_cull_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_err;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_err[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_exp_1z;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_exp_1z[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_f0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[14]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[14]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[14]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[14]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[14]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[14]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[14]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[14]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f0[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_f1t;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_4__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[10]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[10]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[10]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[10]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[10]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[10]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[10]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[10]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[10]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_4__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_5__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_6__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_6__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_4__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_4__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[13]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[14]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_4__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_6__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_6__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_7__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_7__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_7__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_8__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_8__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_8__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_4__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_6__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_4__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_6__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_4__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_6__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_6__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_4__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_5__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_5__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_5__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_6__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_6__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_7__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_7__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_7__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_8__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_8__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[8]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_3__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_3__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_3__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_4__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_4__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_f1t[9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_int_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_int_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_int_mask_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_int_out_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_ivw;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_ivw[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m00;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]r_m00_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[11]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[11]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[11]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[11]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[14]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[14]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[14]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[14]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[14]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[14]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[14]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[3]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[3]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[3]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[3]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[7]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[7]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[7]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[7]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[7]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[7]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m00_reg[7]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m01;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m01[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m01[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m02;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m02[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m02[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m03;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m03[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m03[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m10;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m10[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m10[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m10[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m10[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m11;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m11[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m11[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m12;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m12[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m12[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m13;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m13[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m13[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m20;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m20[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m20[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m21;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m21[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m21[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m22;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m22[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m22[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m23;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m23[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m23[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m30;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m30[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m30[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m31;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m31[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m31[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m32;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m32[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m32[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_m33;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m33[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_m33[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]r_mats_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[11]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[15]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1__3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1__3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1__3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[16]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_mats_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_pixel_color;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_pixel_top_address;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_pixel_top_address[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_pixel_top_address[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_pixel_top_address[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_rd;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[0]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[10]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[10]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[10]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[11]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[11]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[11]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[12]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[12]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[12]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[12]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[13]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[13]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[13]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[13]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[13]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[14]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[14]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[14]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[14]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[14]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[15]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[15]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[15]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[16]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[16]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[16]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[16]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[16]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[17]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[17]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[17]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[17]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[17]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[18]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[18]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[18]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[18]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[18]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[18]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[19]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[19]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[19]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[19]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[19]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[20]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[20]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[20]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[20]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[20]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[21]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[21]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[21]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[21]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[21]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[21]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[21]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[4]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[4]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[5]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[5]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[5]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[6]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[6]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[6]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[7]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[7]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[8]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[8]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[8]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[8]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[9]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[9]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[9]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd[9]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_rd_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd_reg[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd_reg[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd_reg[0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd_reg[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd_reg[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd_reg[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd_reg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd_reg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd_reg[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd_reg[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd_reg[8]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_rd_reg[8]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_req_geo_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_rstr_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_scr_h_m1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_scr_h_m1[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_scr_w;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_scr_w[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_scr_w_m1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_scr_w_m1[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_sign_1z_i_1__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_sign_1z_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_sign_1z_i_2__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_sign_1z_i_2__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_sign_1z_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_size;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]r_size_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[12]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[12]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[12]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[12]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[15]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[15]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[15]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[15]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[4]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[4]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[4]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[4]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[4]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[4]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[4]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[8]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[8]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[8]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[8]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[8]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[8]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_size_reg[8]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_state;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_state[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_state[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_state[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_state[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_state_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_state_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_state_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_sub_i_1__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_sub_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_sub_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_sub_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_sum;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[19]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[19]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[23]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[23]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[23]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]r_sum_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[15]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[15]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[15]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[19]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[19]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[19]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[3]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[3]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[3]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[7]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[7]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_sum_reg[7]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_v0_x;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[10]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[10]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[10]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[10]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[10]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[11]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[11]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[11]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[11]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[7]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x[9]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]r_v0_x_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x_reg[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x_reg[7]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x_reg[7]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_v0_x_reg[7]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_vh;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vh[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vh[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_vw;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vw[21]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vw[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vw[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_vx;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[15]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[16]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[17]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[18]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[19]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[20]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[21]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[21]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]r_vx_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[11]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[11]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[11]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[11]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[14]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[14]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[14]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[14]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[14]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[14]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[14]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[3]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[3]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[3]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[3]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[7]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[7]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[7]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vx_reg[7]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_vy;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[21]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_vy[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_vz_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_x0_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[11]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]r_x_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x_reg[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x_reg[11]_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x_reg[11]_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_x_reg[11]_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y0_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_y[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_y[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_y[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_y[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_y[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_y[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_y[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_y[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_y[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_y[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_y[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_y_flip_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_inferred__1_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_inferred__1_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_inferred__1_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_inferred__1_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_inferred__1_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_inferred__1_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_inferred__1_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_inferred__1_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_inferred__1_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_inferred__1_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_inferred__1_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result0_inferred__1_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__0_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__1_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__2_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__3_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire result3_inferred__4_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rst_i;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire s_wb_ack_o;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:2]s_wb_adr_i;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]s_wb_dat_i;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]s_wb_dat_o;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]s_wb_sel_i;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire s_wb_stb_i;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire s_wb_we_i;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[11]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[11]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[11]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[15]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[15]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[15]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[15]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[3]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[3]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[3]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[7]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[7]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[7]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[7]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd/r_mats[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m01/r_mats[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m0123/r_mats[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fadd_m23/r_mats[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fmul/r_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fmul/r_c[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fmul/r_ce_tmp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fmul/r_ce_tmp_1z[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fmul/r_ce_tmp_1z[1]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fmul/r_ce_tmp_1z[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fmul/r_ce_tmp_1z[2]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fmul/r_ce_tmp_1z[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fmul/r_ce_tmp_1z[3]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fmul/r_ce_tmp_1z[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fmul/r_ce_tmp_1z[4]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_fmul/r_ce_tmp_1z[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_frcp/frcp_rom/r_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/r_int_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/r_int_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/data0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/p_0_in0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/r_bc ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_clip/r_exp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_clip/r_exp_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_clip/r_f0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/r_sign_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/r_sub ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/r_vw_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_clip/r_vz ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_clip/u_fadd/norm/f_incdec_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_clip/u_fadd/r_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/r_sign_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/w_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_clip/u_fadd/w_exp_l ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/w_mag_frac_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/w_mag_frac_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/w_mag_frac_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/w_mag_frac_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/w_mag_frac_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/w_mag_frac_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/w_mag_frac_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_clip/u_fadd/w_sign ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [20:0]\u_geo/u_geo_clip/w_add_in_a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_clip/w_f0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_clip/w_f1t ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_clip/w_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_geo/u_geo_cull/A ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_geo/u_geo_cull/B ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return0_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/f_multi_return_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [23:0]\u_geo/u_geo_cull/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\u_geo/u_geo_cull/r_state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [23:0]\u_geo/u_geo_cull/r_sum0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/r_sum_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_cull/w_set_tri ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/r_lat_cnt ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_matrix/r_vx_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_matrix/r_vy_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_matrix/r_vz_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/r_wait_end_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/r_wait_end_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/r_wait_end_3z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/data0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fadd_m01/norm/w_c_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/u_fadd_m01/r_f0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/u_fadd_m01/r_f1t ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fadd_m01/r_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/r_sign_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/r_sign_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/r_sub ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/w_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fadd_m01/w_exp_l ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/u_fadd_m01/w_f0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/u_fadd_m01/w_f1t ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fadd_m01/w_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/w_sign ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m01/w_sub11_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/data0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fadd_m0123/norm/w_c_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fadd_m0123/r_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/r_sign_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/r_sign_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/r_sub ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/w_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fadd_m0123/w_exp_l ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fadd_m0123/w_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/w_sign ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m0123/w_sub11_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/data0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fadd_m23/norm/w_c_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/u_fadd_m23/r_f0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/u_fadd_m23/r_f1t ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fadd_m23/r_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/r_sign_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/r_sign_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/r_sub ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/w_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fadd_m23/w_exp_l ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/u_fadd_m23/w_f0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/u_fadd_m23/w_f1t ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fadd_m23/w_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/w_sign ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fadd_m23/w_sub11_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fmul_m0/norm/w_c_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [17:0]\u_geo/u_geo_matrix/u_fmul_m0/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[15]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[15]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[15]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[16]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[16]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[16]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_sign_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/r_sign_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_adder_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m0/w_sign ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fmul_m1/norm/w_c_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [17:0]\u_geo/u_geo_matrix/u_fmul_m1/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[15]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[15]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[15]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[16]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[16]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[16]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_sign_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/r_sign_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_adder_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m1/w_sign ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fmul_m2/norm/w_c_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [17:0]\u_geo/u_geo_matrix/u_fmul_m2/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[15]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[15]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[15]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[16]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[16]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[16]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_sign_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/r_sign_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_adder_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m2/w_sign ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fmul_m3/norm/w_c_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [17:0]\u_geo/u_geo_matrix/u_fmul_m3/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[15]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[15]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[15]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[16]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[16]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[16]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_sign_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/r_sign_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_matrix/w_add0123_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_matrix/w_add01_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_matrix/w_add23_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_matrix/w_m0_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_matrix/w_m1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_matrix/w_m2_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_matrix/w_m3_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/w_vx_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/w_vy_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_matrix/w_vz_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_matrix/w_wait_end ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [29:0]\u_geo/u_geo_mem/r_cur_adrs ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\u_geo/u_geo_mem/r_cur_adrs_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[29]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[29]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[29]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[29]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:1]\u_geo/u_geo_mem/r_size ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_mem/r_size__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_vx ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_vy ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/r_vz ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [20:15]\u_geo/u_geo_mem/w_f22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_mem/w_read_end ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [17:0]\u_geo/u_geo_persdiv/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_persdiv/r_ce_tmp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_persdiv/r_ce_tmp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_persdiv/r_ce_tmp_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_persdiv/r_ivw ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/r_sign_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]\u_geo/u_geo_persdiv/r_state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_persdiv/u_fmul/norm/w_c_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[15]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[15]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[15]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[16]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[16]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[16]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/r_sign_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_adder_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_fmul/w_sign ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[31]_inv_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_a_sign ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_persdiv/u_frcp/w_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_persdiv/w_b_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_persdiv/w_cf_tmp2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_persdiv/w_fmul_a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]\u_geo/u_geo_persdiv/w_rom_base ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_tri/exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_tri/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_tri/p_0_in0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_geo/u_geo_tri/p_0_in__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_tri/r_v0_outcode ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_tri/r_v1_outcode ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_tri/r_v2_outcode ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_tri/r_vy ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [12:12]\u_geo/u_geo_tri/u_ftoi/f_ftoi__60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_tri/w_set_v0_x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_tri/w_set_v0_y ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_tri/w_set_v1_x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_tri/w_set_v1_y ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_tri/w_set_v2_x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_tri/w_set_v2_y ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_tri/w_set_y ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_tri/w_tri_outside ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [12:1]\u_geo/u_geo_tri/w_ui_2c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [17:0]\u_geo/u_geo_viewport/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_viewport/r_ce_tmp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_viewport/r_ce_tmp_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_viewport/r_exp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_viewport/r_exp_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_viewport/r_f0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/r_sign_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\u_geo/u_geo_viewport/r_state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/r_sub ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_viewport/sel0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_viewport/u_fadd/norm/w_c_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_viewport/u_fadd/r_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/r_sign_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_viewport/u_fadd/w_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\u_geo/u_geo_viewport/u_fadd/w_exp_l ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fadd/w_mag__7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_viewport/u_fmul/norm/w_c_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_ce_tmp_1z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[15]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[15]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[15]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[16]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[16]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[16]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_sign_1z_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/r_sign_2z ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_adder_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/u_fmul/w_sign ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\u_geo/u_geo_viewport/w_a_exp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_viewport/w_cf_tmp2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/w_f0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_viewport/w_f1t ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/u_geo_viewport/w_fadd_a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/w_fadd_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\u_geo/u_geo_viewport/w_fmul_b ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [16:0]\u_geo/u_geo_viewport/w_mats ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/u_geo_viewport/w_set_vy ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/w_dma_end ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/w_en_clip ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/w_en_dma ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/w_en_mvp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/w_en_tri ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/w_en_view ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/w_outcode_clip ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/w_outcode_pdiv ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:0]\u_geo/w_outcode_view ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/w_state_clip ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/w_state_cull ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/w_state_if ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/w_state_mat ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/w_state_pd ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_geo/w_state_view ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_geo/w_v0_x_tri ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_geo/w_v0_y_tri ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_geo/w_v1_x_tri ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_geo/w_v1_y_tri ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_geo/w_v2_x_tri ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_geo/w_v2_y_tri ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vw_clip ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vw_mvp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vx_clip ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vx_dma ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vx_mvp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vx_pdiv ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vx_view ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vy_clip ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vy_dma ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vy_mvp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vy_pdiv ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vy_view ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vz_dma ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]\u_geo/w_vz_mvp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_mem_arb/r_req_geo ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_mem_arb/r_state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_mem_arb/w_pri__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_ras/B ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:0]\u_ras/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:0]\u_ras/p_2_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/p_2_in[7]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:1]\u_ras/r_e2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:0]\u_ras/r_err ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:0]\u_ras/r_y ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__1_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__1_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__1_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__1_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__5_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__8__0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__8__0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__8__0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__8__0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__8__0_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__8__0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__8__0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__8__0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/_inferred__8__0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_e2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_state_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_state_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_ras/u_ras_line/r_x0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_ras/u_ras_line/r_x1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_x_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_x_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_x_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_x_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_x_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_x_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_x_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_x_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_x_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_x_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_x_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_ras/u_ras_line/r_y0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/r_y1_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_inferred__1_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_inferred__1_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_inferred__1_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/result0_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dx ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym__22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_dym_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_end00_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_end0__3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_end0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_end0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_end0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_end0_inferred__0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_end0_inferred__0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_end0_inferred__0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_err__0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_err__0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_err__0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_err__0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_err__0_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_err__0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_err__0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_err__0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_err__0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject0__7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject1__7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject1_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject1_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject1_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_reject__2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sx_flag1__5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sx_flag1_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sx_flag1_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sx_flag1_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sx_flag1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sx_flag1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sx_flag1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sx_flag1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sy_flag1__5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sy_flag1_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sy_flag1_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sy_flag1_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sy_flag1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sy_flag1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sy_flag1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_line/w_sy_flag1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[25]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[25]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[25]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_adrs_m_reg_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/r_state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\u_ras/u_ras_mem/r_x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_mem/w_y0_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/FSM_sequential_r_state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/FSM_sequential_r_state[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/f_reject0_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/f_reject1_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/f_reject_return ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/p_0_in0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/p_1_in10_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/p_1_in1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/p_1_in8_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\u_ras/u_ras_state/r_state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_state[0]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_state[0]_repN_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_state[0]_repN_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_state[0]_repN_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_state[0]_repN_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_state[1]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_state[1]_repN_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_state[1]_repN_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_state[1]_repN_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_x_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_x_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_x_reg_n_0_[10]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_x_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_x_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_x_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_x_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_x_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_x_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_x_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_x_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_x_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_[10]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_[1]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v0_y_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_x_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_x_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_x_reg_n_0_[10]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_x_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_x_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_x_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_x_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_x_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_x_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_x_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_x_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_x_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[0]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[1]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[5]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[6]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[7]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[8]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v1_y_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_x_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_x_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_x_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_x_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_x_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_x_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_x_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_x_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_x_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_x_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_x_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_y_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_y_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_y_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_y_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_y_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_y_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_y_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_y_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_y_reg_n_0_[6]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_y_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_y_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/r_v2_y_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result115_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result121_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result132_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result141_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result14_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result17_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result316_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result324_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result327_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result333_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result336_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3__7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__1_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__1_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__1_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__2_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__2_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__2_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__2_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__2_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__2_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__2_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__3_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__3_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__3_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__3_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__3_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__3_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__3_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__4_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__4_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__4_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__4_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__4_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__4_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/result3_inferred__4_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/u_ras_state/w_set_vtx ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/w_ack_pix ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_ras/w_dy ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:1]\u_ras/w_e2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/w_en_pix ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:0]\u_ras/w_err ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_ras/w_v0_x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/w_v0_x[10]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_ras/w_v0_y ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/w_v0_y[10]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_ras/w_v1_x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_ras/w_v1_y ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/w_x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:1]\u_ras/w_x0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_ras/w_x1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/w_y ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:1]\u_ras/w_y0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\u_ras/w_y1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/w_y1[1]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras/w_y1[6]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_state[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_x0_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_line/r_y0_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_mem/r_x ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_ras_mem/r_x[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_sys/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [8:0]\u_sys/p_21_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_sys/r_pixel_color ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_sys/r_rstr ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [20:15]\u_sys/w_f22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_sys/w_hit1A_w__2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u_sys/w_int_set ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:7]\u_sys/w_rd ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_ack;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:2]w_adrs_geo;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:2]w_adrs_ras;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_ccw;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_1__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_1__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_2__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_2__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_3__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_3__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_4__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_10__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_10__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_10__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_10__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_11__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_11__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_11__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_11__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_12__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_12__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_12__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_12__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_13__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_13__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_13__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_13__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_14__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_14__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_14__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_14__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_15__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_15__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_15__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_15__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_16__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_16__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_16__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_16__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_1__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_1__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_1__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_2__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_2__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_2__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_33__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_33__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_33__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_34__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_34__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_34__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_35__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_35__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_35__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_36__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_36__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_36__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_37__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_37__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_37__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_38__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_38__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_38__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_39__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_39__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_39__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_3__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_3__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_3__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_40__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_40__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_40__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_41__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_41__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_41__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_42__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_42__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_42__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_43__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_43__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_43__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_44__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_44__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_44__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_45__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_45__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_45__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_46__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_46__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_46__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_47__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_47__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_47__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_47_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_48__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_48__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_48__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_48_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_49_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_4__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_4__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_4__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_50_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_51_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_52_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_53_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_54_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_55_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_56_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_57_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_58_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_59_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_5__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_5__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_5__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_5__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_60_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_61_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_62_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_6__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_6__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_6__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_6__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_7__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_7__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_7__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_7__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_8__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_8__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_8__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_8__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_9__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_9__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_9__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_9__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_cf_tmp_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]w_dma_size;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_dma_start;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [29:0]w_dma_top_address;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_dym_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_dym_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_dym_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_dym_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_dym_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_dym_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_dym_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_dym_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_dym_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_dym_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_dym_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_en;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_en_cull;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_end0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_end0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_end0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_end0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_end0_inferred__0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_end0_inferred__0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_end0_inferred__0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_end0_inferred__0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__0_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__1_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__1_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__1_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__1_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__1_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__1_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry__1_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_err__0_carry_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m00;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m01;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m02;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m03;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m10;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m11;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m12;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m13;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m20;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m21;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m22;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m23;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m30;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m31;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m32;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_m33;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_1__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_1__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_1__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_1__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_1__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_1__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_2__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_2__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_2__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_2__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_2__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_2__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_3__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_3__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_3__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_3__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_3__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_3__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_4__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_4__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_4__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_4__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_4__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_4__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_5__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_5__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_5__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_5__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_5__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_5__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_5__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_6__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_6__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_6__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_6__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_6__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_6__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_6__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_7__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_7__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_7__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_7__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_7__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_7__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_7__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_8__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_8__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_8__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_8__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_8__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_8__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_8__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_mag_frac_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [29:0]w_pixel_top_address;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject0_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_reject1_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_req_geo;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_rom_correct_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]w_scr_h_m1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]w_scr_w;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]w_scr_w_m1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry__0_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry__0_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sx_flag1_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry__0_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry__0_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_sy_flag1_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]w_v0_x;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]w_v0_y;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]w_v1_x;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]w_v1_y;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]w_v2_x;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]w_v2_y;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_vh;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [21:0]w_vw;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y0_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y0_carry_i_1__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y0_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y0_carry_i_2__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y0_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y0_carry_i_3__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y0_carry_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y0_carry_i_4__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_y_flip;

  assign backdoor =  w_y_flip ;

  assign m_wb_dat_o[31:24] = \^m_wb_dat_o [31:24];
  assign m_wb_dat_o[23:16] = \^m_wb_dat_o [31:24];
  assign m_wb_dat_o[15:8] = \^m_wb_dat_o [31:24];
  assign m_wb_dat_o[7:0] = \^m_wb_dat_o [31:24];
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \FSM_onehot_r_state[0]_i_1 
       (.I0(w_dma_start),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\u_geo/w_en_dma ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\FSM_onehot_r_state[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000010111000)) 
    \FSM_onehot_r_state[0]_i_1__0 
       (.I0(\u_geo/u_geo_tri/w_set_v0_y ),
        .I1(\u_geo/u_geo_tri/w_set_v1_y ),
        .I2(\u_geo/u_geo_tri/w_tri_outside ),
        .I3(\u_geo/u_geo_tri/w_set_v2_y ),
        .I4(\u_geo/w_en_tri ),
        .I5(\FSM_onehot_r_state[6]_i_6_n_0 ),
        .O(FSM_onehot_r_state));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00000100)) 
    \FSM_onehot_r_state[1]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I3(\u_geo/w_en_dma ),
        .I4(\u_geo/u_geo_mem/w_read_end ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .O(\FSM_onehot_r_state[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_onehot_r_state[2]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .O(\FSM_onehot_r_state[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_onehot_r_state[2]_i_1__0 
       (.I0(\u_geo/u_geo_tri/w_set_v0_y ),
        .I1(\u_geo/w_state_if ),
        .O(\FSM_onehot_r_state[2]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \FSM_onehot_r_state[3]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .O(\FSM_onehot_r_state[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \FSM_onehot_r_state[3]_i_1__0 
       (.I0(\u_geo/u_geo_tri/w_set_v0_y ),
        .I1(\u_geo/u_geo_tri/p_0_in0_in ),
        .I2(\u_geo/w_state_if ),
        .O(\FSM_onehot_r_state[3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \FSM_onehot_r_state[4]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .O(\FSM_onehot_r_state[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \FSM_onehot_r_state[4]_i_1__0 
       (.I0(\u_geo/u_geo_tri/w_set_v0_y ),
        .I1(\u_geo/u_geo_tri/w_set_v1_y ),
        .I2(\u_geo/u_geo_tri/p_0_in0_in ),
        .I3(\u_geo/w_state_if ),
        .O(\FSM_onehot_r_state[4]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFAEAEAE)) 
    \FSM_onehot_r_state[5]_i_1 
       (.I0(\r_size[15]_i_1_n_0 ),
        .I1(\u_geo/w_dma_end ),
        .I2(w_dma_start),
        .I3(\u_geo/w_en_dma ),
        .I4(\u_geo/w_state_mat ),
        .O(\FSM_onehot_r_state[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_onehot_r_state[5]_i_10 
       (.I0(\u_geo/u_geo_mem/r_size__0 [3]),
        .I1(w_dma_size[3]),
        .I2(w_dma_size[5]),
        .I3(\u_geo/u_geo_mem/r_size__0 [5]),
        .I4(w_dma_size[4]),
        .I5(\u_geo/u_geo_mem/r_size__0 [4]),
        .O(\FSM_onehot_r_state[5]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_onehot_r_state[5]_i_11 
       (.I0(\u_geo/u_geo_mem/r_size__0 [0]),
        .I1(w_dma_size[0]),
        .I2(w_dma_size[2]),
        .I3(\u_geo/u_geo_mem/r_size__0 [2]),
        .I4(w_dma_size[1]),
        .I5(\u_geo/u_geo_mem/r_size__0 [1]),
        .O(\FSM_onehot_r_state[5]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \FSM_onehot_r_state[5]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I2(\FSM_onehot_r_state[5]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .I5(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[4] ),
        .O(\FSM_onehot_r_state[5]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \FSM_onehot_r_state[5]_i_1__1 
       (.I0(\u_geo/u_geo_tri/w_set_v0_y ),
        .I1(\u_geo/u_geo_tri/w_set_v1_y ),
        .I2(\u_geo/u_geo_tri/p_0_in ),
        .I3(\u_geo/u_geo_tri/p_0_in0_in ),
        .I4(\u_geo/w_state_if ),
        .O(\FSM_onehot_r_state[5]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00004540)) 
    \FSM_onehot_r_state[5]_i_2 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(\u_geo/u_geo_mem/w_read_end ),
        .I2(\u_geo/w_en_dma ),
        .I3(w_dma_start),
        .I4(\FSM_onehot_r_state[5]_i_4_n_0 ),
        .O(\FSM_onehot_r_state[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    \FSM_onehot_r_state[5]_i_2__0 
       (.I0(\u_geo/w_en_dma ),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/w_state_clip ),
        .I3(\u_geo/w_en_mvp ),
        .O(\FSM_onehot_r_state[5]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \FSM_onehot_r_state[5]_i_4 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\FSM_onehot_r_state[5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \FSM_onehot_r_state[5]_i_6 
       (.I0(w_dma_size[15]),
        .I1(\u_geo/u_geo_mem/r_size__0 [15]),
        .O(\FSM_onehot_r_state[5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_onehot_r_state[5]_i_7 
       (.I0(\u_geo/u_geo_mem/r_size__0 [12]),
        .I1(w_dma_size[12]),
        .I2(w_dma_size[14]),
        .I3(\u_geo/u_geo_mem/r_size__0 [14]),
        .I4(w_dma_size[13]),
        .I5(\u_geo/u_geo_mem/r_size__0 [13]),
        .O(\FSM_onehot_r_state[5]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_onehot_r_state[5]_i_8 
       (.I0(\u_geo/u_geo_mem/r_size__0 [9]),
        .I1(w_dma_size[9]),
        .I2(w_dma_size[11]),
        .I3(\u_geo/u_geo_mem/r_size__0 [11]),
        .I4(w_dma_size[10]),
        .I5(\u_geo/u_geo_mem/r_size__0 [10]),
        .O(\FSM_onehot_r_state[5]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \FSM_onehot_r_state[5]_i_9 
       (.I0(\u_geo/u_geo_mem/r_size__0 [6]),
        .I1(w_dma_size[6]),
        .I2(w_dma_size[8]),
        .I3(\u_geo/u_geo_mem/r_size__0 [8]),
        .I4(w_dma_size[7]),
        .I5(\u_geo/u_geo_mem/r_size__0 [7]),
        .O(\FSM_onehot_r_state[5]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \FSM_onehot_r_state[6]_i_1 
       (.I0(\u_geo/w_en_tri ),
        .I1(\u_geo/w_state_cull ),
        .I2(\FSM_onehot_r_state[6]_i_4_n_0 ),
        .I3(\u_geo/u_geo_tri/w_set_v2_y ),
        .I4(\u_geo/w_en_view ),
        .I5(\FSM_onehot_r_state[6]_i_6_n_0 ),
        .O(\FSM_onehot_r_state[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \FSM_onehot_r_state[6]_i_10 
       (.I0(\u_geo/u_geo_tri/r_v1_outcode [4]),
        .I1(\u_geo/u_geo_tri/r_v1_outcode [5]),
        .I2(\u_geo/u_geo_tri/r_v2_outcode [4]),
        .I3(\u_geo/u_geo_tri/r_v2_outcode [5]),
        .I4(\u_geo/u_geo_tri/r_v0_outcode [5]),
        .I5(\u_geo/u_geo_tri/r_v0_outcode [4]),
        .O(\FSM_onehot_r_state[6]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \FSM_onehot_r_state[6]_i_2 
       (.I0(\FSM_onehot_r_state[6]_i_4_n_0 ),
        .I1(\u_geo/u_geo_tri/w_set_v2_y ),
        .I2(\u_geo/u_geo_tri/w_tri_outside ),
        .I3(\u_geo/u_geo_tri/p_0_in ),
        .I4(\u_geo/w_state_if ),
        .I5(\u_geo/u_geo_tri/p_0_in0_in ),
        .O(\FSM_onehot_r_state[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_onehot_r_state[6]_i_3 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_state [1]),
        .O(\u_geo/w_state_cull ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_onehot_r_state[6]_i_4 
       (.I0(\u_geo/u_geo_tri/w_set_v0_y ),
        .I1(\u_geo/u_geo_tri/w_set_v1_y ),
        .O(\FSM_onehot_r_state[6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0100)) 
    \FSM_onehot_r_state[6]_i_5 
       (.I0(\u_geo/u_geo_viewport/r_state [0]),
        .I1(\u_geo/u_geo_viewport/r_state [1]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .O(\u_geo/w_en_view ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \FSM_onehot_r_state[6]_i_6 
       (.I0(\u_geo/u_geo_tri/p_0_in0_in ),
        .I1(\u_geo/w_state_if ),
        .I2(\u_geo/u_geo_tri/p_0_in ),
        .O(\FSM_onehot_r_state[6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \FSM_onehot_r_state[6]_i_7 
       (.I0(\FSM_onehot_r_state[6]_i_8_n_0 ),
        .I1(\FSM_onehot_r_state[6]_i_9_n_0 ),
        .I2(\FSM_onehot_r_state[6]_i_10_n_0 ),
        .O(\u_geo/u_geo_tri/w_tri_outside ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF80808080808080)) 
    \FSM_onehot_r_state[6]_i_8 
       (.I0(\u_geo/u_geo_tri/r_v0_outcode [2]),
        .I1(\u_geo/u_geo_tri/r_v2_outcode [2]),
        .I2(\u_geo/u_geo_tri/r_v1_outcode [2]),
        .I3(\u_geo/u_geo_tri/r_v0_outcode [3]),
        .I4(\u_geo/u_geo_tri/r_v2_outcode [3]),
        .I5(\u_geo/u_geo_tri/r_v1_outcode [3]),
        .O(\FSM_onehot_r_state[6]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF80808080808080)) 
    \FSM_onehot_r_state[6]_i_9 
       (.I0(\u_geo/u_geo_tri/r_v0_outcode [0]),
        .I1(\u_geo/u_geo_tri/r_v2_outcode [0]),
        .I2(\u_geo/u_geo_tri/r_v1_outcode [0]),
        .I3(\u_geo/u_geo_tri/r_v0_outcode [1]),
        .I4(\u_geo/u_geo_tri/r_v2_outcode [1]),
        .I5(\u_geo/u_geo_tri/r_v1_outcode [1]),
        .O(\FSM_onehot_r_state[6]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \FSM_onehot_r_state[9]_i_1 
       (.I0(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[7] ),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(\FSM_onehot_r_state[9]_i_2_n_0 ),
        .I5(\FSM_onehot_r_state[9]_i_3_n_0 ),
        .O(\FSM_onehot_r_state[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8888888F88888888)) 
    \FSM_onehot_r_state[9]_i_2 
       (.I0(\u_geo/w_en_mvp ),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .I5(\u_geo/w_en_clip ),
        .O(\FSM_onehot_r_state[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \FSM_onehot_r_state[9]_i_3 
       (.I0(\u_geo/u_geo_clip/r_bc ),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[8] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .O(\FSM_onehot_r_state[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_onehot_r_state_reg[5]_i_3 
       (.CI(FSM_onehot_r_state_reg[3]),
        .CO({\FSM_onehot_r_state_reg[5]_i_3_n_0 ,\FSM_onehot_r_state_reg[5]_i_3_n_1 ,\u_geo/u_geo_mem/w_read_end ,\FSM_onehot_r_state_reg[5]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\FSM_onehot_r_state[5]_i_6_n_0 ,\FSM_onehot_r_state[5]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_onehot_r_state_reg[5]_i_5 
       (.CI(\<const0>__0__0 ),
        .CO(FSM_onehot_r_state_reg),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\FSM_onehot_r_state[5]_i_8_n_0 ,\FSM_onehot_r_state[5]_i_9_n_0 ,\FSM_onehot_r_state[5]_i_10_n_0 ,\FSM_onehot_r_state[5]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44FF00FC)) 
    \FSM_sequential_r_state[0]_i_1 
       (.I0(\u_geo/w_state_view ),
        .I1(\u_geo/u_geo_persdiv/r_state [2]),
        .I2(\u_geo/w_en_clip ),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [1]),
        .O(\FSM_sequential_r_state[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_r_state[0]_i_1__0 
       (.I0(\u_geo/u_geo_viewport/r_state [0]),
        .I1(\u_geo/u_geo_viewport/r_state [3]),
        .O(FSM_sequential_r_state));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \FSM_sequential_r_state[0]_i_1__1 
       (.I0(\u_ras/u_ras_state/r_state [0]),
        .I1(\u_ras/u_ras_state/FSM_sequential_r_state ),
        .O(\FSM_sequential_r_state[0]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4FF0)) 
    \FSM_sequential_r_state[1]_i_1 
       (.I0(\u_geo/w_state_view ),
        .I1(\u_geo/u_geo_persdiv/r_state [2]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .O(\FSM_sequential_r_state[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \FSM_sequential_r_state[1]_i_10 
       (.I0(\u_ras/u_ras_state/p_1_in8_in ),
        .I1(\u_ras/u_ras_state/p_1_in ),
        .I2(\u_ras/u_ras_state/p_1_in10_in ),
        .I3(\u_ras/u_ras_state/p_1_in1_in ),
        .I4(\u_ras/u_ras_state/result121_out ),
        .I5(\u_ras/u_ras_state/result115_out ),
        .O(\u_ras/u_ras_state/f_reject0_return ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h08888808)) 
    \FSM_sequential_r_state[1]_i_11 
       (.I0(\u_geo/u_geo_cull/r_state [1]),
        .I1(\u_geo/u_geo_cull/r_state [0]),
        .I2(w_en_cull),
        .I3(w_ccw),
        .I4(\u_geo/u_geo_cull/p_0_in ),
        .O(w_en));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0400)) 
    \FSM_sequential_r_state[1]_i_12 
       (.I0(\u_ras/u_ras_state/p_1_in10_in ),
        .I1(\u_ras/u_ras_state/result333_in ),
        .I2(\u_ras/u_ras_state/p_1_in1_in ),
        .I3(\u_ras/u_ras_state/result316_in ),
        .O(\u_ras/u_ras_state/result121_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0400)) 
    \FSM_sequential_r_state[1]_i_13 
       (.I0(\u_ras/u_ras_state/p_1_in8_in ),
        .I1(\u_ras/u_ras_state/result324_in ),
        .I2(\u_ras/u_ras_state/p_1_in ),
        .I3(\u_ras/u_ras_state/result3__7 ),
        .O(\u_ras/u_ras_state/result115_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \FSM_sequential_r_state[1]_i_1__0 
       (.I0(\u_ras/u_ras_state/r_state [0]),
        .I1(\u_ras/u_ras_state/r_state [1]),
        .I2(\u_ras/u_ras_state/FSM_sequential_r_state ),
        .O(\FSM_sequential_r_state[1]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h06)) 
    \FSM_sequential_r_state[1]_i_1__1 
       (.I0(\u_geo/u_geo_viewport/r_state [1]),
        .I1(\u_geo/u_geo_viewport/r_state [0]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .O(\FSM_sequential_r_state[1]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \FSM_sequential_r_state[1]_i_3 
       (.I0(\u_ras/u_ras_state/p_1_in ),
        .I1(\u_ras/u_ras_state/p_0_in ),
        .I2(\u_ras/u_ras_state/p_1_in1_in ),
        .I3(\u_ras/u_ras_state/p_0_in0_in ),
        .I4(\u_ras/u_ras_state/result17_out ),
        .I5(\u_ras/u_ras_state/result14_out ),
        .O(\u_ras/u_ras_state/f_reject1_return ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \FSM_sequential_r_state[1]_i_4 
       (.I0(\u_ras/u_ras_state/p_0_in ),
        .I1(\u_ras/u_ras_state/p_1_in8_in ),
        .I2(\u_ras/u_ras_state/p_0_in0_in ),
        .I3(\u_ras/u_ras_state/p_1_in10_in ),
        .I4(\u_ras/u_ras_state/result141_out ),
        .I5(\u_ras/u_ras_state/result132_out ),
        .O(\u_ras/u_ras_state/f_reject_return ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0400)) 
    \FSM_sequential_r_state[1]_i_6 
       (.I0(\u_ras/u_ras_state/p_1_in1_in ),
        .I1(\u_ras/u_ras_state/result316_in ),
        .I2(\u_ras/u_ras_state/p_0_in0_in ),
        .I3(\u_ras/u_ras_state/result336_in ),
        .O(\u_ras/u_ras_state/result17_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0400)) 
    \FSM_sequential_r_state[1]_i_7 
       (.I0(\u_ras/u_ras_state/p_1_in ),
        .I1(\u_ras/u_ras_state/result3__7 ),
        .I2(\u_ras/u_ras_state/p_0_in ),
        .I3(\u_ras/u_ras_state/result327_in ),
        .O(\u_ras/u_ras_state/result14_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0400)) 
    \FSM_sequential_r_state[1]_i_8 
       (.I0(\u_ras/u_ras_state/p_0_in0_in ),
        .I1(\u_ras/u_ras_state/result336_in ),
        .I2(\u_ras/u_ras_state/p_1_in10_in ),
        .I3(\u_ras/u_ras_state/result333_in ),
        .O(\u_ras/u_ras_state/result141_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0400)) 
    \FSM_sequential_r_state[1]_i_9 
       (.I0(\u_ras/u_ras_state/p_0_in ),
        .I1(\u_ras/u_ras_state/result327_in ),
        .I2(\u_ras/u_ras_state/p_1_in8_in ),
        .I3(\u_ras/u_ras_state/result324_in ),
        .O(\u_ras/u_ras_state/result132_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7CCC)) 
    \FSM_sequential_r_state[2]_i_1 
       (.I0(\u_geo/w_state_view ),
        .I1(\u_geo/u_geo_persdiv/r_state [2]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .O(\FSM_sequential_r_state[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h006A)) 
    \FSM_sequential_r_state[2]_i_1__0 
       (.I0(\u_geo/u_geo_viewport/r_state [2]),
        .I1(\u_geo/u_geo_viewport/r_state [0]),
        .I2(\u_geo/u_geo_viewport/r_state [1]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .O(\FSM_sequential_r_state[2]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2000)) 
    \FSM_sequential_r_state[3]_i_2 
       (.I0(\u_geo/u_geo_viewport/r_state [2]),
        .I1(\u_geo/u_geo_viewport/r_state [3]),
        .I2(\u_geo/u_geo_viewport/r_state [0]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .O(\FSM_sequential_r_state[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF80)) 
    \FSM_sequential_r_state[3]_i_3 
       (.I0(\u_geo/u_geo_persdiv/r_state [0]),
        .I1(\u_geo/u_geo_persdiv/r_state [2]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_viewport/r_state [2]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/u_geo_viewport/r_state [1]),
        .O(\FSM_sequential_r_state[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000011111110)) 
    \FSM_sequential_r_state[3]_i_4 
       (.I0(\u_geo/u_geo_viewport/r_state [0]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_tri/p_0_in0_in ),
        .I3(\u_geo/u_geo_tri/p_0_in ),
        .I4(\u_geo/w_state_if ),
        .I5(\u_geo/u_geo_viewport/r_state [1]),
        .O(\FSM_sequential_r_state[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \FSM_sequential_r_state_reg[3]_i_1 
       (.I0(\FSM_sequential_r_state[3]_i_3_n_0 ),
        .I1(\FSM_sequential_r_state[3]_i_4_n_0 ),
        .O(FSM_sequential_r_state_reg),
        .S(\u_geo/u_geo_viewport/r_state [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_1
       (.G(GND_2));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_1
       (.P(VCC_2));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__1_carry__0_i_1
       (.I0(\u_ras/u_ras_line/r_y0 [7]),
        .I1(_inferred__1_carry_i_9__9_n_0),
        .I2(\u_ras/u_ras_line/r_y1_reg_n_0_[7] ),
        .I3(_inferred__1_carry__0_i_9_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_1_in [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__1_carry__0_i_10
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[6] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[6] ),
        .I5(\u_ras/u_ras_state/r_v1_y_reg_n_0_[6] ),
        .O(_inferred__1_carry__0_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__1_carry__0_i_11
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[5] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[5] ),
        .I5(\u_ras/u_ras_state/r_v1_y_reg_n_0_[5] ),
        .O(_inferred__1_carry__0_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__1_carry__0_i_12
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[4] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[4] ),
        .I5(\u_ras/u_ras_state/r_v1_y_reg_n_0_[4] ),
        .O(_inferred__1_carry__0_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    _inferred__1_carry__0_i_13
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_v0_y_reg_n_0_[7] ),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[7] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[7] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__1_carry__0_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    _inferred__1_carry__0_i_14
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_v0_y_reg_n_0_[6] ),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[6] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[6] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__1_carry__0_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    _inferred__1_carry__0_i_15
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_v0_y_reg_n_0_[5] ),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[5] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[5] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__1_carry__0_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    _inferred__1_carry__0_i_16
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_v0_y_reg_n_0_[4] ),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[4] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[4] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__1_carry__0_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__1_carry__0_i_2
       (.I0(\u_ras/u_ras_line/r_y0 [6]),
        .I1(_inferred__1_carry_i_9__9_n_0),
        .I2(\u_ras/u_ras_line/r_y1_reg_n_0_[6] ),
        .I3(_inferred__1_carry__0_i_10_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_1_in [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__1_carry__0_i_3
       (.I0(\u_ras/u_ras_line/r_y0 [5]),
        .I1(_inferred__1_carry_i_9__9_n_0),
        .I2(\u_ras/u_ras_line/r_y1_reg_n_0_[5] ),
        .I3(_inferred__1_carry__0_i_11_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_1_in [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__1_carry__0_i_4
       (.I0(\u_ras/u_ras_line/r_y0 [4]),
        .I1(_inferred__1_carry_i_9__9_n_0),
        .I2(\u_ras/u_ras_line/r_y1_reg_n_0_[4] ),
        .I3(_inferred__1_carry__0_i_12_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_1_in [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDE1212DE)) 
    _inferred__1_carry__0_i_5
       (.I0(_inferred__1_carry__0_i_9_n_0),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(_inferred__1_carry__0_i_13_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [7]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[7] ),
        .O(_inferred__1_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDE1212DE)) 
    _inferred__1_carry__0_i_6
       (.I0(_inferred__1_carry__0_i_10_n_0),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(_inferred__1_carry__0_i_14_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [6]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[6] ),
        .O(_inferred__1_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDE1212DE)) 
    _inferred__1_carry__0_i_7
       (.I0(_inferred__1_carry__0_i_11_n_0),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(_inferred__1_carry__0_i_15_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [5]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[5] ),
        .O(_inferred__1_carry__0_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDE1212DE)) 
    _inferred__1_carry__0_i_8
       (.I0(_inferred__1_carry__0_i_12_n_0),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(_inferred__1_carry__0_i_16_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [4]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[4] ),
        .O(_inferred__1_carry__0_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__1_carry__0_i_9
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[7] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[7] ),
        .I5(\u_ras/u_ras_state/r_v1_y_reg_n_0_[7] ),
        .O(_inferred__1_carry__0_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__1_carry__1_i_1
       (.I0(\u_ras/u_ras_line/r_y0 [10]),
        .I1(_inferred__1_carry_i_9__9_n_0),
        .I2(\u_ras/u_ras_line/r_y1_reg_n_0_[10] ),
        .I3(_inferred__1_carry__1_i_8_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_1_in [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__1_carry__1_i_10
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[8] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[8] ),
        .I5(\u_ras/u_ras_state/r_v1_y_reg_n_0_[8] ),
        .O(_inferred__1_carry__1_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    _inferred__1_carry__1_i_11
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_v0_y_reg_n_0_[10] ),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[10] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[10] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__1_carry__1_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    _inferred__1_carry__1_i_12
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_v0_y_reg_n_0_[9] ),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[9] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[9] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__1_carry__1_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    _inferred__1_carry__1_i_13
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_v0_y_reg_n_0_[8] ),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[8] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[8] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__1_carry__1_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__1_carry__1_i_2
       (.I0(\u_ras/u_ras_line/r_y0 [9]),
        .I1(_inferred__1_carry_i_9__9_n_0),
        .I2(\u_ras/u_ras_line/r_y1_reg_n_0_[9] ),
        .I3(_inferred__1_carry__1_i_9_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_1_in [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__1_carry__1_i_3
       (.I0(\u_ras/u_ras_line/r_y0 [8]),
        .I1(_inferred__1_carry_i_9__9_n_0),
        .I2(\u_ras/u_ras_line/r_y1_reg_n_0_[8] ),
        .I3(_inferred__1_carry__1_i_10_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_1_in [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF90909F9)) 
    _inferred__1_carry__1_i_4
       (.I0(\u_ras/w_v1_y [11]),
        .I1(\u_ras/w_v0_y [11]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_y1_reg_n_0_[11] ),
        .I4(\u_ras/u_ras_line/r_y0 [11]),
        .O(_inferred__1_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDE1212DE)) 
    _inferred__1_carry__1_i_5
       (.I0(_inferred__1_carry__1_i_8_n_0),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(_inferred__1_carry__1_i_11_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [10]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[10] ),
        .O(_inferred__1_carry__1_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDE1212DE)) 
    _inferred__1_carry__1_i_6
       (.I0(_inferred__1_carry__1_i_9_n_0),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(_inferred__1_carry__1_i_12_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [9]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[9] ),
        .O(_inferred__1_carry__1_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDE1212DE)) 
    _inferred__1_carry__1_i_7
       (.I0(_inferred__1_carry__1_i_10_n_0),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(_inferred__1_carry__1_i_13_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [8]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[8] ),
        .O(_inferred__1_carry__1_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__1_carry__1_i_8
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[10] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[10] ),
        .I5(\u_ras/u_ras_state/r_v1_y_reg_n_0_[10] ),
        .O(_inferred__1_carry__1_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__1_carry__1_i_9
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[9] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[9] ),
        .I5(\u_ras/u_ras_state/r_v1_y_reg_n_0_[9] ),
        .O(_inferred__1_carry__1_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [4]),
        .O(_inferred__1_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    _inferred__1_carry_i_10
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [5]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [4]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [7]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [6]),
        .O(_inferred__1_carry_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    _inferred__1_carry_i_10__0
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [5]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [4]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [7]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [6]),
        .O(_inferred__1_carry_i_10__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    _inferred__1_carry_i_10__1
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [5]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [4]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [7]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [6]),
        .O(_inferred__1_carry_i_10__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__1_carry_i_10__10
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[3] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[3] ),
        .I5(\u_ras/u_ras_state/r_v1_y_reg_n_0_[3] ),
        .O(_inferred__1_carry_i_10__10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    _inferred__1_carry_i_10__2
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [5]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [4]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [7]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [6]),
        .O(_inferred__1_carry_i_10__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    _inferred__1_carry_i_10__3
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [5]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [4]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [7]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [6]),
        .O(_inferred__1_carry_i_10__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    _inferred__1_carry_i_10__4
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [5]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [4]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [7]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [6]),
        .O(_inferred__1_carry_i_10__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    _inferred__1_carry_i_10__5
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [5]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [4]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [7]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [6]),
        .O(_inferred__1_carry_i_10__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    _inferred__1_carry_i_10__6
       (.I0(\u_geo/u_geo_clip/r_exp_2z [3]),
        .I1(\u_geo/u_geo_clip/r_exp_2z [2]),
        .I2(\u_geo/u_geo_clip/r_exp_2z [4]),
        .I3(\u_geo/u_geo_clip/u_fadd/r_mats [16]),
        .I4(\u_geo/u_geo_clip/r_exp_2z [1]),
        .I5(\u_geo/u_geo_clip/r_exp_2z [0]),
        .O(_inferred__1_carry_i_10__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    _inferred__1_carry_i_10__7
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [5]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [4]),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [7]),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [6]),
        .O(_inferred__1_carry_i_10__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    _inferred__1_carry_i_10__8
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [9]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [8]),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [11]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [10]),
        .O(_inferred__1_carry_i_10__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    _inferred__1_carry_i_10__9
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [5]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [4]),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [7]),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [6]),
        .O(_inferred__1_carry_i_10__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00FF00FFFFFF0D)) 
    _inferred__1_carry_i_11
       (.I0(_inferred__1_carry_i_14_n_0),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [7]),
        .I2(\u_geo/u_geo_clip/u_fadd/r_mats [8]),
        .I3(_inferred__1_carry_i_15_n_0),
        .I4(\u_geo/u_geo_clip/u_fadd/r_mats [9]),
        .I5(_inferred__1_carry_i_16_n_0),
        .O(_inferred__1_carry_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    _inferred__1_carry_i_11__0
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [5]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [4]),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [7]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [6]),
        .O(_inferred__1_carry_i_11__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__1_carry_i_11__1
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[2] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[2] ),
        .I5(\u_ras/u_ras_state/r_v1_y_reg_n_0_[2] ),
        .O(_inferred__1_carry_i_11__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    _inferred__1_carry_i_12
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [8]),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [9]),
        .O(_inferred__1_carry_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    _inferred__1_carry_i_12__0
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [11]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [10]),
        .I2(_inferred__1_carry_i_13__0_n_0),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [8]),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [9]),
        .O(_inferred__1_carry_i_12__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__1_carry_i_12__1
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[1] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[1] ),
        .I5(\u_ras/u_ras_state/r_v1_y_reg_n_0_[1] ),
        .O(_inferred__1_carry_i_12__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111111110001)) 
    _inferred__1_carry_i_13
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [7]),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [6]),
        .I2(\u_geo/u_geo_clip/u_fadd/r_mats [2]),
        .I3(\u_geo/u_geo_clip/u_fadd/r_mats [3]),
        .I4(\u_geo/u_geo_clip/u_fadd/r_mats [4]),
        .I5(\u_geo/u_geo_clip/u_fadd/r_mats [5]),
        .O(_inferred__1_carry_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111111110001)) 
    _inferred__1_carry_i_13__0
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [7]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [6]),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [3]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [2]),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [4]),
        .I5(\u_geo/u_geo_viewport/u_fadd/r_mats [5]),
        .O(_inferred__1_carry_i_13__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__1_carry_i_13__1
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_ ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_ ),
        .I5(\u_ras/u_ras_state/r_v1_y_reg_n_0_ ),
        .O(_inferred__1_carry_i_13__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBABBBABABABBBABB)) 
    _inferred__1_carry_i_14
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [6]),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [5]),
        .I2(\u_geo/u_geo_clip/u_fadd/r_mats [4]),
        .I3(\u_geo/u_geo_clip/u_fadd/r_mats [3]),
        .I4(\u_geo/u_geo_clip/u_fadd/r_mats [2]),
        .I5(\u_geo/u_geo_clip/u_fadd/r_mats [1]),
        .O(_inferred__1_carry_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    _inferred__1_carry_i_14__0
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_v0_y_reg_n_0_[3] ),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[3] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[3] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__1_carry_i_14__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF0FFF0FFFFFFF4)) 
    _inferred__1_carry_i_15
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [12]),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [11]),
        .I2(\u_geo/u_geo_clip/u_fadd/r_mats [16]),
        .I3(\u_geo/u_geo_clip/u_fadd/r_mats [15]),
        .I4(\u_geo/u_geo_clip/u_fadd/r_mats [13]),
        .I5(\u_geo/u_geo_clip/u_fadd/r_mats [14]),
        .O(_inferred__1_carry_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    _inferred__1_carry_i_15__0
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_v0_y_reg_n_0_[2] ),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[2] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[2] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__1_carry_i_15__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    _inferred__1_carry_i_16
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [10]),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [14]),
        .I2(\u_geo/u_geo_clip/u_fadd/r_mats [12]),
        .O(_inferred__1_carry_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    _inferred__1_carry_i_16__0
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_v0_y_reg_n_0_[1] ),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[1] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_[1] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__1_carry_i_16__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    _inferred__1_carry_i_17
       (.I0(_inferred__1_carry_i_18_n_0),
        .I1(\u_ras/u_ras_state/r_v0_y_reg_n_0_ ),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_ ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_y_reg_n_0_ ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__1_carry_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0FFFA22CEF0CEFA)) 
    _inferred__1_carry_i_18
       (.I0(\u_ras/u_ras_line/w_sy_flag1__5 ),
        .I1(\u_ras/u_ras_state/p_1_in10_in ),
        .I2(\u_ras/u_ras_state/p_1_in1_in ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/p_0_in0_in ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__1_carry_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__0
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .O(_inferred__1_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__1
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [4]),
        .O(_inferred__1_carry_i_1__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__10
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .O(_inferred__1_carry_i_1__10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__11
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [4]),
        .O(_inferred__1_carry_i_1__11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__12
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .O(_inferred__1_carry_i_1__12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__13
       (.I0(\u_geo/u_geo_clip/r_exp_2z [4]),
        .O(_inferred__1_carry_i_1__13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__14
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [16]),
        .O(_inferred__1_carry_i_1__14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__15
       (.I0(\u_geo/u_geo_persdiv/r_ce_tmp_2z [4]),
        .O(_inferred__1_carry_i_1__15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__16
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .O(_inferred__1_carry_i_1__16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__17
       (.I0(\u_geo/u_geo_viewport/r_exp_2z [4]),
        .O(_inferred__1_carry_i_1__17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__18
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .O(_inferred__1_carry_i_1__18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__19
       (.I0(\u_geo/u_geo_viewport/r_ce_tmp_2z [4]),
        .O(_inferred__1_carry_i_1__19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__2
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .O(_inferred__1_carry_i_1__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__20
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .O(_inferred__1_carry_i_1__20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__1_carry_i_1__21
       (.I0(\u_ras/u_ras_line/r_y0 [3]),
        .I1(_inferred__1_carry_i_9__9_n_0),
        .I2(\u_ras/u_ras_line/r_y1_reg_n_0_[3] ),
        .I3(_inferred__1_carry_i_10__10_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_1_in [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__3
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [4]),
        .O(_inferred__1_carry_i_1__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__4
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .O(_inferred__1_carry_i_1__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__5
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [4]),
        .O(_inferred__1_carry_i_1__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__6
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .O(_inferred__1_carry_i_1__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__7
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [4]),
        .O(_inferred__1_carry_i_1__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__8
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .O(_inferred__1_carry_i_1__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    _inferred__1_carry_i_1__9
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [4]),
        .O(_inferred__1_carry_i_1__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    _inferred__1_carry_i_2
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I1(_inferred__1_carry_i_6_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [3]),
        .O(_inferred__1_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    _inferred__1_carry_i_2__0
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I1(_inferred__1_carry_i_6__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [3]),
        .O(_inferred__1_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    _inferred__1_carry_i_2__1
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I1(_inferred__1_carry_i_6__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [3]),
        .O(_inferred__1_carry_i_2__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__1_carry_i_2__10
       (.I0(\u_ras/u_ras_line/r_y0 [2]),
        .I1(_inferred__1_carry_i_9__9_n_0),
        .I2(\u_ras/u_ras_line/r_y1_reg_n_0_[2] ),
        .I3(_inferred__1_carry_i_11__1_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_1_in [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    _inferred__1_carry_i_2__11
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [4]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .O(_inferred__1_carry_i_2__11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    _inferred__1_carry_i_2__12
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [4]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .O(_inferred__1_carry_i_2__12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    _inferred__1_carry_i_2__13
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [4]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .O(_inferred__1_carry_i_2__13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    _inferred__1_carry_i_2__14
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [4]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .O(_inferred__1_carry_i_2__14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    _inferred__1_carry_i_2__15
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [4]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .O(_inferred__1_carry_i_2__15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    _inferred__1_carry_i_2__16
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [4]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .O(_inferred__1_carry_i_2__16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    _inferred__1_carry_i_2__17
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [4]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .O(_inferred__1_carry_i_2__17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    _inferred__1_carry_i_2__18
       (.I0(\u_geo/u_geo_clip/r_exp_2z [4]),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [16]),
        .O(_inferred__1_carry_i_2__18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    _inferred__1_carry_i_2__19
       (.I0(\u_geo/u_geo_persdiv/r_ce_tmp_2z [4]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .O(_inferred__1_carry_i_2__19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    _inferred__1_carry_i_2__2
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I1(_inferred__1_carry_i_6__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [3]),
        .O(_inferred__1_carry_i_2__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    _inferred__1_carry_i_2__20
       (.I0(\u_geo/u_geo_viewport/r_exp_2z [4]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .O(_inferred__1_carry_i_2__20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    _inferred__1_carry_i_2__21
       (.I0(\u_geo/u_geo_viewport/r_ce_tmp_2z [4]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .O(_inferred__1_carry_i_2__21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    _inferred__1_carry_i_2__3
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I1(_inferred__1_carry_i_6__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [3]),
        .O(_inferred__1_carry_i_2__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    _inferred__1_carry_i_2__4
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I1(_inferred__1_carry_i_6__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [3]),
        .O(_inferred__1_carry_i_2__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    _inferred__1_carry_i_2__5
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I1(_inferred__1_carry_i_6__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [3]),
        .O(_inferred__1_carry_i_2__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    _inferred__1_carry_i_2__6
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [16]),
        .I1(\r_c[21]_i_3_n_0 ),
        .I2(\u_geo/u_geo_clip/r_exp_2z [3]),
        .O(_inferred__1_carry_i_2__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    _inferred__1_carry_i_2__7
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I1(_inferred__1_carry_i_6__7_n_0),
        .I2(\u_geo/u_geo_persdiv/r_ce_tmp_2z [3]),
        .O(_inferred__1_carry_i_2__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    _inferred__1_carry_i_2__8
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I1(_inferred__1_carry_i_6__8_n_0),
        .I2(\u_geo/u_geo_viewport/r_exp_2z [3]),
        .O(_inferred__1_carry_i_2__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB4)) 
    _inferred__1_carry_i_2__9
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I1(_inferred__1_carry_i_6__9_n_0),
        .I2(\u_geo/u_geo_viewport/r_ce_tmp_2z [3]),
        .O(_inferred__1_carry_i_2__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_3
       (.I0(_inferred__1_carry_i_7_n_0),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [2]),
        .O(_inferred__1_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_3__0
       (.I0(_inferred__1_carry_i_7__0_n_0),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [2]),
        .O(_inferred__1_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_3__1
       (.I0(_inferred__1_carry_i_7__1_n_0),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [2]),
        .O(_inferred__1_carry_i_3__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__1_carry_i_3__10
       (.I0(\u_ras/u_ras_line/r_y0 [1]),
        .I1(_inferred__1_carry_i_9__9_n_0),
        .I2(\u_ras/u_ras_line/r_y1_reg_n_0_[1] ),
        .I3(_inferred__1_carry_i_12__1_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_1_in [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_3__2
       (.I0(_inferred__1_carry_i_7__2_n_0),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [2]),
        .O(_inferred__1_carry_i_3__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_3__3
       (.I0(_inferred__1_carry_i_7__3_n_0),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [2]),
        .O(_inferred__1_carry_i_3__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_3__4
       (.I0(_inferred__1_carry_i_7__4_n_0),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [2]),
        .O(_inferred__1_carry_i_3__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_3__5
       (.I0(_inferred__1_carry_i_7__5_n_0),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [2]),
        .O(_inferred__1_carry_i_3__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF0700F8)) 
    _inferred__1_carry_i_3__6
       (.I0(_inferred__1_carry_i_6__6_n_0),
        .I1(_inferred__1_carry_i_7__6_n_0),
        .I2(_inferred__1_carry_i_8__6_n_0),
        .I3(\u_geo/u_geo_clip/u_fadd/r_mats [16]),
        .I4(\u_geo/u_geo_clip/r_exp_2z [2]),
        .O(_inferred__1_carry_i_3__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_3__7
       (.I0(_inferred__1_carry_i_7__7_n_0),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I2(\u_geo/u_geo_persdiv/r_ce_tmp_2z [2]),
        .O(_inferred__1_carry_i_3__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_3__8
       (.I0(_inferred__1_carry_i_7__8_n_0),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I2(\u_geo/u_geo_viewport/r_exp_2z [2]),
        .O(_inferred__1_carry_i_3__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_3__9
       (.I0(_inferred__1_carry_i_7__9_n_0),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I2(\u_geo/u_geo_viewport/r_ce_tmp_2z [2]),
        .O(_inferred__1_carry_i_3__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_4
       (.I0(\r_c[1]_i_3_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [1]),
        .O(_inferred__1_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_4__0
       (.I0(\r_c[1]_i_3__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [1]),
        .O(_inferred__1_carry_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_4__1
       (.I0(\r_c[1]_i_3__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [1]),
        .O(_inferred__1_carry_i_4__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__1_carry_i_4__10
       (.I0(\u_ras/u_ras_line/r_y0 [0]),
        .I1(_inferred__1_carry_i_9__9_n_0),
        .I2(\u_ras/u_ras_line/r_y1_reg_n_0_ ),
        .I3(_inferred__1_carry_i_13__1_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_1_in [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_4__2
       (.I0(\r_c[1]_i_3__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [1]),
        .O(_inferred__1_carry_i_4__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_4__3
       (.I0(\r_c[1]_i_3__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [1]),
        .O(_inferred__1_carry_i_4__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_4__4
       (.I0(\r_c[1]_i_3__4_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [1]),
        .O(_inferred__1_carry_i_4__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_4__5
       (.I0(\r_c[1]_i_3__5_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [1]),
        .O(_inferred__1_carry_i_4__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF0200FD)) 
    _inferred__1_carry_i_4__6
       (.I0(_inferred__1_carry_i_9__6_n_0),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [14]),
        .I2(\u_geo/u_geo_clip/u_fadd/r_mats [15]),
        .I3(\u_geo/u_geo_clip/u_fadd/r_mats [16]),
        .I4(\u_geo/u_geo_clip/r_exp_2z [1]),
        .O(_inferred__1_carry_i_4__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_4__7
       (.I0(\r_c[1]_i_3__6_n_0 ),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I2(\u_geo/u_geo_persdiv/r_ce_tmp_2z [1]),
        .O(_inferred__1_carry_i_4__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_4__8
       (.I0(_inferred__1_carry_i_8__8_n_0),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I2(\u_geo/u_geo_viewport/r_exp_2z [1]),
        .O(_inferred__1_carry_i_4__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    _inferred__1_carry_i_4__9
       (.I0(\r_c[1]_i_3__7_n_0 ),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I2(\u_geo/u_geo_viewport/r_ce_tmp_2z [1]),
        .O(_inferred__1_carry_i_4__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDE1212DE)) 
    _inferred__1_carry_i_5
       (.I0(_inferred__1_carry_i_10__10_n_0),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(_inferred__1_carry_i_14__0_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [3]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[3] ),
        .O(_inferred__1_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hD1)) 
    _inferred__1_carry_i_5__0
       (.I0(\r_c[14]_i_4_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I2(_inferred__1_carry_i_8_n_0),
        .O(_inferred__1_carry_i_5__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hD1)) 
    _inferred__1_carry_i_5__1
       (.I0(\r_c[14]_i_4__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I2(_inferred__1_carry_i_8__0_n_0),
        .O(_inferred__1_carry_i_5__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE3)) 
    _inferred__1_carry_i_5__10
       (.I0(w_cf_tmp_i_33__2_n_0),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I2(_inferred__1_carry_i_9__10_n_0),
        .O(_inferred__1_carry_i_5__10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hD1)) 
    _inferred__1_carry_i_5__2
       (.I0(\r_c[14]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I2(_inferred__1_carry_i_8__1_n_0),
        .O(_inferred__1_carry_i_5__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hD1)) 
    _inferred__1_carry_i_5__3
       (.I0(\r_c[14]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I2(_inferred__1_carry_i_8__2_n_0),
        .O(_inferred__1_carry_i_5__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hD1)) 
    _inferred__1_carry_i_5__4
       (.I0(\r_c[14]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I2(_inferred__1_carry_i_8__3_n_0),
        .O(_inferred__1_carry_i_5__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hD1)) 
    _inferred__1_carry_i_5__5
       (.I0(\r_c[14]_i_4__4_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I2(_inferred__1_carry_i_8__4_n_0),
        .O(_inferred__1_carry_i_5__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hD1)) 
    _inferred__1_carry_i_5__6
       (.I0(\r_c[14]_i_4__5_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I2(_inferred__1_carry_i_8__5_n_0),
        .O(_inferred__1_carry_i_5__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h65)) 
    _inferred__1_carry_i_5__7
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [16]),
        .I1(_inferred__1_carry_i_10__6_n_0),
        .I2(_inferred__1_carry_i_11_n_0),
        .O(_inferred__1_carry_i_5__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hD1)) 
    _inferred__1_carry_i_5__8
       (.I0(\r_c[14]_i_4__7_n_0 ),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I2(_inferred__1_carry_i_8__7_n_0),
        .O(_inferred__1_carry_i_5__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hD1)) 
    _inferred__1_carry_i_5__9
       (.I0(\r_c[14]_i_4__8_n_0 ),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I2(_inferred__1_carry_i_8__9_n_0),
        .O(_inferred__1_carry_i_5__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    _inferred__1_carry_i_6
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [13]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [15]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_9_n_0),
        .O(_inferred__1_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    _inferred__1_carry_i_6__0
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [13]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [15]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_9__0_n_0),
        .O(_inferred__1_carry_i_6__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    _inferred__1_carry_i_6__1
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [13]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [15]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_9__1_n_0),
        .O(_inferred__1_carry_i_6__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDE1212DE)) 
    _inferred__1_carry_i_6__10
       (.I0(_inferred__1_carry_i_11__1_n_0),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(_inferred__1_carry_i_15__0_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [2]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[2] ),
        .O(_inferred__1_carry_i_6__10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    _inferred__1_carry_i_6__2
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [13]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [15]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_9__2_n_0),
        .O(_inferred__1_carry_i_6__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    _inferred__1_carry_i_6__3
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [12]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [13]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [15]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [14]),
        .I4(_inferred__1_carry_i_9__3_n_0),
        .O(_inferred__1_carry_i_6__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    _inferred__1_carry_i_6__4
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [12]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [13]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [15]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [14]),
        .I4(_inferred__1_carry_i_9__4_n_0),
        .O(_inferred__1_carry_i_6__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    _inferred__1_carry_i_6__5
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [12]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [13]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [15]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [14]),
        .I4(_inferred__1_carry_i_9__5_n_0),
        .O(_inferred__1_carry_i_6__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    _inferred__1_carry_i_6__6
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [5]),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [4]),
        .I2(\u_geo/u_geo_clip/u_fadd/r_mats [7]),
        .I3(\u_geo/u_geo_clip/u_fadd/r_mats [6]),
        .O(_inferred__1_carry_i_6__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    _inferred__1_carry_i_6__7
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [13]),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [15]),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_9__7_n_0),
        .O(_inferred__1_carry_i_6__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    _inferred__1_carry_i_6__8
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [12]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [13]),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [15]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [14]),
        .I4(_inferred__1_carry_i_10__8_n_0),
        .O(_inferred__1_carry_i_6__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    _inferred__1_carry_i_6__9
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [13]),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [15]),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_9__8_n_0),
        .O(_inferred__1_carry_i_6__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100010001)) 
    _inferred__1_carry_i_7
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [13]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [15]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_10_n_0),
        .I5(_inferred__1_carry_i_9_n_0),
        .O(_inferred__1_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100010001)) 
    _inferred__1_carry_i_7__0
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [13]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [15]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_10__0_n_0),
        .I5(_inferred__1_carry_i_9__0_n_0),
        .O(_inferred__1_carry_i_7__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100010001)) 
    _inferred__1_carry_i_7__1
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [13]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [15]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_10__1_n_0),
        .I5(_inferred__1_carry_i_9__1_n_0),
        .O(_inferred__1_carry_i_7__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDE1212DE)) 
    _inferred__1_carry_i_7__10
       (.I0(_inferred__1_carry_i_12__1_n_0),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(_inferred__1_carry_i_16__0_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [1]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[1] ),
        .O(_inferred__1_carry_i_7__10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100010001)) 
    _inferred__1_carry_i_7__2
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [13]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [15]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_10__2_n_0),
        .I5(_inferred__1_carry_i_9__2_n_0),
        .O(_inferred__1_carry_i_7__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100010001)) 
    _inferred__1_carry_i_7__3
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [12]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [13]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [15]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [14]),
        .I4(_inferred__1_carry_i_10__3_n_0),
        .I5(_inferred__1_carry_i_9__3_n_0),
        .O(_inferred__1_carry_i_7__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100010001)) 
    _inferred__1_carry_i_7__4
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [12]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [13]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [15]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [14]),
        .I4(_inferred__1_carry_i_10__4_n_0),
        .I5(_inferred__1_carry_i_9__4_n_0),
        .O(_inferred__1_carry_i_7__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100010001)) 
    _inferred__1_carry_i_7__5
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [12]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [13]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [15]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [14]),
        .I4(_inferred__1_carry_i_10__5_n_0),
        .I5(_inferred__1_carry_i_9__5_n_0),
        .O(_inferred__1_carry_i_7__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    _inferred__1_carry_i_7__6
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [9]),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [8]),
        .I2(\u_geo/u_geo_clip/u_fadd/r_mats [11]),
        .I3(\u_geo/u_geo_clip/u_fadd/r_mats [10]),
        .O(_inferred__1_carry_i_7__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100010001)) 
    _inferred__1_carry_i_7__7
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [13]),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [15]),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_10__7_n_0),
        .I5(_inferred__1_carry_i_9__7_n_0),
        .O(_inferred__1_carry_i_7__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100010001)) 
    _inferred__1_carry_i_7__8
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [12]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [13]),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [15]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [14]),
        .I4(_inferred__1_carry_i_11__0_n_0),
        .I5(_inferred__1_carry_i_10__8_n_0),
        .O(_inferred__1_carry_i_7__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100010001)) 
    _inferred__1_carry_i_7__9
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [13]),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [15]),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_10__9_n_0),
        .I5(_inferred__1_carry_i_9__8_n_0),
        .O(_inferred__1_carry_i_7__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    _inferred__1_carry_i_8
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [3]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [4]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [1]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [0]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [2]),
        .O(_inferred__1_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    _inferred__1_carry_i_8__0
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [3]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [4]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [1]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [0]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [2]),
        .O(_inferred__1_carry_i_8__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    _inferred__1_carry_i_8__1
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [3]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [4]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [1]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [0]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [2]),
        .O(_inferred__1_carry_i_8__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDE1212DE)) 
    _inferred__1_carry_i_8__10
       (.I0(_inferred__1_carry_i_13__1_n_0),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(_inferred__1_carry_i_17_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [0]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_ ),
        .O(_inferred__1_carry_i_8__10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    _inferred__1_carry_i_8__2
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [3]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [4]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [1]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [0]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [2]),
        .O(_inferred__1_carry_i_8__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    _inferred__1_carry_i_8__3
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [3]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [4]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [1]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [0]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [2]),
        .O(_inferred__1_carry_i_8__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    _inferred__1_carry_i_8__4
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [3]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [4]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [1]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [0]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [2]),
        .O(_inferred__1_carry_i_8__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    _inferred__1_carry_i_8__5
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [3]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [4]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [1]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [0]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [2]),
        .O(_inferred__1_carry_i_8__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    _inferred__1_carry_i_8__6
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [13]),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [12]),
        .I2(\u_geo/u_geo_clip/u_fadd/r_mats [14]),
        .I3(\u_geo/u_geo_clip/u_fadd/r_mats [15]),
        .O(_inferred__1_carry_i_8__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    _inferred__1_carry_i_8__7
       (.I0(\u_geo/u_geo_persdiv/r_ce_tmp_2z [0]),
        .I1(\u_geo/u_geo_persdiv/r_ce_tmp_2z [4]),
        .I2(\u_geo/u_geo_persdiv/r_ce_tmp_2z [3]),
        .I3(\u_geo/u_geo_persdiv/r_ce_tmp_2z [1]),
        .I4(\u_geo/u_geo_persdiv/r_ce_tmp_2z [2]),
        .O(_inferred__1_carry_i_8__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    _inferred__1_carry_i_8__8
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [14]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [15]),
        .I2(_inferred__1_carry_i_12__0_n_0),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [12]),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [13]),
        .O(_inferred__1_carry_i_8__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    _inferred__1_carry_i_8__9
       (.I0(\u_geo/u_geo_viewport/r_ce_tmp_2z [0]),
        .I1(\u_geo/u_geo_viewport/r_ce_tmp_2z [4]),
        .I2(\u_geo/u_geo_viewport/r_ce_tmp_2z [3]),
        .I3(\u_geo/u_geo_viewport/r_ce_tmp_2z [1]),
        .I4(\u_geo/u_geo_viewport/r_ce_tmp_2z [2]),
        .O(_inferred__1_carry_i_8__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    _inferred__1_carry_i_9
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [8]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [11]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [10]),
        .O(_inferred__1_carry_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    _inferred__1_carry_i_9__0
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [8]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [11]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [10]),
        .O(_inferred__1_carry_i_9__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    _inferred__1_carry_i_9__1
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [8]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [11]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [10]),
        .O(_inferred__1_carry_i_9__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    _inferred__1_carry_i_9__10
       (.I0(\u_geo/u_geo_viewport/r_exp_2z [2]),
        .I1(\u_geo/u_geo_viewport/r_exp_2z [1]),
        .I2(\u_geo/u_geo_viewport/r_exp_2z [3]),
        .I3(\u_geo/u_geo_viewport/r_exp_2z [4]),
        .I4(\u_geo/u_geo_viewport/r_exp_2z [0]),
        .I5(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .O(_inferred__1_carry_i_9__10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    _inferred__1_carry_i_9__2
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [8]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [11]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [10]),
        .O(_inferred__1_carry_i_9__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    _inferred__1_carry_i_9__3
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [9]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [8]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [11]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [10]),
        .O(_inferred__1_carry_i_9__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    _inferred__1_carry_i_9__4
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [9]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [8]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [11]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [10]),
        .O(_inferred__1_carry_i_9__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    _inferred__1_carry_i_9__5
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [9]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [8]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [11]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [10]),
        .O(_inferred__1_carry_i_9__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEEEEEEFFEF)) 
    _inferred__1_carry_i_9__6
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [13]),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [12]),
        .I2(_inferred__1_carry_i_12_n_0),
        .I3(_inferred__1_carry_i_13_n_0),
        .I4(\u_geo/u_geo_clip/u_fadd/r_mats [10]),
        .I5(\u_geo/u_geo_clip/u_fadd/r_mats [11]),
        .O(_inferred__1_carry_i_9__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    _inferred__1_carry_i_9__7
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [8]),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [11]),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [10]),
        .O(_inferred__1_carry_i_9__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    _inferred__1_carry_i_9__8
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [8]),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [11]),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [10]),
        .O(_inferred__1_carry_i_9__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAE)) 
    _inferred__1_carry_i_9__9
       (.I0(\u_ras/u_ras_line/r_y0 [11]),
        .I1(\u_ras/u_ras_line/w_sy_flag1__5 ),
        .I2(\u_ras/u_ras_line/r_y1_reg_n_0_[11] ),
        .O(_inferred__1_carry_i_9__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__5_carry__0_i_1
       (.I0(\u_ras/u_ras_line/r_x0 [7]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x1 [7]),
        .I3(_inferred__5_carry__0_i_9_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_2_in [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__5_carry__0_i_10
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[6] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[6] ),
        .I5(\u_ras/u_ras_state/r_v1_x_reg_n_0_[6] ),
        .O(_inferred__5_carry__0_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__5_carry__0_i_11
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[5] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[5] ),
        .I5(\u_ras/u_ras_state/r_v1_x_reg_n_0_[5] ),
        .O(_inferred__5_carry__0_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__5_carry__0_i_12
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[4] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[4] ),
        .I5(\u_ras/u_ras_state/r_v1_x_reg_n_0_[4] ),
        .O(_inferred__5_carry__0_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "_inferred__5_carry__0_i_1" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__5_carry__0_i_1_replica
       (.I0(\u_ras/u_ras_line/r_x0 [7]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x1 [7]),
        .I3(_inferred__5_carry__0_i_9_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_2_in[7]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__5_carry__0_i_2
       (.I0(\u_ras/u_ras_line/r_x0 [6]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x1 [6]),
        .I3(_inferred__5_carry__0_i_10_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_2_in [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__5_carry__0_i_3
       (.I0(\u_ras/u_ras_line/r_x0 [5]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x1 [5]),
        .I3(_inferred__5_carry__0_i_11_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_2_in [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__5_carry__0_i_4
       (.I0(\u_ras/u_ras_line/r_x0 [4]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x1 [4]),
        .I3(_inferred__5_carry__0_i_12_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_2_in [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    _inferred__5_carry__0_i_5
       (.I0(\u_ras/p_2_in[7]_repN ),
        .I1(w_err__0_carry__0_i_12_n_0),
        .O(_inferred__5_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    _inferred__5_carry__0_i_6
       (.I0(\u_ras/p_2_in [6]),
        .I1(w_err__0_carry__0_i_9_n_0),
        .O(_inferred__5_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    _inferred__5_carry__0_i_7
       (.I0(\u_ras/p_2_in [5]),
        .I1(w_err__0_carry__0_i_10_n_0),
        .O(_inferred__5_carry__0_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    _inferred__5_carry__0_i_8
       (.I0(\u_ras/p_2_in [4]),
        .I1(w_err__0_carry__0_i_11_n_0),
        .O(_inferred__5_carry__0_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__5_carry__0_i_9
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[7] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[7] ),
        .I5(\u_ras/u_ras_state/r_v1_x_reg_n_0_[7] ),
        .O(_inferred__5_carry__0_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__5_carry__1_i_1
       (.I0(\u_ras/u_ras_line/r_x0 [10]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x1 [10]),
        .I3(_inferred__5_carry__1_i_8_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_2_in [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__5_carry__1_i_10
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[8] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[8] ),
        .I5(\u_ras/u_ras_state/r_v1_x_reg_n_0_[8] ),
        .O(_inferred__5_carry__1_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__5_carry__1_i_2
       (.I0(\u_ras/u_ras_line/r_x0 [9]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x1 [9]),
        .I3(_inferred__5_carry__1_i_9_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_2_in [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__5_carry__1_i_3
       (.I0(\u_ras/u_ras_line/r_x0 [8]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x1 [8]),
        .I3(_inferred__5_carry__1_i_10_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_2_in [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF90909F9)) 
    _inferred__5_carry__1_i_4
       (.I0(\u_ras/w_v1_x [11]),
        .I1(\u_ras/w_v0_x [11]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_x1 [11]),
        .I4(\u_ras/u_ras_line/r_x0 [11]),
        .O(_inferred__5_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    _inferred__5_carry__1_i_5
       (.I0(\u_ras/p_2_in [10]),
        .I1(w_err__0_carry__1_i_8_n_0),
        .O(_inferred__5_carry__1_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    _inferred__5_carry__1_i_6
       (.I0(\u_ras/p_2_in [9]),
        .I1(w_err__0_carry__1_i_7_n_0),
        .O(_inferred__5_carry__1_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    _inferred__5_carry__1_i_7
       (.I0(\u_ras/p_2_in [8]),
        .I1(w_err__0_carry__1_i_6_n_0),
        .O(_inferred__5_carry__1_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__5_carry__1_i_8
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[10] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[10] ),
        .I5(\u_ras/u_ras_state/r_v1_x_reg_n_0_[10] ),
        .O(_inferred__5_carry__1_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__5_carry__1_i_9
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[9] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[9] ),
        .I5(\u_ras/u_ras_state/r_v1_x_reg_n_0_[9] ),
        .O(_inferred__5_carry__1_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__5_carry_i_1
       (.I0(\u_ras/u_ras_line/r_x0 [3]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x1 [3]),
        .I3(_inferred__5_carry_i_10_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_2_in [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__5_carry_i_10
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[3] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[3] ),
        .I5(\u_ras/u_ras_state/r_v1_x_reg_n_0_[3] ),
        .O(_inferred__5_carry_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__5_carry_i_11
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[2] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[2] ),
        .I5(\u_ras/u_ras_state/r_v1_x_reg_n_0_[2] ),
        .O(_inferred__5_carry_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__5_carry_i_12
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[1] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[1] ),
        .I5(\u_ras/u_ras_state/r_v1_x_reg_n_0_[1] ),
        .O(_inferred__5_carry_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04099D2B264DBF6F)) 
    _inferred__5_carry_i_13
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_ ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_ ),
        .I5(\u_ras/u_ras_state/r_v1_x_reg_n_0_ ),
        .O(_inferred__5_carry_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0FFFA22CEF0CEFA)) 
    _inferred__5_carry_i_14
       (.I0(\u_ras/u_ras_line/w_sx_flag1__5 ),
        .I1(\u_ras/u_ras_state/p_1_in8_in ),
        .I2(\u_ras/u_ras_state/p_1_in ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/p_0_in ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(_inferred__5_carry_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__5_carry_i_2
       (.I0(\u_ras/u_ras_line/r_x0 [2]),
        .I1(_inferred__5_carry_i_9_n_0_repN),
        .I2(\u_ras/u_ras_line/r_x1 [2]),
        .I3(_inferred__5_carry_i_11_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_2_in [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__5_carry_i_3
       (.I0(\u_ras/u_ras_line/r_x0 [1]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x1 [1]),
        .I3(_inferred__5_carry_i_12_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_2_in [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4747FF00)) 
    _inferred__5_carry_i_4
       (.I0(\u_ras/u_ras_line/r_x0 [0]),
        .I1(_inferred__5_carry_i_9_n_0_repN),
        .I2(\u_ras/u_ras_line/r_x1 [0]),
        .I3(_inferred__5_carry_i_13_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/p_2_in [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    _inferred__5_carry_i_5
       (.I0(\u_ras/p_2_in [3]),
        .I1(w_err__0_carry_i_11_n_0),
        .O(_inferred__5_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    _inferred__5_carry_i_6
       (.I0(\u_ras/p_2_in [2]),
        .I1(w_err__0_carry_i_8_n_0),
        .O(_inferred__5_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    _inferred__5_carry_i_7
       (.I0(\u_ras/p_2_in [1]),
        .I1(w_err__0_carry_i_9_n_0),
        .O(_inferred__5_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    _inferred__5_carry_i_8
       (.I0(\u_ras/p_2_in [0]),
        .I1(w_err__0_carry_i_10_n_0),
        .O(_inferred__5_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAE)) 
    _inferred__5_carry_i_9
       (.I0(\u_ras/u_ras_line/r_x0 [11]),
        .I1(\u_ras/u_ras_line/w_sx_flag1__5 ),
        .I2(\u_ras/u_ras_line/r_x1 [11]),
        .O(_inferred__5_carry_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "_inferred__5_carry_i_9" *) 
  LUT3 #(
    .INIT(8'hAE)) 
    _inferred__5_carry_i_9_replica
       (.I0(\u_ras/u_ras_line/r_x0 [11]),
        .I1(\u_ras/u_ras_line/w_sx_flag1__5 ),
        .I2(\u_ras/u_ras_line/r_x1 [11]),
        .O(_inferred__5_carry_i_9_n_0_repN));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8080000A808AAAA)) 
    _inferred__8__0_carry__0_i_1
       (.I0(\u_ras/w_e2 [7]),
        .I1(\u_ras/w_err [6]),
        .I2(_inferred__8__0_carry_i_8_n_0),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__0_n_5 ),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .I5(\u_ras/w_dy [6]),
        .O(_inferred__8__0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD400D4D4D4000000)) 
    _inferred__8__0_carry__0_i_10
       (.I0(\u_ras/u_ras_line/w_dx ),
        .I1(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I2(\u_ras/u_ras_line/r_e2 ),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__0_n_5 ),
        .I4(_inferred__8__0_carry_i_8_n_0),
        .I5(\u_ras/w_err [6]),
        .O(_inferred__8__0_carry__0_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD400D4D4D4000000)) 
    _inferred__8__0_carry__0_i_11
       (.I0(\u_ras/u_ras_line/w_dx ),
        .I1(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I2(\u_ras/u_ras_line/r_e2 ),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__0_n_6 ),
        .I4(_inferred__8__0_carry_i_8_n_0),
        .I5(\u_ras/w_err [5]),
        .O(_inferred__8__0_carry__0_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD400D4D4D4000000)) 
    _inferred__8__0_carry__0_i_12
       (.I0(\u_ras/u_ras_line/w_dx ),
        .I1(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I2(\u_ras/u_ras_line/r_e2 ),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__0_n_7 ),
        .I4(_inferred__8__0_carry_i_8_n_0),
        .I5(\u_ras/w_err [4]),
        .O(_inferred__8__0_carry__0_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8080000A808AAAA)) 
    _inferred__8__0_carry__0_i_2
       (.I0(\u_ras/w_e2 [6]),
        .I1(\u_ras/w_err [5]),
        .I2(_inferred__8__0_carry_i_8_n_0),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__0_n_6 ),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .I5(\u_ras/w_dy [5]),
        .O(_inferred__8__0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8080000A808AAAA)) 
    _inferred__8__0_carry__0_i_3
       (.I0(\u_ras/w_e2 [5]),
        .I1(\u_ras/w_err [4]),
        .I2(_inferred__8__0_carry_i_8_n_0),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__0_n_7 ),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .I5(\u_ras/w_dy [4]),
        .O(_inferred__8__0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8080000A808AAAA)) 
    _inferred__8__0_carry__0_i_4
       (.I0(\u_ras/w_e2 [4]),
        .I1(\u_ras/w_err [3]),
        .I2(_inferred__8__0_carry_i_8_n_0),
        .I3(\u_ras/u_ras_line/_inferred__5_carry_n_4 ),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .I5(\u_ras/w_dy [3]),
        .O(_inferred__8__0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96969669)) 
    _inferred__8__0_carry__0_i_5
       (.I0(_inferred__8__0_carry__0_i_1_n_0),
        .I1(_inferred__8__0_carry__0_i_9_n_0),
        .I2(\u_ras/w_e2 [8]),
        .I3(\u_ras/w_dy [7]),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .O(_inferred__8__0_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96969669)) 
    _inferred__8__0_carry__0_i_6
       (.I0(_inferred__8__0_carry__0_i_2_n_0),
        .I1(_inferred__8__0_carry__0_i_10_n_0),
        .I2(\u_ras/w_e2 [7]),
        .I3(\u_ras/w_dy [6]),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .O(_inferred__8__0_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96969669)) 
    _inferred__8__0_carry__0_i_7
       (.I0(_inferred__8__0_carry__0_i_3_n_0),
        .I1(_inferred__8__0_carry__0_i_11_n_0),
        .I2(\u_ras/w_e2 [6]),
        .I3(\u_ras/w_dy [5]),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .O(_inferred__8__0_carry__0_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96969669)) 
    _inferred__8__0_carry__0_i_8
       (.I0(_inferred__8__0_carry__0_i_4_n_0),
        .I1(_inferred__8__0_carry__0_i_12_n_0),
        .I2(\u_ras/w_e2 [5]),
        .I3(\u_ras/w_dy [4]),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .O(_inferred__8__0_carry__0_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD400D4D4D4000000)) 
    _inferred__8__0_carry__0_i_9
       (.I0(\u_ras/u_ras_line/w_dx ),
        .I1(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I2(\u_ras/u_ras_line/r_e2 ),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__0_n_4 ),
        .I4(_inferred__8__0_carry_i_8_n_0),
        .I5(\u_ras/w_err [7]),
        .O(_inferred__8__0_carry__0_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8080000A808AAAA)) 
    _inferred__8__0_carry__1_i_1
       (.I0(\u_ras/w_e2 [9]),
        .I1(\u_ras/w_err [8]),
        .I2(_inferred__8__0_carry_i_8_n_0),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__1_n_7 ),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .I5(\u_ras/w_dy [8]),
        .O(_inferred__8__0_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8080000A808AAAA)) 
    _inferred__8__0_carry__1_i_2
       (.I0(\u_ras/w_e2 [8]),
        .I1(\u_ras/w_err [7]),
        .I2(_inferred__8__0_carry_i_8_n_0),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__0_n_4 ),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .I5(\u_ras/w_dy [7]),
        .O(_inferred__8__0_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0EEFF110)) 
    _inferred__8__0_carry__1_i_3
       (.I0(\u_ras/w_dy [9]),
        .I1(\u_ras/u_ras_line/p_0_in ),
        .I2(_inferred__8__0_carry__1_i_6_n_0),
        .I3(\u_ras/w_e2 [10]),
        .I4(_inferred__8__0_carry__1_i_7_n_0),
        .O(_inferred__8__0_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96969669)) 
    _inferred__8__0_carry__1_i_4
       (.I0(_inferred__8__0_carry__1_i_1_n_0),
        .I1(_inferred__8__0_carry__1_i_6_n_0),
        .I2(\u_ras/w_e2 [10]),
        .I3(\u_ras/w_dy [9]),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .O(_inferred__8__0_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96969669)) 
    _inferred__8__0_carry__1_i_5
       (.I0(_inferred__8__0_carry__1_i_2_n_0),
        .I1(_inferred__8__0_carry__1_i_8_n_0),
        .I2(\u_ras/w_e2 [9]),
        .I3(\u_ras/w_dy [8]),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .O(_inferred__8__0_carry__1_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD400D4D4D4000000)) 
    _inferred__8__0_carry__1_i_6
       (.I0(\u_ras/u_ras_line/w_dx ),
        .I1(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I2(\u_ras/u_ras_line/r_e2 ),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__1_n_6 ),
        .I4(_inferred__8__0_carry_i_8_n_0),
        .I5(\u_ras/w_err [9]),
        .O(_inferred__8__0_carry__1_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h39C9393939C9C9C9)) 
    _inferred__8__0_carry__1_i_7
       (.I0(\u_ras/w_dy [10]),
        .I1(\u_ras/w_e2 [11]),
        .I2(\u_ras/u_ras_line/p_0_in ),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__1_n_5 ),
        .I4(_inferred__8__0_carry_i_8_n_0),
        .I5(\u_ras/w_err [10]),
        .O(_inferred__8__0_carry__1_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD400D4D4D4000000)) 
    _inferred__8__0_carry__1_i_8
       (.I0(\u_ras/u_ras_line/w_dx ),
        .I1(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I2(\u_ras/u_ras_line/r_e2 ),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__1_n_7 ),
        .I4(_inferred__8__0_carry_i_8_n_0),
        .I5(\u_ras/w_err [8]),
        .O(_inferred__8__0_carry__1_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8080000A808AAAA)) 
    _inferred__8__0_carry_i_1
       (.I0(\u_ras/w_e2 [3]),
        .I1(\u_ras/w_err [2]),
        .I2(_inferred__8__0_carry_i_8_n_0),
        .I3(\u_ras/u_ras_line/_inferred__5_carry_n_5 ),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .I5(\u_ras/w_dy [2]),
        .O(_inferred__8__0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD400D4D4D4000000)) 
    _inferred__8__0_carry_i_10
       (.I0(\u_ras/u_ras_line/w_dx ),
        .I1(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I2(\u_ras/u_ras_line/r_e2 ),
        .I3(\u_ras/u_ras_line/_inferred__5_carry_n_4 ),
        .I4(_inferred__8__0_carry_i_8_n_0),
        .I5(\u_ras/w_err [3]),
        .O(_inferred__8__0_carry_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD400D4D4D4000000)) 
    _inferred__8__0_carry_i_11
       (.I0(\u_ras/u_ras_line/w_dx ),
        .I1(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I2(\u_ras/u_ras_line/r_e2 ),
        .I3(\u_ras/u_ras_line/_inferred__5_carry_n_5 ),
        .I4(_inferred__8__0_carry_i_8_n_0),
        .I5(\u_ras/w_err [2]),
        .O(_inferred__8__0_carry_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD400D4D4D4000000)) 
    _inferred__8__0_carry_i_12
       (.I0(\u_ras/u_ras_line/w_dx ),
        .I1(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I2(\u_ras/u_ras_line/r_e2 ),
        .I3(\u_ras/u_ras_line/_inferred__5_carry_n_6 ),
        .I4(_inferred__8__0_carry_i_8_n_0),
        .I5(\u_ras/w_err [1]),
        .O(_inferred__8__0_carry_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8080000A808AAAA)) 
    _inferred__8__0_carry_i_2
       (.I0(\u_ras/w_e2 [2]),
        .I1(\u_ras/w_err [1]),
        .I2(_inferred__8__0_carry_i_8_n_0),
        .I3(\u_ras/u_ras_line/_inferred__5_carry_n_6 ),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .I5(\u_ras/w_dy [1]),
        .O(_inferred__8__0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA808AAAAA808FFFF)) 
    _inferred__8__0_carry_i_3
       (.I0(\u_ras/w_e2 [1]),
        .I1(\u_ras/w_err [0]),
        .I2(_inferred__8__0_carry_i_8_n_0),
        .I3(\u_ras/u_ras_line/_inferred__5_carry_n_7 ),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .I5(\u_ras/w_dy [0]),
        .O(_inferred__8__0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96969669)) 
    _inferred__8__0_carry_i_4
       (.I0(_inferred__8__0_carry_i_1_n_0),
        .I1(_inferred__8__0_carry_i_10_n_0),
        .I2(\u_ras/w_e2 [4]),
        .I3(\u_ras/w_dy [3]),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .O(_inferred__8__0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96969669)) 
    _inferred__8__0_carry_i_5
       (.I0(_inferred__8__0_carry_i_2_n_0),
        .I1(_inferred__8__0_carry_i_11_n_0),
        .I2(\u_ras/w_e2 [3]),
        .I3(\u_ras/w_dy [2]),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .O(_inferred__8__0_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96969669)) 
    _inferred__8__0_carry_i_6
       (.I0(_inferred__8__0_carry_i_3_n_0),
        .I1(_inferred__8__0_carry_i_12_n_0),
        .I2(\u_ras/w_e2 [2]),
        .I3(\u_ras/w_dy [1]),
        .I4(\u_ras/u_ras_line/p_0_in ),
        .O(_inferred__8__0_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h36C6363636C6C6C6)) 
    _inferred__8__0_carry_i_7
       (.I0(\u_ras/w_dy [0]),
        .I1(\u_ras/w_e2 [1]),
        .I2(\u_ras/u_ras_line/p_0_in ),
        .I3(\u_ras/u_ras_line/_inferred__5_carry_n_7 ),
        .I4(_inferred__8__0_carry_i_8_n_0),
        .I5(\u_ras/w_err [0]),
        .O(_inferred__8__0_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h30F5)) 
    _inferred__8__0_carry_i_8
       (.I0(r_x_reg[1]),
        .I1(\u_ras/u_ras_line/result0_carry__0_n_2 ),
        .I2(\u_ras/u_ras_line/r_e2 ),
        .I3(\u_ras/u_ras_line/w_dym__22 ),
        .O(_inferred__8__0_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8E)) 
    _inferred__8__0_carry_i_9
       (.I0(\u_ras/u_ras_line/r_e2 ),
        .I1(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I2(\u_ras/u_ras_line/w_dx ),
        .O(\u_ras/u_ras_line/p_0_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_1
       (.I0(w_v1_y[11]),
        .I1(w_v2_y[11]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_y_tri [11]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/B [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_10
       (.I0(w_v1_y[2]),
        .I1(w_v2_y[2]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_y_tri [2]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/B [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_11
       (.I0(w_v1_y[1]),
        .I1(w_v2_y[1]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_y_tri [1]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/B [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_12
       (.I0(w_v1_y[0]),
        .I1(w_v2_y[0]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_y_tri [0]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/B [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_13
       (.I0(w_v2_x[11]),
        .I1(w_v0_x[11]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_x_tri [11]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/A [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_14
       (.I0(w_v2_x[10]),
        .I1(w_v0_x[10]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_x_tri [10]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/A [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_15
       (.I0(w_v2_x[9]),
        .I1(w_v0_x[9]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_x_tri [9]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/A [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_16
       (.I0(w_v2_x[8]),
        .I1(w_v0_x[8]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_x_tri [8]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/A [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_17
       (.I0(w_v2_x[7]),
        .I1(w_v0_x[7]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_x_tri [7]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/A [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_18
       (.I0(w_v2_x[6]),
        .I1(w_v0_x[6]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_x_tri [6]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/A [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_19
       (.I0(w_v2_x[5]),
        .I1(w_v0_x[5]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_x_tri [5]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/A [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_2
       (.I0(w_v1_y[10]),
        .I1(w_v2_y[10]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_y_tri [10]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/B [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_20
       (.I0(w_v2_x[4]),
        .I1(w_v0_x[4]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_x_tri [4]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/A [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_21
       (.I0(w_v2_x[3]),
        .I1(w_v0_x[3]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_x_tri [3]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/A [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_22
       (.I0(w_v2_x[2]),
        .I1(w_v0_x[2]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_x_tri [2]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/A [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_23
       (.I0(w_v2_x[1]),
        .I1(w_v0_x[1]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_x_tri [1]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/A [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_24
       (.I0(w_v2_x[0]),
        .I1(w_v0_x[0]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_x_tri [0]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/A [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_3
       (.I0(w_v1_y[9]),
        .I1(w_v2_y[9]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_y_tri [9]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/B [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_4
       (.I0(w_v1_y[8]),
        .I1(w_v2_y[8]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_y_tri [8]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/B [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_5
       (.I0(w_v1_y[7]),
        .I1(w_v2_y[7]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_y_tri [7]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/B [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_6
       (.I0(w_v1_y[6]),
        .I1(w_v2_y[6]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_y_tri [6]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/B [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_7
       (.I0(w_v1_y[5]),
        .I1(w_v2_y[5]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_y_tri [5]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/B [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_8
       (.I0(w_v1_y[4]),
        .I1(w_v2_y[4]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_y_tri [4]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/B [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return0_i_9
       (.I0(w_v1_y[3]),
        .I1(w_v2_y[3]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_y_tri [3]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(\u_geo/u_geo_cull/B [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_1
       (.I0(w_v2_y[11]),
        .I1(w_v0_y[11]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_y_tri [11]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_10
       (.I0(w_v2_y[2]),
        .I1(w_v0_y[2]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_y_tri [2]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_11
       (.I0(w_v2_y[1]),
        .I1(w_v0_y[1]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_y_tri [1]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_12
       (.I0(w_v2_y[0]),
        .I1(w_v0_y[0]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_y_tri [0]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_13
       (.I0(w_v1_x[11]),
        .I1(w_v2_x[11]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_x_tri [11]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_14
       (.I0(w_v1_x[10]),
        .I1(w_v2_x[10]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_x_tri [10]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_15
       (.I0(w_v1_x[9]),
        .I1(w_v2_x[9]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_x_tri [9]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_16
       (.I0(w_v1_x[8]),
        .I1(w_v2_x[8]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_x_tri [8]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_17
       (.I0(w_v1_x[7]),
        .I1(w_v2_x[7]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_x_tri [7]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_18
       (.I0(w_v1_x[6]),
        .I1(w_v2_x[6]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_x_tri [6]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_19
       (.I0(w_v1_x[5]),
        .I1(w_v2_x[5]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_x_tri [5]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_2
       (.I0(w_v2_y[10]),
        .I1(w_v0_y[10]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_y_tri [10]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_20
       (.I0(w_v1_x[4]),
        .I1(w_v2_x[4]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_x_tri [4]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_21
       (.I0(w_v1_x[3]),
        .I1(w_v2_x[3]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_x_tri [3]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_22
       (.I0(w_v1_x[2]),
        .I1(w_v2_x[2]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_x_tri [2]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_23
       (.I0(w_v1_x[1]),
        .I1(w_v2_x[1]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_x_tri [1]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_24
       (.I0(w_v1_x[0]),
        .I1(w_v2_x[0]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v0_x_tri [0]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_3
       (.I0(w_v2_y[9]),
        .I1(w_v0_y[9]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_y_tri [9]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_4
       (.I0(w_v2_y[8]),
        .I1(w_v0_y[8]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_y_tri [8]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_5
       (.I0(w_v2_y[7]),
        .I1(w_v0_y[7]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_y_tri [7]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_6
       (.I0(w_v2_y[6]),
        .I1(w_v0_y[6]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_y_tri [6]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_7
       (.I0(w_v2_y[5]),
        .I1(w_v0_y[5]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_y_tri [5]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_8
       (.I0(w_v2_y[4]),
        .I1(w_v0_y[4]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_y_tri [4]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    f_multi_return_i_9
       (.I0(w_v2_y[3]),
        .I1(w_v0_y[3]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/w_v1_y_tri [3]),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .O(f_multi_return_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h66D55B0FC4A9CE58)) 
    g0_b0
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B6663F03C64AB60)) 
    g0_b1
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCBDDD09AA631561E)) 
    g0_b16
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD78D83DFF553BA14)) 
    g0_b17
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9EF9A1311A2B1AD4)) 
    g0_b18
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B04C0A0A1460D90)) 
    g0_b19
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD92D295556B6CC7F)) 
    g0_b2
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6C03AAC06A7EAFB8)) 
    g0_b20
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h700066554C7E6520)) 
    g0_b21
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h80001E33252B49C0)) 
    g0_b22
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAB5A49B38E00)) 
    g0_b23
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99999936DB695AAA)) 
    g0_b24
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h787878F1C718C666)) 
    g0_b25
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF807F80FC0F83E1E)) 
    g0_b26
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h07FFF8003FF801FE)) 
    g0_b27
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF8000007FFFE)) 
    g0_b28
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000007FFFFFFFFFE)) 
    g0_b29
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h38E318CCCD925AD5)) 
    g0_b3
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    g0_b30
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    g0_b31
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h07E0F83C3C71C633)) 
    g0_b4
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFE007FC03F03E0F)) 
    g0_b5
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFE00003FFF001FF)) 
    g0_b6
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFE00000000FFFFF)) 
    g0_b7
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001FFFFFFFFFFFFF)) 
    g0_b8
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g0_b8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h552B5B64C61E003C)) 
    g1_b0
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3366C92DAD4AAAA9)) 
    g1_b1
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4436E2AA54600F59)) 
    g1_b16
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2866412425688770)) 
    g1_b17
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AB9D5DD44CFA8DF)) 
    g1_b18
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h066A99FCD1706560)) 
    g1_b19
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F1E38E39CC66664)) 
    g1_b2
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h01E64B5699801CD5)) 
    g1_b20
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h001E38CDB4AAA966)) 
    g1_b21
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAB5296D9333187)) 
    g1_b22
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6666C9B24B696B52)) 
    g1_b23
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1E1E3871C718E731)) 
    g1_b24
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h01FE07F03F07E0F0)) 
    g1_b25
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001FFF000FFE00F)) 
    g1_b26
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000FFFFFE000)) 
    g1_b27
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000001FFF)) 
    g1_b28
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FE07E07C3E1E1C)) 
    g1_b3
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001FFE003FE01FC)) 
    g1_b4
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000001FFFFE0003)) 
    g1_b5
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000001FFFF)) 
    g1_b6
       (.I0(\u_geo/w_vw_clip [8]),
        .I1(\u_geo/w_vw_clip [9]),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\u_geo/w_vw_clip [11]),
        .I4(\u_geo/w_vw_clip [12]),
        .I5(\u_geo/w_vw_clip [13]),
        .O(g1_b6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[10]_INST_0 
       (.I0(w_adrs_geo[10]),
        .I1(w_adrs_ras[10]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[11]_INST_0 
       (.I0(w_adrs_geo[11]),
        .I1(w_adrs_ras[11]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[12]_INST_0 
       (.I0(w_adrs_geo[12]),
        .I1(w_adrs_ras[12]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[13]_INST_0 
       (.I0(w_adrs_geo[13]),
        .I1(w_adrs_ras[13]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \m_wb_adr_o[13]_INST_0_i_1 
       (.CI(\m_wb_adr_o[9]_INST_0_i_1_n_0 ),
        .CO({\m_wb_adr_o[13]_INST_0_i_1_n_0 ,\m_wb_adr_o[13]_INST_0_i_1_n_1 ,\m_wb_adr_o[13]_INST_0_i_1_n_2 ,\m_wb_adr_o[13]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(w_pixel_top_address[11:8]),
        .O(w_adrs_ras[13:10]),
        .S({\u_ras/u_ras_mem/m_wb_adr_o ,\u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_3_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_4_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[14]_INST_0 
       (.I0(w_adrs_geo[14]),
        .I1(w_adrs_ras[14]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[15]_INST_0 
       (.I0(w_adrs_geo[15]),
        .I1(w_adrs_ras[15]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[16]_INST_0 
       (.I0(w_adrs_geo[16]),
        .I1(w_adrs_ras[16]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[17]_INST_0 
       (.I0(w_adrs_geo[17]),
        .I1(w_adrs_ras[17]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \m_wb_adr_o[17]_INST_0_i_1 
       (.CI(\m_wb_adr_o[13]_INST_0_i_1_n_0 ),
        .CO({\m_wb_adr_o[17]_INST_0_i_1_n_0 ,\m_wb_adr_o[17]_INST_0_i_1_n_1 ,\m_wb_adr_o[17]_INST_0_i_1_n_2 ,\m_wb_adr_o[17]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(w_pixel_top_address[15:12]),
        .O(w_adrs_ras[17:14]),
        .S({\u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_2_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_3_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_4_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[18]_INST_0 
       (.I0(w_adrs_geo[18]),
        .I1(w_adrs_ras[18]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[19]_INST_0 
       (.I0(w_adrs_geo[19]),
        .I1(w_adrs_ras[19]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[20]_INST_0 
       (.I0(w_adrs_geo[20]),
        .I1(w_adrs_ras[20]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[21]_INST_0 
       (.I0(w_adrs_geo[21]),
        .I1(w_adrs_ras[21]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \m_wb_adr_o[21]_INST_0_i_1 
       (.CI(\m_wb_adr_o[17]_INST_0_i_1_n_0 ),
        .CO({\m_wb_adr_o[21]_INST_0_i_1_n_0 ,\m_wb_adr_o[21]_INST_0_i_1_n_1 ,\m_wb_adr_o[21]_INST_0_i_1_n_2 ,\m_wb_adr_o[21]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(w_pixel_top_address[19:16]),
        .O(w_adrs_ras[21:18]),
        .S({\u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_2_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_3_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_4_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[22]_INST_0 
       (.I0(w_adrs_geo[22]),
        .I1(w_adrs_ras[22]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[23]_INST_0 
       (.I0(w_adrs_geo[23]),
        .I1(w_adrs_ras[23]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[24]_INST_0 
       (.I0(w_adrs_geo[24]),
        .I1(w_adrs_ras[24]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[25]_INST_0 
       (.I0(w_adrs_geo[25]),
        .I1(w_adrs_ras[25]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \m_wb_adr_o[25]_INST_0_i_1 
       (.CI(\m_wb_adr_o[21]_INST_0_i_1_n_0 ),
        .CO({\m_wb_adr_o[25]_INST_0_i_1_n_0 ,\m_wb_adr_o[25]_INST_0_i_1_n_1 ,\m_wb_adr_o[25]_INST_0_i_1_n_2 ,\m_wb_adr_o[25]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,w_pixel_top_address[22:20]}),
        .O(w_adrs_ras[25:22]),
        .S({w_pixel_top_address[23],\u_ras/u_ras_mem/m_wb_adr_o[25]_INST_0_i_3_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[25]_INST_0_i_4_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[25]_INST_0_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[26]_INST_0 
       (.I0(w_adrs_geo[26]),
        .I1(w_adrs_ras[26]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[27]_INST_0 
       (.I0(w_adrs_geo[27]),
        .I1(w_adrs_ras[27]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[28]_INST_0 
       (.I0(w_adrs_geo[28]),
        .I1(w_adrs_ras[28]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[29]_INST_0 
       (.I0(w_adrs_geo[29]),
        .I1(w_adrs_ras[29]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \m_wb_adr_o[29]_INST_0_i_1 
       (.CI(\m_wb_adr_o[25]_INST_0_i_1_n_0 ),
        .CO({\m_wb_adr_o[29]_INST_0_i_1_n_0 ,\m_wb_adr_o[29]_INST_0_i_1_n_1 ,\m_wb_adr_o[29]_INST_0_i_1_n_2 ,\m_wb_adr_o[29]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(w_adrs_ras[29:26]),
        .S(w_pixel_top_address[27:24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[2]_INST_0 
       (.I0(w_adrs_geo[2]),
        .I1(w_adrs_ras[2]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[30]_INST_0 
       (.I0(w_adrs_geo[30]),
        .I1(w_adrs_ras[30]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[31]_INST_0 
       (.I0(w_adrs_geo[31]),
        .I1(w_adrs_ras[31]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \m_wb_adr_o[31]_INST_0_i_1 
       (.CI(\m_wb_adr_o[29]_INST_0_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\m_wb_adr_o[31]_INST_0_i_1_n_4 ,\m_wb_adr_o[31]_INST_0_i_1_n_5 ,w_adrs_ras[31:30]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,w_pixel_top_address[29:28]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBBBB8)) 
    \m_wb_adr_o[31]_INST_0_i_2 
       (.I0(\u_mem_arb/r_req_geo ),
        .I1(\u_mem_arb/r_state ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\u_mem_arb/w_pri__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[3]_INST_0 
       (.I0(w_adrs_geo[3]),
        .I1(w_adrs_ras[3]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[4]_INST_0 
       (.I0(w_adrs_geo[4]),
        .I1(w_adrs_ras[4]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[5]_INST_0 
       (.I0(w_adrs_geo[5]),
        .I1(w_adrs_ras[5]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \m_wb_adr_o[5]_INST_0_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\m_wb_adr_o[5]_INST_0_i_1_n_0 ,\m_wb_adr_o[5]_INST_0_i_1_n_1 ,\m_wb_adr_o[5]_INST_0_i_1_n_2 ,\m_wb_adr_o[5]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(w_pixel_top_address[3:0]),
        .O(w_adrs_ras[5:2]),
        .S({\u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_2_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_3_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_4_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[6]_INST_0 
       (.I0(w_adrs_geo[6]),
        .I1(w_adrs_ras[6]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[7]_INST_0 
       (.I0(w_adrs_geo[7]),
        .I1(w_adrs_ras[7]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[8]_INST_0 
       (.I0(w_adrs_geo[8]),
        .I1(w_adrs_ras[8]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \m_wb_adr_o[9]_INST_0 
       (.I0(w_adrs_geo[9]),
        .I1(w_adrs_ras[9]),
        .I2(\u_mem_arb/w_pri__0 ),
        .O(m_wb_adr_o[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \m_wb_adr_o[9]_INST_0_i_1 
       (.CI(\m_wb_adr_o[5]_INST_0_i_1_n_0 ),
        .CO({\m_wb_adr_o[9]_INST_0_i_1_n_0 ,\m_wb_adr_o[9]_INST_0_i_1_n_1 ,\m_wb_adr_o[9]_INST_0_i_1_n_2 ,\m_wb_adr_o[9]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(w_pixel_top_address[7:4]),
        .O(w_adrs_ras[9:6]),
        .S({\u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_2_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_3_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_4_n_0 ,\u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \m_wb_sel_o[1]_INST_0 
       (.I0(\u_ras/u_ras_mem/r_x [0]),
        .I1(\u_ras/u_ras_mem/r_x [1]),
        .O(m_wb_sel_o[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \m_wb_sel_o[2]_INST_0 
       (.I0(\u_ras/u_ras_mem/r_x [1]),
        .I1(\u_ras/u_ras_mem/r_x [0]),
        .O(m_wb_sel_o[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    m_wb_stb_o_INST_0
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I3(\u_ras/u_ras_mem/r_state ),
        .O(m_wb_stb_o));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0001FF01)) 
    m_wb_we_o_INST_0
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I3(\u_mem_arb/r_state ),
        .I4(\u_mem_arb/r_req_geo ),
        .O(m_wb_we_o));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \o_v0_x[11]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [1]),
        .I1(\u_geo/u_geo_cull/r_state [0]),
        .I2(\u_geo/w_en_tri ),
        .O(\u_geo/u_geo_cull/w_set_tri ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h20FF)) 
    r_adrs_m_reg_i_1
       (.I0(\u_ras/w_en_pix ),
        .I1(\u_mem_arb/w_pri__0 ),
        .I2(m_wb_ack_i),
        .I3(\u_ras/u_ras_mem/r_state ),
        .O(r_adrs_m_reg_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    r_adrs_m_reg_i_10
       (.I0(\u_ras/u_ras_mem/w_y0_carry_n_4 ),
        .I1(\u_ras/r_y [3]),
        .I2(w_y_flip),
        .O(\u_ras/B [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    r_adrs_m_reg_i_11
       (.I0(\u_ras/u_ras_mem/w_y0_carry_n_5 ),
        .I1(\u_ras/r_y [2]),
        .I2(w_y_flip),
        .O(\u_ras/B [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    r_adrs_m_reg_i_12
       (.I0(\u_ras/u_ras_mem/w_y0_carry_n_6 ),
        .I1(\u_ras/r_y [1]),
        .I2(w_y_flip),
        .O(\u_ras/B [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    r_adrs_m_reg_i_13
       (.I0(\u_ras/u_ras_mem/w_y0_carry_n_7 ),
        .I1(\u_ras/r_y [0]),
        .I2(w_y_flip),
        .O(\u_ras/B [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    r_adrs_m_reg_i_14
       (.I0(\u_ras/u_ras_line/r_state_reg_n_0_ ),
        .I1(\u_ras/w_y ),
        .I2(\u_ras/u_ras_line/w_reject1__7 ),
        .I3(\u_ras/w_x ),
        .I4(\u_ras/u_ras_line/w_reject0__7 ),
        .I5(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\u_ras/w_en_pix ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    r_adrs_m_reg_i_2
       (.I0(\u_ras/u_ras_mem/w_y0_carry__1_n_4 ),
        .I1(\u_ras/w_y ),
        .I2(w_y_flip),
        .O(\u_ras/B [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    r_adrs_m_reg_i_3
       (.I0(\u_ras/u_ras_mem/w_y0_carry__1_n_5 ),
        .I1(\u_ras/r_y [10]),
        .I2(w_y_flip),
        .O(\u_ras/B [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    r_adrs_m_reg_i_4
       (.I0(\u_ras/u_ras_mem/w_y0_carry__1_n_6 ),
        .I1(\u_ras/r_y [9]),
        .I2(w_y_flip),
        .O(\u_ras/B [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    r_adrs_m_reg_i_5
       (.I0(\u_ras/u_ras_mem/w_y0_carry__1_n_7 ),
        .I1(\u_ras/r_y [8]),
        .I2(w_y_flip),
        .O(\u_ras/B [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    r_adrs_m_reg_i_6
       (.I0(\u_ras/u_ras_mem/w_y0_carry__0_n_4 ),
        .I1(\u_ras/r_y [7]),
        .I2(w_y_flip),
        .O(\u_ras/B [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    r_adrs_m_reg_i_7
       (.I0(\u_ras/u_ras_mem/w_y0_carry__0_n_5 ),
        .I1(\u_ras/r_y [6]),
        .I2(w_y_flip),
        .O(\u_ras/B [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    r_adrs_m_reg_i_8
       (.I0(\u_ras/u_ras_mem/w_y0_carry__0_n_6 ),
        .I1(\u_ras/r_y [5]),
        .I2(w_y_flip),
        .O(\u_ras/B [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    r_adrs_m_reg_i_9
       (.I0(\u_ras/u_ras_mem/w_y0_carry__0_n_7 ),
        .I1(\u_ras/r_y [4]),
        .I2(w_y_flip),
        .O(\u_ras/B [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_bc[0]_i_1 
       (.I0(\u_geo/u_geo_clip/p_0_in0 ),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I2(\u_geo/w_outcode_clip [0]),
        .O(r_bc));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_bc[1]_i_1 
       (.I0(\u_geo/u_geo_clip/p_0_in0 ),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/w_outcode_clip [1]),
        .O(\r_bc[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_bc[2]_i_1 
       (.I0(\u_geo/u_geo_clip/p_0_in0 ),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I2(\u_geo/w_outcode_clip [2]),
        .O(\r_bc[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_bc[3]_i_1 
       (.I0(\u_geo/u_geo_clip/p_0_in0 ),
        .I1(\u_geo/u_geo_clip/r_bc ),
        .I2(\u_geo/w_outcode_clip [3]),
        .O(\r_bc[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_bc[4]_i_1 
       (.I0(\u_geo/u_geo_clip/p_0_in0 ),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[7] ),
        .I2(\u_geo/w_outcode_clip [4]),
        .O(\r_bc[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_bc[5]_i_1 
       (.I0(\u_geo/u_geo_clip/p_0_in0 ),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[8] ),
        .I2(\u_geo/w_outcode_clip [5]),
        .O(\r_bc[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FE00)) 
    \r_c[0]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[17]_i_2_n_0 ),
        .I4(\r_c[0]_i_2_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACA0)) 
    \r_c[0]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [1]),
        .I1(\r_c[0]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I3(\r_c[14]_i_4_n_0 ),
        .O(r_c));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACA0)) 
    \r_c[0]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [1]),
        .I1(\r_c[0]_i_2__3_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I3(\r_c[14]_i_4__0_n_0 ),
        .O(\r_c[0]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACA0)) 
    \r_c[0]_i_1__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [1]),
        .I1(\r_c[0]_i_2__4_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I3(\r_c[14]_i_4__1_n_0 ),
        .O(\r_c[0]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACA0)) 
    \r_c[0]_i_1__3 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [1]),
        .I1(\r_c[0]_i_2__5_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I3(\r_c[14]_i_4__2_n_0 ),
        .O(\r_c[0]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACA0)) 
    \r_c[0]_i_1__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [1]),
        .I1(\r_c[0]_i_2__6_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I3(\r_c[14]_i_4__3_n_0 ),
        .O(\r_c[0]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACA0)) 
    \r_c[0]_i_1__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [1]),
        .I1(\r_c[0]_i_2__7_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I3(\r_c[14]_i_4__4_n_0 ),
        .O(\r_c[0]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACA0)) 
    \r_c[0]_i_1__6 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [1]),
        .I1(\r_c[0]_i_2__8_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I3(\r_c[14]_i_4__5_n_0 ),
        .O(\r_c[0]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA0E4)) 
    \r_c[0]_i_1__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I1(\r_c[14]_i_4__7_n_0 ),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [1]),
        .I3(\r_c[0]_i_2__0_n_0 ),
        .O(\r_c[0]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA0E4)) 
    \r_c[0]_i_1__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I1(\r_c[14]_i_4__8_n_0 ),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [1]),
        .I3(\r_c[0]_i_2__1_n_0 ),
        .O(\r_c[0]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    \r_c[0]_i_2 
       (.I0(\r_c[17]_i_3_n_0 ),
        .I1(\r_c[20]_i_2__6_n_0 ),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [0]),
        .I3(\r_c[18]_i_3_n_0 ),
        .O(\r_c[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFBF)) 
    \r_c[0]_i_2__0 
       (.I0(\r_c[1]_i_3__6_n_0 ),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [0]),
        .I2(_inferred__1_carry_i_6__7_n_0),
        .I3(_inferred__1_carry_i_7__7_n_0),
        .O(\r_c[0]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFBF)) 
    \r_c[0]_i_2__1 
       (.I0(\r_c[1]_i_3__7_n_0 ),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [0]),
        .I2(_inferred__1_carry_i_6__9_n_0),
        .I3(_inferred__1_carry_i_7__9_n_0),
        .O(\r_c[0]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[0]_i_2__2 
       (.I0(\r_c[1]_i_3_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [0]),
        .I2(_inferred__1_carry_i_6_n_0),
        .I3(_inferred__1_carry_i_7_n_0),
        .O(\r_c[0]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[0]_i_2__3 
       (.I0(\r_c[1]_i_3__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [0]),
        .I2(_inferred__1_carry_i_6__0_n_0),
        .I3(_inferred__1_carry_i_7__0_n_0),
        .O(\r_c[0]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[0]_i_2__4 
       (.I0(\r_c[1]_i_3__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [0]),
        .I2(_inferred__1_carry_i_6__1_n_0),
        .I3(_inferred__1_carry_i_7__1_n_0),
        .O(\r_c[0]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[0]_i_2__5 
       (.I0(\r_c[1]_i_3__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [0]),
        .I2(_inferred__1_carry_i_6__2_n_0),
        .I3(_inferred__1_carry_i_7__2_n_0),
        .O(\r_c[0]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[0]_i_2__6 
       (.I0(\r_c[1]_i_3__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [0]),
        .I2(_inferred__1_carry_i_6__3_n_0),
        .I3(_inferred__1_carry_i_7__3_n_0),
        .O(\r_c[0]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[0]_i_2__7 
       (.I0(\r_c[1]_i_3__4_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [0]),
        .I2(_inferred__1_carry_i_6__4_n_0),
        .I3(_inferred__1_carry_i_7__4_n_0),
        .O(\r_c[0]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[0]_i_2__8 
       (.I0(\r_c[1]_i_3__5_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [0]),
        .I2(_inferred__1_carry_i_6__5_n_0),
        .I3(_inferred__1_carry_i_7__5_n_0),
        .O(\r_c[0]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[10]_i_1 
       (.I0(\r_c[10]_i_2_n_0 ),
        .I1(\r_c[14]_i_4_n_0 ),
        .I2(\r_c[11]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [11]),
        .O(\r_c[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[10]_i_1__0 
       (.I0(\r_c[10]_i_2__0_n_0 ),
        .I1(\r_c[14]_i_4__0_n_0 ),
        .I2(\r_c[11]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [11]),
        .O(\r_c[10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[10]_i_1__1 
       (.I0(\r_c[10]_i_2__1_n_0 ),
        .I1(\r_c[14]_i_4__1_n_0 ),
        .I2(\r_c[11]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [11]),
        .O(\r_c[10]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[10]_i_1__2 
       (.I0(\r_c[10]_i_2__2_n_0 ),
        .I1(\r_c[14]_i_4__2_n_0 ),
        .I2(\r_c[11]_i_2__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [11]),
        .O(\r_c[10]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[10]_i_1__3 
       (.I0(\r_c[10]_i_2__3_n_0 ),
        .I1(\r_c[14]_i_4__3_n_0 ),
        .I2(\r_c[11]_i_2__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [11]),
        .O(\r_c[10]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[10]_i_1__4 
       (.I0(\r_c[10]_i_2__4_n_0 ),
        .I1(\r_c[14]_i_4__4_n_0 ),
        .I2(\r_c[11]_i_2__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [11]),
        .O(\r_c[10]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[10]_i_1__5 
       (.I0(\r_c[10]_i_2__5_n_0 ),
        .I1(\r_c[14]_i_4__5_n_0 ),
        .I2(\r_c[11]_i_2__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [11]),
        .O(\r_c[10]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[10]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[10]_i_2__6_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[11]_i_2__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCC55)) 
    \r_c[10]_i_1__7 
       (.I0(\r_c[10]_i_2__7_n_0 ),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [11]),
        .I2(\r_c[11]_i_2__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\r_c[14]_i_4__7_n_0 ),
        .O(\r_c[10]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCC55)) 
    \r_c[10]_i_1__8 
       (.I0(\r_c[10]_i_2__8_n_0 ),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [11]),
        .I2(\r_c[11]_i_2__8_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\r_c[14]_i_4__8_n_0 ),
        .O(\r_c[10]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[10]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [3]),
        .I1(_inferred__1_carry_i_7_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [7]),
        .I3(_inferred__1_carry_i_6_n_0),
        .I4(\r_c[1]_i_3_n_0 ),
        .I5(\r_c[12]_i_3_n_0 ),
        .O(\r_c[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[10]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [3]),
        .I1(_inferred__1_carry_i_7__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [7]),
        .I3(_inferred__1_carry_i_6__0_n_0),
        .I4(\r_c[1]_i_3__0_n_0 ),
        .I5(\r_c[12]_i_3__0_n_0 ),
        .O(\r_c[10]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[10]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [3]),
        .I1(_inferred__1_carry_i_7__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [7]),
        .I3(_inferred__1_carry_i_6__1_n_0),
        .I4(\r_c[1]_i_3__1_n_0 ),
        .I5(\r_c[12]_i_3__1_n_0 ),
        .O(\r_c[10]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[10]_i_2__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [3]),
        .I1(_inferred__1_carry_i_7__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [7]),
        .I3(_inferred__1_carry_i_6__2_n_0),
        .I4(\r_c[1]_i_3__2_n_0 ),
        .I5(\r_c[12]_i_3__2_n_0 ),
        .O(\r_c[10]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[10]_i_2__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [3]),
        .I1(_inferred__1_carry_i_7__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [7]),
        .I3(_inferred__1_carry_i_6__3_n_0),
        .I4(\r_c[1]_i_3__3_n_0 ),
        .I5(\r_c[12]_i_3__3_n_0 ),
        .O(\r_c[10]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[10]_i_2__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [3]),
        .I1(_inferred__1_carry_i_7__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [7]),
        .I3(_inferred__1_carry_i_6__4_n_0),
        .I4(\r_c[1]_i_3__4_n_0 ),
        .I5(\r_c[12]_i_3__4_n_0 ),
        .O(\r_c[10]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[10]_i_2__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [3]),
        .I1(_inferred__1_carry_i_7__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [7]),
        .I3(_inferred__1_carry_i_6__5_n_0),
        .I4(\r_c[1]_i_3__5_n_0 ),
        .I5(\r_c[12]_i_3__5_n_0 ),
        .O(\r_c[10]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \r_c[10]_i_2__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [3]),
        .I1(\r_c[18]_i_3_n_0 ),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [7]),
        .I4(\r_c[17]_i_3_n_0 ),
        .I5(\r_c[12]_i_3__6_n_0 ),
        .O(\r_c[10]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[10]_i_2__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [3]),
        .I1(_inferred__1_carry_i_7__7_n_0),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [7]),
        .I3(_inferred__1_carry_i_6__7_n_0),
        .I4(\r_c[1]_i_3__6_n_0 ),
        .I5(\r_c[12]_i_3__7_n_0 ),
        .O(\r_c[10]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[10]_i_2__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [3]),
        .I1(_inferred__1_carry_i_7__9_n_0),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [7]),
        .I3(_inferred__1_carry_i_6__9_n_0),
        .I4(\r_c[1]_i_3__7_n_0 ),
        .I5(\r_c[12]_i_3__8_n_0 ),
        .O(\r_c[10]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[11]_i_1 
       (.I0(\r_c[11]_i_2_n_0 ),
        .I1(\r_c[14]_i_4_n_0 ),
        .I2(\r_c[12]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [12]),
        .O(\r_c[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[11]_i_1__0 
       (.I0(\r_c[11]_i_2__0_n_0 ),
        .I1(\r_c[14]_i_4__0_n_0 ),
        .I2(\r_c[12]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [12]),
        .O(\r_c[11]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[11]_i_1__1 
       (.I0(\r_c[11]_i_2__1_n_0 ),
        .I1(\r_c[14]_i_4__1_n_0 ),
        .I2(\r_c[12]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [12]),
        .O(\r_c[11]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[11]_i_1__2 
       (.I0(\r_c[11]_i_2__2_n_0 ),
        .I1(\r_c[14]_i_4__2_n_0 ),
        .I2(\r_c[12]_i_2__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [12]),
        .O(\r_c[11]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[11]_i_1__3 
       (.I0(\r_c[11]_i_2__3_n_0 ),
        .I1(\r_c[14]_i_4__3_n_0 ),
        .I2(\r_c[12]_i_2__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [12]),
        .O(\r_c[11]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[11]_i_1__4 
       (.I0(\r_c[11]_i_2__4_n_0 ),
        .I1(\r_c[14]_i_4__4_n_0 ),
        .I2(\r_c[12]_i_2__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [12]),
        .O(\r_c[11]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[11]_i_1__5 
       (.I0(\r_c[11]_i_2__5_n_0 ),
        .I1(\r_c[14]_i_4__5_n_0 ),
        .I2(\r_c[12]_i_2__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [12]),
        .O(\r_c[11]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[11]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[11]_i_2__6_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[12]_i_2__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[11]_i_1__7 
       (.I0(\r_c[11]_i_2__7_n_0 ),
        .I1(\r_c[14]_i_4__7_n_0 ),
        .I2(\r_c[12]_i_2__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [12]),
        .O(\r_c[11]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[11]_i_1__8 
       (.I0(\r_c[11]_i_2__8_n_0 ),
        .I1(\r_c[14]_i_4__8_n_0 ),
        .I2(\r_c[12]_i_2__8_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [12]),
        .O(\r_c[11]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[11]_i_2 
       (.I0(\r_c[11]_i_3_n_0 ),
        .I1(\r_c[1]_i_3_n_0 ),
        .I2(\r_c[13]_i_3_n_0 ),
        .O(\r_c[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[11]_i_2__0 
       (.I0(\r_c[11]_i_3__0_n_0 ),
        .I1(\r_c[1]_i_3__0_n_0 ),
        .I2(\r_c[13]_i_3__0_n_0 ),
        .O(\r_c[11]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[11]_i_2__1 
       (.I0(\r_c[11]_i_3__1_n_0 ),
        .I1(\r_c[1]_i_3__1_n_0 ),
        .I2(\r_c[13]_i_3__1_n_0 ),
        .O(\r_c[11]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[11]_i_2__2 
       (.I0(\r_c[11]_i_3__2_n_0 ),
        .I1(\r_c[1]_i_3__2_n_0 ),
        .I2(\r_c[13]_i_3__2_n_0 ),
        .O(\r_c[11]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[11]_i_2__3 
       (.I0(\r_c[11]_i_3__3_n_0 ),
        .I1(\r_c[1]_i_3__3_n_0 ),
        .I2(\r_c[13]_i_3__3_n_0 ),
        .O(\r_c[11]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[11]_i_2__4 
       (.I0(\r_c[11]_i_3__4_n_0 ),
        .I1(\r_c[1]_i_3__4_n_0 ),
        .I2(\r_c[13]_i_3__4_n_0 ),
        .O(\r_c[11]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[11]_i_2__5 
       (.I0(\r_c[11]_i_3__5_n_0 ),
        .I1(\r_c[1]_i_3__5_n_0 ),
        .I2(\r_c[13]_i_3__5_n_0 ),
        .O(\r_c[11]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[11]_i_2__6 
       (.I0(\r_c[11]_i_3__6_n_0 ),
        .I1(\r_c[17]_i_3_n_0 ),
        .I2(\r_c[13]_i_3__6_n_0 ),
        .O(\r_c[11]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[11]_i_2__7 
       (.I0(\r_c[11]_i_3__7_n_0 ),
        .I1(\r_c[1]_i_3__6_n_0 ),
        .I2(\r_c[13]_i_3__7_n_0 ),
        .O(\r_c[11]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[11]_i_2__8 
       (.I0(\r_c[11]_i_3__8_n_0 ),
        .I1(\r_c[1]_i_3__7_n_0 ),
        .I2(\r_c[13]_i_3__8_n_0 ),
        .O(\r_c[11]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[11]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [4]),
        .I1(_inferred__1_carry_i_7_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [8]),
        .I3(_inferred__1_carry_i_6_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [0]),
        .O(\r_c[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[11]_i_3__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [4]),
        .I1(_inferred__1_carry_i_7__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [8]),
        .I3(_inferred__1_carry_i_6__0_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [0]),
        .O(\r_c[11]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[11]_i_3__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [4]),
        .I1(_inferred__1_carry_i_7__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [8]),
        .I3(_inferred__1_carry_i_6__1_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [0]),
        .O(\r_c[11]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[11]_i_3__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [4]),
        .I1(_inferred__1_carry_i_7__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [8]),
        .I3(_inferred__1_carry_i_6__2_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [0]),
        .O(\r_c[11]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[11]_i_3__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [4]),
        .I1(_inferred__1_carry_i_7__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [8]),
        .I3(_inferred__1_carry_i_6__3_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [0]),
        .O(\r_c[11]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[11]_i_3__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [4]),
        .I1(_inferred__1_carry_i_7__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [8]),
        .I3(_inferred__1_carry_i_6__4_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [0]),
        .O(\r_c[11]_i_3__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[11]_i_3__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [4]),
        .I1(_inferred__1_carry_i_7__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [8]),
        .I3(_inferred__1_carry_i_6__5_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [0]),
        .O(\r_c[11]_i_3__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC4C4C7F7)) 
    \r_c[11]_i_3__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [4]),
        .I1(\r_c[18]_i_3_n_0 ),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [0]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [8]),
        .O(\r_c[11]_i_3__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[11]_i_3__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [4]),
        .I1(_inferred__1_carry_i_7__7_n_0),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [8]),
        .I3(_inferred__1_carry_i_6__7_n_0),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [0]),
        .O(\r_c[11]_i_3__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[11]_i_3__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [4]),
        .I1(_inferred__1_carry_i_7__9_n_0),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [8]),
        .I3(_inferred__1_carry_i_6__9_n_0),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [0]),
        .O(\r_c[11]_i_3__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[12]_i_1 
       (.I0(\r_c[12]_i_2_n_0 ),
        .I1(\r_c[14]_i_4_n_0 ),
        .I2(\r_c[13]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [13]),
        .O(\r_c[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[12]_i_1__0 
       (.I0(\r_c[12]_i_2__0_n_0 ),
        .I1(\r_c[14]_i_4__0_n_0 ),
        .I2(\r_c[13]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [13]),
        .O(\r_c[12]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[12]_i_1__1 
       (.I0(\r_c[12]_i_2__1_n_0 ),
        .I1(\r_c[14]_i_4__1_n_0 ),
        .I2(\r_c[13]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [13]),
        .O(\r_c[12]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[12]_i_1__2 
       (.I0(\r_c[12]_i_2__2_n_0 ),
        .I1(\r_c[14]_i_4__2_n_0 ),
        .I2(\r_c[13]_i_2__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [13]),
        .O(\r_c[12]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[12]_i_1__3 
       (.I0(\r_c[12]_i_2__3_n_0 ),
        .I1(\r_c[14]_i_4__3_n_0 ),
        .I2(\r_c[13]_i_2__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [13]),
        .O(\r_c[12]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[12]_i_1__4 
       (.I0(\r_c[12]_i_2__4_n_0 ),
        .I1(\r_c[14]_i_4__4_n_0 ),
        .I2(\r_c[13]_i_2__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [13]),
        .O(\r_c[12]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[12]_i_1__5 
       (.I0(\r_c[12]_i_2__5_n_0 ),
        .I1(\r_c[14]_i_4__5_n_0 ),
        .I2(\r_c[13]_i_2__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [13]),
        .O(\r_c[12]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[12]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[12]_i_2__6_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[13]_i_2__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[12]_i_1__7 
       (.I0(\r_c[12]_i_2__7_n_0 ),
        .I1(\r_c[14]_i_4__7_n_0 ),
        .I2(\r_c[13]_i_2__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [13]),
        .O(\r_c[12]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[12]_i_1__8 
       (.I0(\r_c[12]_i_2__8_n_0 ),
        .I1(\r_c[14]_i_4__8_n_0 ),
        .I2(\r_c[13]_i_2__8_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [13]),
        .O(\r_c[12]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[12]_i_2 
       (.I0(\r_c[12]_i_3_n_0 ),
        .I1(\r_c[1]_i_3_n_0 ),
        .I2(\r_c[14]_i_5_n_0 ),
        .O(\r_c[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[12]_i_2__0 
       (.I0(\r_c[12]_i_3__0_n_0 ),
        .I1(\r_c[1]_i_3__0_n_0 ),
        .I2(\r_c[14]_i_5__0_n_0 ),
        .O(\r_c[12]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[12]_i_2__1 
       (.I0(\r_c[12]_i_3__1_n_0 ),
        .I1(\r_c[1]_i_3__1_n_0 ),
        .I2(\r_c[14]_i_5__1_n_0 ),
        .O(\r_c[12]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[12]_i_2__2 
       (.I0(\r_c[12]_i_3__2_n_0 ),
        .I1(\r_c[1]_i_3__2_n_0 ),
        .I2(\r_c[14]_i_5__2_n_0 ),
        .O(\r_c[12]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[12]_i_2__3 
       (.I0(\r_c[12]_i_3__3_n_0 ),
        .I1(\r_c[1]_i_3__3_n_0 ),
        .I2(\r_c[14]_i_5__3_n_0 ),
        .O(\r_c[12]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[12]_i_2__4 
       (.I0(\r_c[12]_i_3__4_n_0 ),
        .I1(\r_c[1]_i_3__4_n_0 ),
        .I2(\r_c[14]_i_5__4_n_0 ),
        .O(\r_c[12]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[12]_i_2__5 
       (.I0(\r_c[12]_i_3__5_n_0 ),
        .I1(\r_c[1]_i_3__5_n_0 ),
        .I2(\r_c[14]_i_5__5_n_0 ),
        .O(\r_c[12]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[12]_i_2__6 
       (.I0(\r_c[12]_i_3__6_n_0 ),
        .I1(\r_c[17]_i_3_n_0 ),
        .I2(\r_c[14]_i_7__6_n_0 ),
        .O(\r_c[12]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[12]_i_2__7 
       (.I0(\r_c[12]_i_3__7_n_0 ),
        .I1(\r_c[1]_i_3__6_n_0 ),
        .I2(\r_c[14]_i_5__7_n_0 ),
        .O(\r_c[12]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[12]_i_2__8 
       (.I0(\r_c[12]_i_3__8_n_0 ),
        .I1(\r_c[1]_i_3__7_n_0 ),
        .I2(\r_c[14]_i_5__8_n_0 ),
        .O(\r_c[12]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[12]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [5]),
        .I1(_inferred__1_carry_i_7_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [9]),
        .I3(_inferred__1_carry_i_6_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [1]),
        .O(\r_c[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[12]_i_3__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [5]),
        .I1(_inferred__1_carry_i_7__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [9]),
        .I3(_inferred__1_carry_i_6__0_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [1]),
        .O(\r_c[12]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[12]_i_3__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [5]),
        .I1(_inferred__1_carry_i_7__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [9]),
        .I3(_inferred__1_carry_i_6__1_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [1]),
        .O(\r_c[12]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[12]_i_3__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [5]),
        .I1(_inferred__1_carry_i_7__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [9]),
        .I3(_inferred__1_carry_i_6__2_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [1]),
        .O(\r_c[12]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[12]_i_3__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [5]),
        .I1(_inferred__1_carry_i_7__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [9]),
        .I3(_inferred__1_carry_i_6__3_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [1]),
        .O(\r_c[12]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[12]_i_3__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [5]),
        .I1(_inferred__1_carry_i_7__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [9]),
        .I3(_inferred__1_carry_i_6__4_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [1]),
        .O(\r_c[12]_i_3__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[12]_i_3__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [5]),
        .I1(_inferred__1_carry_i_7__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [9]),
        .I3(_inferred__1_carry_i_6__5_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [1]),
        .O(\r_c[12]_i_3__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC4C4C7F7)) 
    \r_c[12]_i_3__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [5]),
        .I1(\r_c[18]_i_3_n_0 ),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [1]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [9]),
        .O(\r_c[12]_i_3__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[12]_i_3__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [5]),
        .I1(_inferred__1_carry_i_7__7_n_0),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [9]),
        .I3(_inferred__1_carry_i_6__7_n_0),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [1]),
        .O(\r_c[12]_i_3__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[12]_i_3__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [5]),
        .I1(_inferred__1_carry_i_7__9_n_0),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [9]),
        .I3(_inferred__1_carry_i_6__9_n_0),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [1]),
        .O(\r_c[12]_i_3__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[13]_i_1 
       (.I0(\r_c[13]_i_2_n_0 ),
        .I1(\r_c[14]_i_4_n_0 ),
        .I2(\r_c[14]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [14]),
        .O(\r_c[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[13]_i_1__0 
       (.I0(\r_c[13]_i_2__0_n_0 ),
        .I1(\r_c[14]_i_4__0_n_0 ),
        .I2(\r_c[14]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [14]),
        .O(\r_c[13]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[13]_i_1__1 
       (.I0(\r_c[13]_i_2__1_n_0 ),
        .I1(\r_c[14]_i_4__1_n_0 ),
        .I2(\r_c[14]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [14]),
        .O(\r_c[13]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[13]_i_1__2 
       (.I0(\r_c[13]_i_2__2_n_0 ),
        .I1(\r_c[14]_i_4__2_n_0 ),
        .I2(\r_c[14]_i_2__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [14]),
        .O(\r_c[13]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[13]_i_1__3 
       (.I0(\r_c[13]_i_2__3_n_0 ),
        .I1(\r_c[14]_i_4__3_n_0 ),
        .I2(\r_c[14]_i_2__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [14]),
        .O(\r_c[13]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[13]_i_1__4 
       (.I0(\r_c[13]_i_2__4_n_0 ),
        .I1(\r_c[14]_i_4__4_n_0 ),
        .I2(\r_c[14]_i_2__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [14]),
        .O(\r_c[13]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[13]_i_1__5 
       (.I0(\r_c[13]_i_2__5_n_0 ),
        .I1(\r_c[14]_i_4__5_n_0 ),
        .I2(\r_c[14]_i_2__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [14]),
        .O(\r_c[13]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[13]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[13]_i_2__6_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[14]_i_3__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[13]_i_1__7 
       (.I0(\r_c[13]_i_2__7_n_0 ),
        .I1(\r_c[14]_i_4__7_n_0 ),
        .I2(\r_c[14]_i_2__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [14]),
        .O(\r_c[13]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[13]_i_1__8 
       (.I0(\r_c[13]_i_2__8_n_0 ),
        .I1(\r_c[14]_i_4__8_n_0 ),
        .I2(\r_c[14]_i_2__8_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [14]),
        .O(\r_c[13]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[13]_i_2 
       (.I0(\r_c[13]_i_3_n_0 ),
        .I1(\r_c[1]_i_3_n_0 ),
        .I2(\r_c[14]_i_8_n_0 ),
        .O(\r_c[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[13]_i_2__0 
       (.I0(\r_c[13]_i_3__0_n_0 ),
        .I1(\r_c[1]_i_3__0_n_0 ),
        .I2(\r_c[14]_i_8__0_n_0 ),
        .O(\r_c[13]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[13]_i_2__1 
       (.I0(\r_c[13]_i_3__1_n_0 ),
        .I1(\r_c[1]_i_3__1_n_0 ),
        .I2(\r_c[14]_i_8__1_n_0 ),
        .O(\r_c[13]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[13]_i_2__2 
       (.I0(\r_c[13]_i_3__2_n_0 ),
        .I1(\r_c[1]_i_3__2_n_0 ),
        .I2(\r_c[14]_i_8__2_n_0 ),
        .O(\r_c[13]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[13]_i_2__3 
       (.I0(\r_c[13]_i_3__3_n_0 ),
        .I1(\r_c[1]_i_3__3_n_0 ),
        .I2(\r_c[14]_i_8__3_n_0 ),
        .O(\r_c[13]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[13]_i_2__4 
       (.I0(\r_c[13]_i_3__4_n_0 ),
        .I1(\r_c[1]_i_3__4_n_0 ),
        .I2(\r_c[14]_i_8__4_n_0 ),
        .O(\r_c[13]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[13]_i_2__5 
       (.I0(\r_c[13]_i_3__5_n_0 ),
        .I1(\r_c[1]_i_3__5_n_0 ),
        .I2(\r_c[14]_i_8__5_n_0 ),
        .O(\r_c[13]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[13]_i_2__6 
       (.I0(\r_c[13]_i_3__6_n_0 ),
        .I1(\r_c[17]_i_3_n_0 ),
        .I2(\r_c[20]_i_6_n_0 ),
        .O(\r_c[13]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[13]_i_2__7 
       (.I0(\r_c[13]_i_3__7_n_0 ),
        .I1(\r_c[1]_i_3__6_n_0 ),
        .I2(\r_c[14]_i_8__7_n_0 ),
        .O(\r_c[13]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[13]_i_2__8 
       (.I0(\r_c[13]_i_3__8_n_0 ),
        .I1(\r_c[1]_i_3__7_n_0 ),
        .I2(\r_c[14]_i_8__8_n_0 ),
        .O(\r_c[13]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[13]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [6]),
        .I1(_inferred__1_carry_i_7_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [10]),
        .I3(_inferred__1_carry_i_6_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [2]),
        .O(\r_c[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[13]_i_3__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [6]),
        .I1(_inferred__1_carry_i_7__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [10]),
        .I3(_inferred__1_carry_i_6__0_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [2]),
        .O(\r_c[13]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[13]_i_3__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [6]),
        .I1(_inferred__1_carry_i_7__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [10]),
        .I3(_inferred__1_carry_i_6__1_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [2]),
        .O(\r_c[13]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[13]_i_3__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [6]),
        .I1(_inferred__1_carry_i_7__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [10]),
        .I3(_inferred__1_carry_i_6__2_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [2]),
        .O(\r_c[13]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[13]_i_3__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [6]),
        .I1(_inferred__1_carry_i_7__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [10]),
        .I3(_inferred__1_carry_i_6__3_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [2]),
        .O(\r_c[13]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[13]_i_3__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [6]),
        .I1(_inferred__1_carry_i_7__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [10]),
        .I3(_inferred__1_carry_i_6__4_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [2]),
        .O(\r_c[13]_i_3__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[13]_i_3__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [6]),
        .I1(_inferred__1_carry_i_7__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [10]),
        .I3(_inferred__1_carry_i_6__5_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [2]),
        .O(\r_c[13]_i_3__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC4C4C7F7)) 
    \r_c[13]_i_3__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [6]),
        .I1(\r_c[18]_i_3_n_0 ),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [2]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [10]),
        .O(\r_c[13]_i_3__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[13]_i_3__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [6]),
        .I1(_inferred__1_carry_i_7__7_n_0),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [10]),
        .I3(_inferred__1_carry_i_6__7_n_0),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [2]),
        .O(\r_c[13]_i_3__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[13]_i_3__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [6]),
        .I1(_inferred__1_carry_i_7__9_n_0),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [10]),
        .I3(_inferred__1_carry_i_6__9_n_0),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [2]),
        .O(\r_c[13]_i_3__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[14]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[14]_i_3__6_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[14]_i_4__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00F4)) 
    \r_c[14]_i_10 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [11]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [13]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [14]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [15]),
        .O(\r_c[14]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00F4)) 
    \r_c[14]_i_10__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [11]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [13]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [14]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [15]),
        .O(\r_c[14]_i_10__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00F4)) 
    \r_c[14]_i_10__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [11]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [13]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [14]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [15]),
        .O(\r_c[14]_i_10__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00F4)) 
    \r_c[14]_i_10__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [11]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [13]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [14]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [15]),
        .O(\r_c[14]_i_10__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00F4)) 
    \r_c[14]_i_10__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [12]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [11]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [13]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [14]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [15]),
        .O(\r_c[14]_i_10__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00F4)) 
    \r_c[14]_i_10__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [12]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [11]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [13]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [14]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [15]),
        .O(\r_c[14]_i_10__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00F4)) 
    \r_c[14]_i_10__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [12]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [11]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [13]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [14]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [15]),
        .O(\r_c[14]_i_10__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00F4)) 
    \r_c[14]_i_10__6 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [11]),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [13]),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [14]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [15]),
        .O(\r_c[14]_i_10__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00F4)) 
    \r_c[14]_i_10__7 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [12]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [11]),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [13]),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [14]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [15]),
        .O(\r_c[14]_i_10__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r_c[14]_i_11 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [8]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [12]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [14]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [10]),
        .O(\r_c[14]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r_c[14]_i_11__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [8]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [12]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [14]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [10]),
        .O(\r_c[14]_i_11__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r_c[14]_i_11__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [8]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [12]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [14]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [10]),
        .O(\r_c[14]_i_11__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r_c[14]_i_11__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [8]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [12]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [14]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [10]),
        .O(\r_c[14]_i_11__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r_c[14]_i_11__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [8]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [12]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [14]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [10]),
        .O(\r_c[14]_i_11__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r_c[14]_i_11__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [8]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [12]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [14]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [10]),
        .O(\r_c[14]_i_11__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r_c[14]_i_11__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [8]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [12]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [14]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [10]),
        .O(\r_c[14]_i_11__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r_c[14]_i_11__6 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [8]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [12]),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [14]),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [10]),
        .O(\r_c[14]_i_11__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r_c[14]_i_11__7 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [8]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [12]),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [14]),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [10]),
        .O(\r_c[14]_i_11__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551011)) 
    \r_c[14]_i_12 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [5]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [3]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [2]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [1]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [4]),
        .O(\r_c[14]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551011)) 
    \r_c[14]_i_12__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [5]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [3]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [2]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [1]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [4]),
        .O(\r_c[14]_i_12__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551011)) 
    \r_c[14]_i_12__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [5]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [3]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [2]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [1]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [4]),
        .O(\r_c[14]_i_12__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551011)) 
    \r_c[14]_i_12__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [5]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [3]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [2]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [1]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [4]),
        .O(\r_c[14]_i_12__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551011)) 
    \r_c[14]_i_12__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [5]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [3]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [2]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [1]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [4]),
        .O(\r_c[14]_i_12__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551011)) 
    \r_c[14]_i_12__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [5]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [3]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [2]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [1]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [4]),
        .O(\r_c[14]_i_12__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551011)) 
    \r_c[14]_i_12__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [5]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [3]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [2]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [1]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [4]),
        .O(\r_c[14]_i_12__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551011)) 
    \r_c[14]_i_12__6 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [5]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [3]),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [2]),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [1]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [4]),
        .O(\r_c[14]_i_12__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551011)) 
    \r_c[14]_i_12__7 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [5]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [3]),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [2]),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [1]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [4]),
        .O(\r_c[14]_i_12__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCC55)) 
    \r_c[14]_i_1__0 
       (.I0(\r_c[14]_i_2_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [15]),
        .I2(\r_c[14]_i_3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I4(\r_c[14]_i_4_n_0 ),
        .O(\r_c[14]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCC55)) 
    \r_c[14]_i_1__1 
       (.I0(\r_c[14]_i_2__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [15]),
        .I2(\r_c[14]_i_3__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I4(\r_c[14]_i_4__0_n_0 ),
        .O(\r_c[14]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCC55)) 
    \r_c[14]_i_1__2 
       (.I0(\r_c[14]_i_2__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [15]),
        .I2(\r_c[14]_i_3__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I4(\r_c[14]_i_4__1_n_0 ),
        .O(\r_c[14]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCC55)) 
    \r_c[14]_i_1__3 
       (.I0(\r_c[14]_i_2__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [15]),
        .I2(\r_c[14]_i_3__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I4(\r_c[14]_i_4__2_n_0 ),
        .O(\r_c[14]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCC55)) 
    \r_c[14]_i_1__4 
       (.I0(\r_c[14]_i_2__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [15]),
        .I2(\r_c[14]_i_3__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I4(\r_c[14]_i_4__3_n_0 ),
        .O(\r_c[14]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCC55)) 
    \r_c[14]_i_1__5 
       (.I0(\r_c[14]_i_2__4_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [15]),
        .I2(\r_c[14]_i_3__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I4(\r_c[14]_i_4__4_n_0 ),
        .O(\r_c[14]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCC55)) 
    \r_c[14]_i_1__6 
       (.I0(\r_c[14]_i_2__5_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [15]),
        .I2(\r_c[14]_i_3__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I4(\r_c[14]_i_4__5_n_0 ),
        .O(\r_c[14]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCC55)) 
    \r_c[14]_i_1__7 
       (.I0(\r_c[14]_i_2__7_n_0 ),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [15]),
        .I2(\r_c[14]_i_3__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\r_c[14]_i_4__7_n_0 ),
        .O(\r_c[14]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCC55)) 
    \r_c[14]_i_1__8 
       (.I0(\r_c[14]_i_2__8_n_0 ),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [15]),
        .I2(\r_c[14]_i_3__8_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\r_c[14]_i_4__8_n_0 ),
        .O(\r_c[14]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[14]_i_2 
       (.I0(\r_c[14]_i_5_n_0 ),
        .I1(\r_c[1]_i_3_n_0 ),
        .I2(\r_c[14]_i_6_n_0 ),
        .O(\r_c[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[14]_i_2__0 
       (.I0(\r_c[14]_i_5__0_n_0 ),
        .I1(\r_c[1]_i_3__0_n_0 ),
        .I2(\r_c[14]_i_6__0_n_0 ),
        .O(\r_c[14]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[14]_i_2__1 
       (.I0(\r_c[14]_i_5__1_n_0 ),
        .I1(\r_c[1]_i_3__1_n_0 ),
        .I2(\r_c[14]_i_6__1_n_0 ),
        .O(\r_c[14]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[14]_i_2__2 
       (.I0(\r_c[14]_i_5__2_n_0 ),
        .I1(\r_c[1]_i_3__2_n_0 ),
        .I2(\r_c[14]_i_6__2_n_0 ),
        .O(\r_c[14]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[14]_i_2__3 
       (.I0(\r_c[14]_i_5__3_n_0 ),
        .I1(\r_c[1]_i_3__3_n_0 ),
        .I2(\r_c[14]_i_6__3_n_0 ),
        .O(\r_c[14]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[14]_i_2__4 
       (.I0(\r_c[14]_i_5__4_n_0 ),
        .I1(\r_c[1]_i_3__4_n_0 ),
        .I2(\r_c[14]_i_6__4_n_0 ),
        .O(\r_c[14]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[14]_i_2__5 
       (.I0(\r_c[14]_i_5__5_n_0 ),
        .I1(\r_c[1]_i_3__5_n_0 ),
        .I2(\r_c[14]_i_6__5_n_0 ),
        .O(\r_c[14]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0E08080E0E0E0E0E)) 
    \r_c[14]_i_2__6 
       (.I0(\r_c[14]_i_5__6_n_0 ),
        .I1(\u_geo/u_geo_persdiv/r_ce_tmp [4]),
        .I2(\r_c[20]_i_4_n_0 ),
        .I3(\r_c[17]_i_2_n_0 ),
        .I4(\u_geo/u_geo_persdiv/r_ce_tmp [0]),
        .I5(\r_c[14]_i_6__8_n_0 ),
        .O(\r_c[14]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[14]_i_2__7 
       (.I0(\r_c[14]_i_5__7_n_0 ),
        .I1(\r_c[1]_i_3__6_n_0 ),
        .I2(\r_c[14]_i_6__6_n_0 ),
        .O(\r_c[14]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[14]_i_2__8 
       (.I0(\r_c[14]_i_5__8_n_0 ),
        .I1(\r_c[1]_i_3__7_n_0 ),
        .I2(\r_c[14]_i_6__7_n_0 ),
        .O(\r_c[14]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \r_c[14]_i_3 
       (.I0(\r_c[14]_i_7_n_0 ),
        .I1(\r_c[14]_i_8_n_0 ),
        .I2(\r_c[1]_i_3_n_0 ),
        .O(\r_c[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \r_c[14]_i_3__0 
       (.I0(\r_c[14]_i_7__0_n_0 ),
        .I1(\r_c[14]_i_8__0_n_0 ),
        .I2(\r_c[1]_i_3__0_n_0 ),
        .O(\r_c[14]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \r_c[14]_i_3__1 
       (.I0(\r_c[14]_i_7__1_n_0 ),
        .I1(\r_c[14]_i_8__1_n_0 ),
        .I2(\r_c[1]_i_3__1_n_0 ),
        .O(\r_c[14]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \r_c[14]_i_3__2 
       (.I0(\r_c[14]_i_7__2_n_0 ),
        .I1(\r_c[14]_i_8__2_n_0 ),
        .I2(\r_c[1]_i_3__2_n_0 ),
        .O(\r_c[14]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \r_c[14]_i_3__3 
       (.I0(\r_c[14]_i_7__3_n_0 ),
        .I1(\r_c[14]_i_8__3_n_0 ),
        .I2(\r_c[1]_i_3__3_n_0 ),
        .O(\r_c[14]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \r_c[14]_i_3__4 
       (.I0(\r_c[14]_i_7__4_n_0 ),
        .I1(\r_c[14]_i_8__4_n_0 ),
        .I2(\r_c[1]_i_3__4_n_0 ),
        .O(\r_c[14]_i_3__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \r_c[14]_i_3__5 
       (.I0(\r_c[14]_i_7__5_n_0 ),
        .I1(\r_c[14]_i_8__5_n_0 ),
        .I2(\r_c[1]_i_3__5_n_0 ),
        .O(\r_c[14]_i_3__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_c[14]_i_3__6 
       (.I0(\r_c[14]_i_7__6_n_0 ),
        .I1(\r_c[17]_i_3_n_0 ),
        .I2(\r_c[14]_i_8__6_n_0 ),
        .O(\r_c[14]_i_3__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \r_c[14]_i_3__7 
       (.I0(\r_c[14]_i_7__7_n_0 ),
        .I1(\r_c[14]_i_8__7_n_0 ),
        .I2(\r_c[1]_i_3__6_n_0 ),
        .O(\r_c[14]_i_3__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \r_c[14]_i_3__8 
       (.I0(\r_c[14]_i_7__8_n_0 ),
        .I1(\r_c[14]_i_8__8_n_0 ),
        .I2(\r_c[1]_i_3__7_n_0 ),
        .O(\r_c[14]_i_3__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEFEFEEEEEFEFF)) 
    \r_c[14]_i_4 
       (.I0(\r_c[14]_i_9_n_0 ),
        .I1(\r_c[14]_i_10_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [7]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [6]),
        .I4(\r_c[14]_i_11_n_0 ),
        .I5(\r_c[14]_i_12_n_0 ),
        .O(\r_c[14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEFEFEEEEEFEFF)) 
    \r_c[14]_i_4__0 
       (.I0(\r_c[14]_i_9__0_n_0 ),
        .I1(\r_c[14]_i_10__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [7]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [6]),
        .I4(\r_c[14]_i_11__0_n_0 ),
        .I5(\r_c[14]_i_12__0_n_0 ),
        .O(\r_c[14]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEFEFEEEEEFEFF)) 
    \r_c[14]_i_4__1 
       (.I0(\r_c[14]_i_9__1_n_0 ),
        .I1(\r_c[14]_i_10__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [7]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [6]),
        .I4(\r_c[14]_i_11__1_n_0 ),
        .I5(\r_c[14]_i_12__1_n_0 ),
        .O(\r_c[14]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEFEFEEEEEFEFF)) 
    \r_c[14]_i_4__2 
       (.I0(\r_c[14]_i_9__2_n_0 ),
        .I1(\r_c[14]_i_10__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [7]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [6]),
        .I4(\r_c[14]_i_11__2_n_0 ),
        .I5(\r_c[14]_i_12__2_n_0 ),
        .O(\r_c[14]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEFEFEEEEEFEFF)) 
    \r_c[14]_i_4__3 
       (.I0(\r_c[14]_i_9__3_n_0 ),
        .I1(\r_c[14]_i_10__3_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [7]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [6]),
        .I4(\r_c[14]_i_11__3_n_0 ),
        .I5(\r_c[14]_i_12__3_n_0 ),
        .O(\r_c[14]_i_4__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEFEFEEEEEFEFF)) 
    \r_c[14]_i_4__4 
       (.I0(\r_c[14]_i_9__4_n_0 ),
        .I1(\r_c[14]_i_10__4_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [7]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [6]),
        .I4(\r_c[14]_i_11__4_n_0 ),
        .I5(\r_c[14]_i_12__4_n_0 ),
        .O(\r_c[14]_i_4__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEFEFEEEEEFEFF)) 
    \r_c[14]_i_4__5 
       (.I0(\r_c[14]_i_9__5_n_0 ),
        .I1(\r_c[14]_i_10__5_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [7]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [6]),
        .I4(\r_c[14]_i_11__5_n_0 ),
        .I5(\r_c[14]_i_12__5_n_0 ),
        .O(\r_c[14]_i_4__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8A)) 
    \r_c[14]_i_4__6 
       (.I0(\r_c[20]_i_7_n_0 ),
        .I1(\r_c[20]_i_6_n_0 ),
        .I2(\r_c[17]_i_3_n_0 ),
        .O(\r_c[14]_i_4__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEFEFEEEEEFEFF)) 
    \r_c[14]_i_4__7 
       (.I0(\r_c[14]_i_9__6_n_0 ),
        .I1(\r_c[14]_i_10__6_n_0 ),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [7]),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [6]),
        .I4(\r_c[14]_i_11__6_n_0 ),
        .I5(\r_c[14]_i_12__6_n_0 ),
        .O(\r_c[14]_i_4__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEFEFEEEEEFEFF)) 
    \r_c[14]_i_4__8 
       (.I0(\r_c[14]_i_9__7_n_0 ),
        .I1(\r_c[14]_i_10__7_n_0 ),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [7]),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [6]),
        .I4(\r_c[14]_i_11__7_n_0 ),
        .I5(\r_c[14]_i_12__7_n_0 ),
        .O(\r_c[14]_i_4__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[14]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [7]),
        .I1(_inferred__1_carry_i_7_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [11]),
        .I3(_inferred__1_carry_i_6_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [3]),
        .O(\r_c[14]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[14]_i_5__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [7]),
        .I1(_inferred__1_carry_i_7__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [11]),
        .I3(_inferred__1_carry_i_6__0_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [3]),
        .O(\r_c[14]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[14]_i_5__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [7]),
        .I1(_inferred__1_carry_i_7__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [11]),
        .I3(_inferred__1_carry_i_6__1_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [3]),
        .O(\r_c[14]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[14]_i_5__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [7]),
        .I1(_inferred__1_carry_i_7__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [11]),
        .I3(_inferred__1_carry_i_6__2_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [3]),
        .O(\r_c[14]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[14]_i_5__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [7]),
        .I1(_inferred__1_carry_i_7__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [11]),
        .I3(_inferred__1_carry_i_6__3_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [3]),
        .O(\r_c[14]_i_5__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[14]_i_5__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [7]),
        .I1(_inferred__1_carry_i_7__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [11]),
        .I3(_inferred__1_carry_i_6__4_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [3]),
        .O(\r_c[14]_i_5__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    \r_c[14]_i_5__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [7]),
        .I1(_inferred__1_carry_i_7__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [11]),
        .I3(_inferred__1_carry_i_6__5_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [3]),
        .O(\r_c[14]_i_5__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    \r_c[14]_i_5__6 
       (.I0(\r_c[20]_i_3__6_n_0 ),
        .I1(\r_c[20]_i_2__6_n_0 ),
        .I2(\u_geo/u_geo_persdiv/r_ce_tmp [3]),
        .O(\r_c[14]_i_5__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44CC77CF)) 
    \r_c[14]_i_5__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [7]),
        .I1(_inferred__1_carry_i_7__7_n_0),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [3]),
        .I3(_inferred__1_carry_i_6__7_n_0),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [11]),
        .O(\r_c[14]_i_5__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44CC77CF)) 
    \r_c[14]_i_5__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [7]),
        .I1(_inferred__1_carry_i_7__9_n_0),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [3]),
        .I3(_inferred__1_carry_i_6__9_n_0),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [11]),
        .O(\r_c[14]_i_5__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_6 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [1]),
        .I2(_inferred__1_carry_i_7_n_0),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [13]),
        .I4(_inferred__1_carry_i_6_n_0),
        .I5(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [5]),
        .O(\r_c[14]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_6__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [1]),
        .I2(_inferred__1_carry_i_7__0_n_0),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [13]),
        .I4(_inferred__1_carry_i_6__0_n_0),
        .I5(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [5]),
        .O(\r_c[14]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_6__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [1]),
        .I2(_inferred__1_carry_i_7__1_n_0),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [13]),
        .I4(_inferred__1_carry_i_6__1_n_0),
        .I5(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [5]),
        .O(\r_c[14]_i_6__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_6__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [1]),
        .I2(_inferred__1_carry_i_7__2_n_0),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [13]),
        .I4(_inferred__1_carry_i_6__2_n_0),
        .I5(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [5]),
        .O(\r_c[14]_i_6__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_6__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [9]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [1]),
        .I2(_inferred__1_carry_i_7__3_n_0),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [13]),
        .I4(_inferred__1_carry_i_6__3_n_0),
        .I5(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [5]),
        .O(\r_c[14]_i_6__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_6__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [9]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [1]),
        .I2(_inferred__1_carry_i_7__4_n_0),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [13]),
        .I4(_inferred__1_carry_i_6__4_n_0),
        .I5(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [5]),
        .O(\r_c[14]_i_6__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_6__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [9]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [1]),
        .I2(_inferred__1_carry_i_7__5_n_0),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [13]),
        .I4(_inferred__1_carry_i_6__5_n_0),
        .I5(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [5]),
        .O(\r_c[14]_i_6__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_6__6 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [1]),
        .I2(_inferred__1_carry_i_7__7_n_0),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [13]),
        .I4(_inferred__1_carry_i_6__7_n_0),
        .I5(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [5]),
        .O(\r_c[14]_i_6__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_6__7 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [1]),
        .I2(_inferred__1_carry_i_7__9_n_0),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [13]),
        .I4(_inferred__1_carry_i_6__9_n_0),
        .I5(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [5]),
        .O(\r_c[14]_i_6__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r_c[14]_i_6__8 
       (.I0(\u_geo/u_geo_persdiv/r_ce_tmp [1]),
        .I1(\r_c[17]_i_3_n_0 ),
        .O(\r_c[14]_i_6__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_7 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [10]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [2]),
        .I2(_inferred__1_carry_i_7_n_0),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_6_n_0),
        .I5(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [6]),
        .O(\r_c[14]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_7__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [10]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [2]),
        .I2(_inferred__1_carry_i_7__0_n_0),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_6__0_n_0),
        .I5(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [6]),
        .O(\r_c[14]_i_7__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_7__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [10]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [2]),
        .I2(_inferred__1_carry_i_7__1_n_0),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_6__1_n_0),
        .I5(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [6]),
        .O(\r_c[14]_i_7__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_7__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [10]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [2]),
        .I2(_inferred__1_carry_i_7__2_n_0),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_6__2_n_0),
        .I5(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [6]),
        .O(\r_c[14]_i_7__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_7__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [10]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [2]),
        .I2(_inferred__1_carry_i_7__3_n_0),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [14]),
        .I4(_inferred__1_carry_i_6__3_n_0),
        .I5(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [6]),
        .O(\r_c[14]_i_7__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_7__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [10]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [2]),
        .I2(_inferred__1_carry_i_7__4_n_0),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [14]),
        .I4(_inferred__1_carry_i_6__4_n_0),
        .I5(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [6]),
        .O(\r_c[14]_i_7__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_7__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [10]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [2]),
        .I2(_inferred__1_carry_i_7__5_n_0),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [14]),
        .I4(_inferred__1_carry_i_6__5_n_0),
        .I5(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [6]),
        .O(\r_c[14]_i_7__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC4C4C7F7)) 
    \r_c[14]_i_7__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [7]),
        .I1(\r_c[18]_i_3_n_0 ),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [3]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [11]),
        .O(\r_c[14]_i_7__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_7__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [10]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [2]),
        .I2(_inferred__1_carry_i_7__7_n_0),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_6__7_n_0),
        .I5(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [6]),
        .O(\r_c[14]_i_7__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_7__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [10]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [2]),
        .I2(_inferred__1_carry_i_7__9_n_0),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [14]),
        .I4(_inferred__1_carry_i_6__9_n_0),
        .I5(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [6]),
        .O(\r_c[14]_i_7__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_8 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [8]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [0]),
        .I2(_inferred__1_carry_i_7_n_0),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [12]),
        .I4(_inferred__1_carry_i_6_n_0),
        .I5(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [4]),
        .O(\r_c[14]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_8__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [8]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [0]),
        .I2(_inferred__1_carry_i_7__0_n_0),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [12]),
        .I4(_inferred__1_carry_i_6__0_n_0),
        .I5(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [4]),
        .O(\r_c[14]_i_8__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_8__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [8]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [0]),
        .I2(_inferred__1_carry_i_7__1_n_0),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [12]),
        .I4(_inferred__1_carry_i_6__1_n_0),
        .I5(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [4]),
        .O(\r_c[14]_i_8__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_8__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [8]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [0]),
        .I2(_inferred__1_carry_i_7__2_n_0),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [12]),
        .I4(_inferred__1_carry_i_6__2_n_0),
        .I5(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [4]),
        .O(\r_c[14]_i_8__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_8__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [8]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [0]),
        .I2(_inferred__1_carry_i_7__3_n_0),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [12]),
        .I4(_inferred__1_carry_i_6__3_n_0),
        .I5(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [4]),
        .O(\r_c[14]_i_8__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_8__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [8]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [0]),
        .I2(_inferred__1_carry_i_7__4_n_0),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [12]),
        .I4(_inferred__1_carry_i_6__4_n_0),
        .I5(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [4]),
        .O(\r_c[14]_i_8__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_8__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [8]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [0]),
        .I2(_inferred__1_carry_i_7__5_n_0),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [12]),
        .I4(_inferred__1_carry_i_6__5_n_0),
        .I5(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [4]),
        .O(\r_c[14]_i_8__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000051515151515)) 
    \r_c[14]_i_8__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [13]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [5]),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [1]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [9]),
        .I5(\r_c[18]_i_3_n_0 ),
        .O(\r_c[14]_i_8__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_8__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [8]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [0]),
        .I2(_inferred__1_carry_i_7__7_n_0),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [12]),
        .I4(_inferred__1_carry_i_6__7_n_0),
        .I5(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [4]),
        .O(\r_c[14]_i_8__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F1010505F101F)) 
    \r_c[14]_i_8__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [8]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [0]),
        .I2(_inferred__1_carry_i_7__9_n_0),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [12]),
        .I4(_inferred__1_carry_i_6__9_n_0),
        .I5(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [4]),
        .O(\r_c[14]_i_8__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \r_c[14]_i_9 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [12]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [14]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [10]),
        .O(\r_c[14]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \r_c[14]_i_9__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [12]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [14]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [10]),
        .O(\r_c[14]_i_9__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \r_c[14]_i_9__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [12]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [14]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [10]),
        .O(\r_c[14]_i_9__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \r_c[14]_i_9__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [12]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [14]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [10]),
        .O(\r_c[14]_i_9__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \r_c[14]_i_9__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [9]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [12]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [14]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [10]),
        .O(\r_c[14]_i_9__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \r_c[14]_i_9__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [9]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [12]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [14]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [10]),
        .O(\r_c[14]_i_9__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \r_c[14]_i_9__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [9]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [12]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [14]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [10]),
        .O(\r_c[14]_i_9__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \r_c[14]_i_9__6 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [12]),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [14]),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [10]),
        .O(\r_c[14]_i_9__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \r_c[14]_i_9__7 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [9]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [12]),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [14]),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [10]),
        .O(\r_c[14]_i_9__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF00FF00FF00FE)) 
    \r_c[15]_i_1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [4]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [0]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [2]),
        .I3(\r_c[20]_i_2_n_0 ),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [3]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [1]),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/w_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF00FF00FF00FE)) 
    \r_c[15]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [4]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [0]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [2]),
        .I3(\r_c[20]_i_2__0_n_0 ),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [3]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [1]),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/w_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF00FF00FF00FE)) 
    \r_c[15]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [4]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [0]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [2]),
        .I3(\r_c[20]_i_2__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [3]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [1]),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/w_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF00FF00FF00FE)) 
    \r_c[15]_i_1__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [4]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [0]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [2]),
        .I3(\r_c[20]_i_2__2_n_0 ),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [3]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [1]),
        .O(\u_geo/u_geo_matrix/u_fmul_m3/w_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF00FF00FF00FE)) 
    \r_c[15]_i_1__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [4]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [0]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [2]),
        .I3(\r_c[20]_i_2__3_n_0 ),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [3]),
        .I5(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [1]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF00FF00FF00FE)) 
    \r_c[15]_i_1__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [4]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [0]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [2]),
        .I3(\r_c[20]_i_2__4_n_0 ),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [3]),
        .I5(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [1]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF00FF00FF00FE)) 
    \r_c[15]_i_1__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [4]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [0]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [2]),
        .I3(\r_c[20]_i_2__5_n_0 ),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [3]),
        .I5(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [1]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \r_c[15]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [1]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [4]),
        .I2(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [0]),
        .I3(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF00FF00FF00FE)) 
    \r_c[15]_i_1__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [0]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [2]),
        .I2(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [1]),
        .I3(\r_c[20]_i_2__7_n_0 ),
        .I4(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [4]),
        .I5(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [3]),
        .O(\u_geo/u_geo_persdiv/u_fmul/w_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF00FF00FF00FE)) 
    \r_c[15]_i_1__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [0]),
        .I1(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [2]),
        .I2(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [1]),
        .I3(\r_c[20]_i_2__9_n_0 ),
        .I4(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [4]),
        .I5(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [3]),
        .O(\u_geo/u_geo_viewport/u_fmul/w_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair297" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[16]_i_1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [0]),
        .I1(\r_c[20]_i_2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/norm/w_c_exp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair294" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[16]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [0]),
        .I1(\r_c[20]_i_2__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/norm/w_c_exp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair292" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[16]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [0]),
        .I1(\r_c[20]_i_2__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/norm/w_c_exp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair289" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[16]_i_1__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [0]),
        .I1(\r_c[20]_i_2__2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m3/norm/w_c_exp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[16]_i_1__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [0]),
        .I1(\r_c[20]_i_2__3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/norm/w_c_exp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[16]_i_1__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [0]),
        .I1(\r_c[20]_i_2__4_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/norm/w_c_exp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair285" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[16]_i_1__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [0]),
        .I1(\r_c[20]_i_2__5_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/norm/w_c_exp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1001)) 
    \r_c[16]_i_1__6 
       (.I0(\r_c[18]_i_2_n_0 ),
        .I1(\r_c[20]_i_4_n_0 ),
        .I2(\r_c[17]_i_2_n_0 ),
        .I3(\u_geo/u_geo_persdiv/r_ce_tmp [0]),
        .O(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[16]_i_1__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [0]),
        .I1(\r_c[20]_i_2__7_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_fmul/norm/w_c_exp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair287" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[16]_i_1__8 
       (.I0(\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [0]),
        .I1(\r_c[20]_i_2__8_n_0 ),
        .O(\u_geo/u_geo_viewport/u_fadd/norm/w_c_exp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[16]_i_1__9 
       (.I0(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [0]),
        .I1(\r_c[20]_i_2__9_n_0 ),
        .O(\u_geo/u_geo_viewport/u_fmul/norm/w_c_exp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[17]_i_1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [1]),
        .I1(\r_c[20]_i_2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/norm/w_c_exp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r_c[17]_i_10 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [8]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [9]),
        .O(\r_c[17]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r_c[17]_i_11 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [12]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [13]),
        .O(\r_c[17]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[17]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [1]),
        .I1(\r_c[20]_i_2__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/norm/w_c_exp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[17]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [1]),
        .I1(\r_c[20]_i_2__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/norm/w_c_exp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[17]_i_1__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [1]),
        .I1(\r_c[20]_i_2__2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m3/norm/w_c_exp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[17]_i_1__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [1]),
        .I1(\r_c[20]_i_2__3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/norm/w_c_exp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair296" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[17]_i_1__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [1]),
        .I1(\r_c[20]_i_2__4_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/norm/w_c_exp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair285" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[17]_i_1__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [1]),
        .I1(\r_c[20]_i_2__5_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/norm/w_c_exp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000001EE1)) 
    \r_c[17]_i_1__6 
       (.I0(\r_c[17]_i_2_n_0 ),
        .I1(\u_geo/u_geo_persdiv/r_ce_tmp [0]),
        .I2(\r_c[17]_i_3_n_0 ),
        .I3(\u_geo/u_geo_persdiv/r_ce_tmp [1]),
        .I4(\r_c[20]_i_4_n_0 ),
        .I5(\r_c[18]_i_2_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair288" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[17]_i_1__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [1]),
        .I1(\r_c[20]_i_2__7_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_fmul/norm/w_c_exp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair287" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[17]_i_1__8 
       (.I0(\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [1]),
        .I1(\r_c[20]_i_2__8_n_0 ),
        .O(\u_geo/u_geo_viewport/u_fadd/norm/w_c_exp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[17]_i_1__9 
       (.I0(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [1]),
        .I1(\r_c[20]_i_2__9_n_0 ),
        .O(\u_geo/u_geo_viewport/u_fmul/norm/w_c_exp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF0FFF0FFFFFFF1)) 
    \r_c[17]_i_2 
       (.I0(\r_c[17]_i_4_n_0 ),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [6]),
        .I2(\r_c[17]_i_5_n_0 ),
        .I3(\r_c[17]_i_6_n_0 ),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [7]),
        .I5(\r_c[17]_i_7_n_0 ),
        .O(\r_c[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000101011111111)) 
    \r_c[17]_i_3 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [14]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [15]),
        .I2(\r_c[17]_i_8_n_0 ),
        .I3(\r_c[17]_i_9_n_0 ),
        .I4(\r_c[17]_i_10_n_0 ),
        .I5(\r_c[17]_i_11_n_0 ),
        .O(\r_c[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551011)) 
    \r_c[17]_i_4 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [5]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [3]),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [2]),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [1]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [4]),
        .O(\r_c[17]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \r_c[17]_i_5 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [9]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [12]),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [14]),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [10]),
        .O(\r_c[17]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00F4)) 
    \r_c[17]_i_6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [12]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [11]),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [13]),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [14]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [15]),
        .O(\r_c[17]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r_c[17]_i_7 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [8]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [12]),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [14]),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [10]),
        .O(\r_c[17]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r_c[17]_i_8 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [10]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [11]),
        .O(\r_c[17]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1110111011101111)) 
    \r_c[17]_i_9 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [7]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [6]),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [4]),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [5]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [2]),
        .I5(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [3]),
        .O(\r_c[17]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair298" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[18]_i_1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [2]),
        .I1(\r_c[20]_i_2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/norm/w_c_exp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair295" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[18]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [2]),
        .I1(\r_c[20]_i_2__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/norm/w_c_exp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[18]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [2]),
        .I1(\r_c[20]_i_2__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/norm/w_c_exp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[18]_i_1__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [2]),
        .I1(\r_c[20]_i_2__2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m3/norm/w_c_exp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[18]_i_1__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [2]),
        .I1(\r_c[20]_i_2__3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/norm/w_c_exp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[18]_i_1__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [2]),
        .I1(\r_c[20]_i_2__4_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/norm/w_c_exp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair299" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[18]_i_1__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [2]),
        .I1(\r_c[20]_i_2__5_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/norm/w_c_exp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h01101001)) 
    \r_c[18]_i_1__6 
       (.I0(\r_c[18]_i_2_n_0 ),
        .I1(\r_c[20]_i_4_n_0 ),
        .I2(\u_geo/u_geo_persdiv/r_ce_tmp [2]),
        .I3(\r_c[18]_i_3_n_0 ),
        .I4(\r_c[18]_i_4_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair288" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[18]_i_1__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [2]),
        .I1(\r_c[20]_i_2__7_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_fmul/norm/w_c_exp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair286" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[18]_i_1__8 
       (.I0(\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [2]),
        .I1(\r_c[20]_i_2__8_n_0 ),
        .O(\u_geo/u_geo_viewport/u_fadd/norm/w_c_exp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[18]_i_1__9 
       (.I0(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [2]),
        .I1(\r_c[20]_i_2__9_n_0 ),
        .O(\u_geo/u_geo_viewport/u_fmul/norm/w_c_exp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1051)) 
    \r_c[18]_i_2 
       (.I0(\u_geo/u_geo_persdiv/r_ce_tmp [4]),
        .I1(\u_geo/u_geo_persdiv/r_ce_tmp [3]),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\r_c[20]_i_3__6_n_0 ),
        .O(\r_c[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000155555555)) 
    \r_c[18]_i_3 
       (.I0(\r_c[20]_i_5_n_0 ),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [7]),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [6]),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [5]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [4]),
        .I5(\r_c[18]_i_5_n_0 ),
        .O(\r_c[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBBB2)) 
    \r_c[18]_i_4 
       (.I0(\u_geo/u_geo_persdiv/r_ce_tmp [1]),
        .I1(\r_c[17]_i_3_n_0 ),
        .I2(\u_geo/u_geo_persdiv/r_ce_tmp [0]),
        .I3(\r_c[17]_i_2_n_0 ),
        .O(\r_c[18]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \r_c[18]_i_5 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [9]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [8]),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [11]),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [10]),
        .O(\r_c[18]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair297" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[19]_i_1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [3]),
        .I1(\r_c[20]_i_2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/norm/w_c_exp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair294" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[19]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [3]),
        .I1(\r_c[20]_i_2__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/norm/w_c_exp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair292" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[19]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [3]),
        .I1(\r_c[20]_i_2__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/norm/w_c_exp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair289" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[19]_i_1__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [3]),
        .I1(\r_c[20]_i_2__2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m3/norm/w_c_exp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[19]_i_1__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [3]),
        .I1(\r_c[20]_i_2__3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/norm/w_c_exp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[19]_i_1__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [3]),
        .I1(\r_c[20]_i_2__4_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/norm/w_c_exp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[19]_i_1__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [3]),
        .I1(\r_c[20]_i_2__5_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/norm/w_c_exp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h14410400)) 
    \r_c[19]_i_1__6 
       (.I0(\r_c[20]_i_4_n_0 ),
        .I1(\r_c[20]_i_3__6_n_0 ),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/r_ce_tmp [3]),
        .I4(\u_geo/u_geo_persdiv/r_ce_tmp [4]),
        .O(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[19]_i_1__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [3]),
        .I1(\r_c[20]_i_2__7_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_fmul/norm/w_c_exp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[19]_i_1__8 
       (.I0(\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [3]),
        .I1(\r_c[20]_i_2__8_n_0 ),
        .O(\u_geo/u_geo_viewport/u_fadd/norm/w_c_exp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[19]_i_1__9 
       (.I0(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [3]),
        .I1(\r_c[20]_i_2__9_n_0 ),
        .O(\u_geo/u_geo_viewport/u_fmul/norm/w_c_exp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888B8888888BBB)) 
    \r_c[1]_i_1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [2]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I2(\r_c[1]_i_2_n_0 ),
        .I3(\r_c[14]_i_4_n_0 ),
        .I4(\r_c[1]_i_3_n_0 ),
        .I5(\r_c[1]_i_4_n_0 ),
        .O(\r_c[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888B8888888BBB)) 
    \r_c[1]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [2]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I2(\r_c[1]_i_2__0_n_0 ),
        .I3(\r_c[14]_i_4__0_n_0 ),
        .I4(\r_c[1]_i_3__0_n_0 ),
        .I5(\r_c[1]_i_4__0_n_0 ),
        .O(\r_c[1]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888B8888888BBB)) 
    \r_c[1]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [2]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I2(\r_c[1]_i_2__1_n_0 ),
        .I3(\r_c[14]_i_4__1_n_0 ),
        .I4(\r_c[1]_i_3__1_n_0 ),
        .I5(\r_c[1]_i_4__1_n_0 ),
        .O(\r_c[1]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888B8888888BBB)) 
    \r_c[1]_i_1__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [2]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I2(\r_c[1]_i_2__2_n_0 ),
        .I3(\r_c[14]_i_4__2_n_0 ),
        .I4(\r_c[1]_i_3__2_n_0 ),
        .I5(\r_c[1]_i_4__2_n_0 ),
        .O(\r_c[1]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888B8888888BBB)) 
    \r_c[1]_i_1__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [2]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I2(\r_c[1]_i_2__3_n_0 ),
        .I3(\r_c[14]_i_4__3_n_0 ),
        .I4(\r_c[1]_i_3__3_n_0 ),
        .I5(\r_c[1]_i_4__3_n_0 ),
        .O(\r_c[1]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888B8888888BBB)) 
    \r_c[1]_i_1__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [2]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I2(\r_c[1]_i_2__4_n_0 ),
        .I3(\r_c[14]_i_4__4_n_0 ),
        .I4(\r_c[1]_i_3__4_n_0 ),
        .I5(\r_c[1]_i_4__4_n_0 ),
        .O(\r_c[1]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888B8888888BBB)) 
    \r_c[1]_i_1__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [2]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I2(\r_c[1]_i_2__5_n_0 ),
        .I3(\r_c[14]_i_4__5_n_0 ),
        .I4(\r_c[1]_i_3__5_n_0 ),
        .I5(\r_c[1]_i_4__5_n_0 ),
        .O(\r_c[1]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFFFFE)) 
    \r_c[1]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [0]),
        .I3(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [4]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [1]),
        .I5(\r_c[1]_i_2__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCC000FCCCC0505)) 
    \r_c[1]_i_1__7 
       (.I0(\r_c[1]_i_2__7_n_0 ),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [2]),
        .I2(\r_c[1]_i_3__6_n_0 ),
        .I3(\r_c[1]_i_4__6_n_0 ),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I5(\r_c[14]_i_4__7_n_0 ),
        .O(\r_c[1]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCC000FCCCC0505)) 
    \r_c[1]_i_1__8 
       (.I0(\r_c[1]_i_2__8_n_0 ),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [2]),
        .I2(\r_c[1]_i_3__7_n_0 ),
        .I3(\r_c[1]_i_4__7_n_0 ),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I5(\r_c[14]_i_4__8_n_0 ),
        .O(\r_c[1]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_2 
       (.I0(_inferred__1_carry_i_7_n_0),
        .I1(_inferred__1_carry_i_6_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [1]),
        .O(\r_c[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_2__0 
       (.I0(_inferred__1_carry_i_7__0_n_0),
        .I1(_inferred__1_carry_i_6__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [1]),
        .O(\r_c[1]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_2__1 
       (.I0(_inferred__1_carry_i_7__1_n_0),
        .I1(_inferred__1_carry_i_6__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [1]),
        .O(\r_c[1]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_2__2 
       (.I0(_inferred__1_carry_i_7__2_n_0),
        .I1(_inferred__1_carry_i_6__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [1]),
        .O(\r_c[1]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_2__3 
       (.I0(_inferred__1_carry_i_7__3_n_0),
        .I1(_inferred__1_carry_i_6__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [1]),
        .O(\r_c[1]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_2__4 
       (.I0(_inferred__1_carry_i_7__4_n_0),
        .I1(_inferred__1_carry_i_6__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [1]),
        .O(\r_c[1]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_2__5 
       (.I0(_inferred__1_carry_i_7__5_n_0),
        .I1(_inferred__1_carry_i_6__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [1]),
        .O(\r_c[1]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF4FFF7)) 
    \r_c[1]_i_2__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [1]),
        .I1(\r_c[17]_i_2_n_0 ),
        .I2(\r_c[17]_i_3_n_0 ),
        .I3(\r_c[20]_i_2__6_n_0 ),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [0]),
        .I5(\r_c[18]_i_3_n_0 ),
        .O(\r_c[1]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_2__7 
       (.I0(_inferred__1_carry_i_7__7_n_0),
        .I1(_inferred__1_carry_i_6__7_n_0),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [0]),
        .O(\r_c[1]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_2__8 
       (.I0(_inferred__1_carry_i_7__9_n_0),
        .I1(_inferred__1_carry_i_6__9_n_0),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [0]),
        .O(\r_c[1]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [14]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [15]),
        .I2(\r_c[1]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [12]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [13]),
        .O(\r_c[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_3__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [14]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [15]),
        .I2(\r_c[1]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [12]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [13]),
        .O(\r_c[1]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_3__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [14]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [15]),
        .I2(\r_c[1]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [12]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [13]),
        .O(\r_c[1]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_3__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [14]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [15]),
        .I2(\r_c[1]_i_5__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [12]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [13]),
        .O(\r_c[1]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_3__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [14]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [15]),
        .I2(\r_c[1]_i_5__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [12]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [13]),
        .O(\r_c[1]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_3__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [14]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [15]),
        .I2(\r_c[1]_i_5__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [12]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [13]),
        .O(\r_c[1]_i_3__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_3__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [14]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [15]),
        .I2(\r_c[1]_i_5__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [12]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [13]),
        .O(\r_c[1]_i_3__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_3__6 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [14]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [15]),
        .I2(\r_c[1]_i_5__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [12]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [13]),
        .O(\r_c[1]_i_3__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_3__7 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [14]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [15]),
        .I2(\r_c[1]_i_5__7_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [12]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [13]),
        .O(\r_c[1]_i_3__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_4 
       (.I0(_inferred__1_carry_i_7_n_0),
        .I1(_inferred__1_carry_i_6_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [0]),
        .O(\r_c[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_4__0 
       (.I0(_inferred__1_carry_i_7__0_n_0),
        .I1(_inferred__1_carry_i_6__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [0]),
        .O(\r_c[1]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_4__1 
       (.I0(_inferred__1_carry_i_7__1_n_0),
        .I1(_inferred__1_carry_i_6__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [0]),
        .O(\r_c[1]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_4__2 
       (.I0(_inferred__1_carry_i_7__2_n_0),
        .I1(_inferred__1_carry_i_6__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [0]),
        .O(\r_c[1]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_4__3 
       (.I0(_inferred__1_carry_i_7__3_n_0),
        .I1(_inferred__1_carry_i_6__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [0]),
        .O(\r_c[1]_i_4__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_4__4 
       (.I0(_inferred__1_carry_i_7__4_n_0),
        .I1(_inferred__1_carry_i_6__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [0]),
        .O(\r_c[1]_i_4__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_4__5 
       (.I0(_inferred__1_carry_i_7__5_n_0),
        .I1(_inferred__1_carry_i_6__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [0]),
        .O(\r_c[1]_i_4__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_4__6 
       (.I0(_inferred__1_carry_i_7__7_n_0),
        .I1(_inferred__1_carry_i_6__7_n_0),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [1]),
        .O(\r_c[1]_i_4__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r_c[1]_i_4__7 
       (.I0(_inferred__1_carry_i_7__9_n_0),
        .I1(_inferred__1_carry_i_6__9_n_0),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [1]),
        .O(\r_c[1]_i_4__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [11]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [10]),
        .I2(\r_c[1]_i_6_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [8]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [9]),
        .O(\r_c[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_5__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [11]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [10]),
        .I2(\r_c[1]_i_6__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [8]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [9]),
        .O(\r_c[1]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_5__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [11]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [10]),
        .I2(\r_c[1]_i_6__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [8]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [9]),
        .O(\r_c[1]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_5__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [11]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [10]),
        .I2(\r_c[1]_i_6__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [8]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [9]),
        .O(\r_c[1]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_5__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [11]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [10]),
        .I2(\r_c[1]_i_6__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [8]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [9]),
        .O(\r_c[1]_i_5__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_5__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [11]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [10]),
        .I2(\r_c[1]_i_6__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [8]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [9]),
        .O(\r_c[1]_i_5__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_5__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [11]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [10]),
        .I2(\r_c[1]_i_6__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [8]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [9]),
        .O(\r_c[1]_i_5__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_5__6 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [11]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [10]),
        .I2(\r_c[1]_i_6__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [8]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [9]),
        .O(\r_c[1]_i_5__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11111110)) 
    \r_c[1]_i_5__7 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [11]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [10]),
        .I2(\r_c[1]_i_6__7_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [8]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [9]),
        .O(\r_c[1]_i_5__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111111110001)) 
    \r_c[1]_i_6 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [7]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [6]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [2]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [3]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [4]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [5]),
        .O(\r_c[1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111111110001)) 
    \r_c[1]_i_6__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [7]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [6]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [2]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [3]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [4]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [5]),
        .O(\r_c[1]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111111110001)) 
    \r_c[1]_i_6__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [7]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [6]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [2]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [3]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [4]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [5]),
        .O(\r_c[1]_i_6__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111111110001)) 
    \r_c[1]_i_6__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [7]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [6]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [2]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [3]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [4]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [5]),
        .O(\r_c[1]_i_6__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111111110001)) 
    \r_c[1]_i_6__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [7]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [6]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [2]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [3]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [4]),
        .I5(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [5]),
        .O(\r_c[1]_i_6__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111111110001)) 
    \r_c[1]_i_6__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [7]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [6]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [2]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [3]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [4]),
        .I5(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [5]),
        .O(\r_c[1]_i_6__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111111110001)) 
    \r_c[1]_i_6__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [7]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [6]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [2]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [3]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [4]),
        .I5(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [5]),
        .O(\r_c[1]_i_6__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111111110001)) 
    \r_c[1]_i_6__6 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [7]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [6]),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [2]),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [3]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [4]),
        .I5(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [5]),
        .O(\r_c[1]_i_6__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111111110001)) 
    \r_c[1]_i_6__7 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [7]),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [6]),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [2]),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [3]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [4]),
        .I5(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [5]),
        .O(\r_c[1]_i_6__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair298" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[20]_i_1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [4]),
        .I1(\r_c[20]_i_2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/norm/w_c_exp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair295" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[20]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [4]),
        .I1(\r_c[20]_i_2__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/norm/w_c_exp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[20]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [4]),
        .I1(\r_c[20]_i_2__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/norm/w_c_exp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[20]_i_1__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [4]),
        .I1(\r_c[20]_i_2__2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m3/norm/w_c_exp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[20]_i_1__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [4]),
        .I1(\r_c[20]_i_2__3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/norm/w_c_exp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair296" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[20]_i_1__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [4]),
        .I1(\r_c[20]_i_2__4_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/norm/w_c_exp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair299" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[20]_i_1__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [4]),
        .I1(\r_c[20]_i_2__5_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/norm/w_c_exp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000B200)) 
    \r_c[20]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/r_ce_tmp [3]),
        .I1(\r_c[20]_i_2__6_n_0 ),
        .I2(\r_c[20]_i_3__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/r_ce_tmp [4]),
        .I4(\r_c[20]_i_4_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[20]_i_1__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [4]),
        .I1(\r_c[20]_i_2__7_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_fmul/norm/w_c_exp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair286" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[20]_i_1__8 
       (.I0(\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [4]),
        .I1(\r_c[20]_i_2__8_n_0 ),
        .O(\u_geo/u_geo_viewport/u_fadd/norm/w_c_exp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[20]_i_1__9 
       (.I0(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [4]),
        .I1(\r_c[20]_i_2__9_n_0 ),
        .O(\u_geo/u_geo_viewport/u_fmul/norm/w_c_exp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \r_c[20]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [5]),
        .I1(\r_c[20]_i_3_n_0 ),
        .I2(_inferred__1_carry_i_6_n_0),
        .O(\r_c[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \r_c[20]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [5]),
        .I1(\r_c[20]_i_3__0_n_0 ),
        .I2(_inferred__1_carry_i_6__0_n_0),
        .O(\r_c[20]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \r_c[20]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [5]),
        .I1(\r_c[20]_i_3__1_n_0 ),
        .I2(_inferred__1_carry_i_6__1_n_0),
        .O(\r_c[20]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \r_c[20]_i_2__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [5]),
        .I1(\r_c[20]_i_3__2_n_0 ),
        .I2(_inferred__1_carry_i_6__2_n_0),
        .O(\r_c[20]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \r_c[20]_i_2__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [5]),
        .I1(\r_c[20]_i_3__3_n_0 ),
        .I2(_inferred__1_carry_i_6__3_n_0),
        .O(\r_c[20]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \r_c[20]_i_2__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [5]),
        .I1(\r_c[20]_i_3__4_n_0 ),
        .I2(_inferred__1_carry_i_6__4_n_0),
        .O(\r_c[20]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \r_c[20]_i_2__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [5]),
        .I1(\r_c[20]_i_3__5_n_0 ),
        .I2(_inferred__1_carry_i_6__5_n_0),
        .O(\r_c[20]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \r_c[20]_i_2__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [10]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [11]),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [8]),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [9]),
        .I4(\r_c[20]_i_5_n_0 ),
        .O(\r_c[20]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \r_c[20]_i_2__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [5]),
        .I1(\r_c[20]_i_3__7_n_0 ),
        .I2(_inferred__1_carry_i_6__7_n_0),
        .O(\r_c[20]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \r_c[20]_i_2__8 
       (.I0(\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [5]),
        .I1(\r_c[20]_i_3__8_n_0 ),
        .I2(_inferred__1_carry_i_6__8_n_0),
        .O(\r_c[20]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \r_c[20]_i_2__9 
       (.I0(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [5]),
        .I1(\r_c[20]_i_3__9_n_0 ),
        .I2(_inferred__1_carry_i_6__9_n_0),
        .O(\r_c[20]_i_2__9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r_c[20]_i_3 
       (.I0(_inferred__1_carry_i_10_n_0),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [0]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [1]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [2]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [3]),
        .O(\r_c[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r_c[20]_i_3__0 
       (.I0(_inferred__1_carry_i_10__0_n_0),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [0]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [1]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [2]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [3]),
        .O(\r_c[20]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r_c[20]_i_3__1 
       (.I0(_inferred__1_carry_i_10__1_n_0),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [0]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [1]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [2]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [3]),
        .O(\r_c[20]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r_c[20]_i_3__2 
       (.I0(_inferred__1_carry_i_10__2_n_0),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [0]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [1]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [2]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [3]),
        .O(\r_c[20]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r_c[20]_i_3__3 
       (.I0(_inferred__1_carry_i_10__3_n_0),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [0]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [1]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [2]),
        .I5(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [3]),
        .O(\r_c[20]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r_c[20]_i_3__4 
       (.I0(_inferred__1_carry_i_10__4_n_0),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [0]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [1]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [2]),
        .I5(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [3]),
        .O(\r_c[20]_i_3__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r_c[20]_i_3__5 
       (.I0(_inferred__1_carry_i_10__5_n_0),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [0]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [1]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [2]),
        .I5(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [3]),
        .O(\r_c[20]_i_3__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB2FFFF0000BBB2)) 
    \r_c[20]_i_3__6 
       (.I0(\u_geo/u_geo_persdiv/r_ce_tmp [1]),
        .I1(\r_c[17]_i_3_n_0 ),
        .I2(\u_geo/u_geo_persdiv/r_ce_tmp [0]),
        .I3(\r_c[17]_i_2_n_0 ),
        .I4(\r_c[18]_i_3_n_0 ),
        .I5(\u_geo/u_geo_persdiv/r_ce_tmp [2]),
        .O(\r_c[20]_i_3__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r_c[20]_i_3__7 
       (.I0(_inferred__1_carry_i_10__7_n_0),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [0]),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [1]),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [2]),
        .I5(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [3]),
        .O(\r_c[20]_i_3__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r_c[20]_i_3__8 
       (.I0(_inferred__1_carry_i_11__0_n_0),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [0]),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [1]),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [3]),
        .I5(\u_geo/u_geo_viewport/u_fadd/r_mats [2]),
        .O(\r_c[20]_i_3__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r_c[20]_i_3__9 
       (.I0(_inferred__1_carry_i_10__9_n_0),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [0]),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [1]),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [2]),
        .I5(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [3]),
        .O(\r_c[20]_i_3__9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00D0)) 
    \r_c[20]_i_4 
       (.I0(\r_c[17]_i_3_n_0 ),
        .I1(\r_c[20]_i_6_n_0 ),
        .I2(\r_c[20]_i_7_n_0 ),
        .I3(\r_c[17]_i_2_n_0 ),
        .O(\r_c[20]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r_c[20]_i_5 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [14]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [15]),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [13]),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [12]),
        .O(\r_c[20]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000051515151515)) 
    \r_c[20]_i_6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [12]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [4]),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [0]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [8]),
        .I5(\r_c[18]_i_3_n_0 ),
        .O(\r_c[20]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h10301030103F1F3F)) 
    \r_c[20]_i_7 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [10]),
        .I2(\r_c[18]_i_3_n_0 ),
        .I3(\r_c[20]_i_2__6_n_0 ),
        .I4(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [6]),
        .I5(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [14]),
        .O(\r_c[20]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0F0F0F0F0F1)) 
    \r_c[21]_i_1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [1]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [3]),
        .I2(\r_c[20]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [2]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [0]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [4]),
        .O(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0F0F0F0F0F1)) 
    \r_c[21]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [1]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [3]),
        .I2(\r_c[20]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [2]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [0]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [4]),
        .O(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0F0F0F0F0F1)) 
    \r_c[21]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [1]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [3]),
        .I2(\r_c[20]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [2]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [0]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [4]),
        .O(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0F0F0F0F0F1)) 
    \r_c[21]_i_1__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [1]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [3]),
        .I2(\r_c[20]_i_2__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [2]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [0]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [4]),
        .O(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0F0F0F0F0F1)) 
    \r_c[21]_i_1__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [1]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [3]),
        .I2(\r_c[20]_i_2__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [2]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [0]),
        .I5(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [4]),
        .O(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0F0F0F0F0F1)) 
    \r_c[21]_i_1__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [1]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [3]),
        .I2(\r_c[20]_i_2__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [2]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [0]),
        .I5(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [4]),
        .O(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0F0F0F0F0F1)) 
    \r_c[21]_i_1__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [1]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [3]),
        .I2(\r_c[20]_i_2__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [2]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [0]),
        .I5(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [4]),
        .O(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000E00)) 
    \r_c[21]_i_1__6 
       (.I0(\r_c[21]_i_2_n_0 ),
        .I1(\r_c[21]_i_3_n_0 ),
        .I2(\u_geo/u_geo_clip/u_fadd/norm/f_incdec_return [5]),
        .I3(\u_geo/u_geo_clip/u_fadd/r_sign_2z ),
        .I4(\r_c[21]_i_4_n_0 ),
        .O(\u_geo/u_geo_clip/u_fadd/w_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    \r_c[21]_i_1__7 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_a_sign ),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I2(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I3(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [0]),
        .I4(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [4]),
        .I5(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [1]),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r_c[21]_i_1__8 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_sign_2z ),
        .I1(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r_c[21]_i_2 
       (.I0(_inferred__1_carry_i_6__6_n_0),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [1]),
        .I2(\u_geo/u_geo_clip/u_fadd/r_mats [0]),
        .I3(\u_geo/u_geo_clip/u_fadd/r_mats [16]),
        .I4(\u_geo/u_geo_clip/u_fadd/r_mats [2]),
        .I5(\u_geo/u_geo_clip/u_fadd/r_mats [3]),
        .O(\r_c[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    \r_c[21]_i_3 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_mats [15]),
        .I1(\u_geo/u_geo_clip/u_fadd/r_mats [14]),
        .I2(\u_geo/u_geo_clip/u_fadd/r_mats [12]),
        .I3(\u_geo/u_geo_clip/u_fadd/r_mats [13]),
        .I4(_inferred__1_carry_i_7__6_n_0),
        .O(\r_c[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \r_c[21]_i_4 
       (.I0(\u_geo/u_geo_clip/u_fadd/norm/f_incdec_return [2]),
        .I1(\u_geo/u_geo_clip/u_fadd/norm/f_incdec_return [0]),
        .I2(\u_geo/u_geo_clip/u_fadd/norm/f_incdec_return [1]),
        .I3(\u_geo/u_geo_clip/u_fadd/norm/f_incdec_return [4]),
        .I4(\u_geo/u_geo_clip/u_fadd/norm/f_incdec_return [3]),
        .O(\r_c[21]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_c[29]_i_1 
       (.I0(g0_b29_n_0),
        .I1(\u_geo/w_vw_clip [14]),
        .O(\r_c[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[2]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[2]_i_2_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[3]_i_2__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[2]_i_1__0 
       (.I0(\r_c[2]_i_2__0_n_0 ),
        .I1(\r_c[14]_i_4__7_n_0 ),
        .I2(\r_c[3]_i_2__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [3]),
        .O(\r_c[2]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[2]_i_1__1 
       (.I0(\r_c[2]_i_2__1_n_0 ),
        .I1(\r_c[14]_i_4__8_n_0 ),
        .I2(\r_c[3]_i_2__8_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [3]),
        .O(\r_c[2]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCCAA)) 
    \r_c[2]_i_1__2 
       (.I0(\r_c[2]_i_2__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [3]),
        .I2(\r_c[3]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I4(\r_c[14]_i_4_n_0 ),
        .O(\r_c[2]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCCAA)) 
    \r_c[2]_i_1__3 
       (.I0(\r_c[2]_i_2__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [3]),
        .I2(\r_c[3]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I4(\r_c[14]_i_4__0_n_0 ),
        .O(\r_c[2]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCCAA)) 
    \r_c[2]_i_1__4 
       (.I0(\r_c[2]_i_2__4_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [3]),
        .I2(\r_c[3]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I4(\r_c[14]_i_4__1_n_0 ),
        .O(\r_c[2]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCCAA)) 
    \r_c[2]_i_1__5 
       (.I0(\r_c[2]_i_2__5_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [3]),
        .I2(\r_c[3]_i_2__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I4(\r_c[14]_i_4__2_n_0 ),
        .O(\r_c[2]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCCAA)) 
    \r_c[2]_i_1__6 
       (.I0(\r_c[2]_i_2__6_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [3]),
        .I2(\r_c[3]_i_2__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I4(\r_c[14]_i_4__3_n_0 ),
        .O(\r_c[2]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCCAA)) 
    \r_c[2]_i_1__7 
       (.I0(\r_c[2]_i_2__7_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [3]),
        .I2(\r_c[3]_i_2__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I4(\r_c[14]_i_4__4_n_0 ),
        .O(\r_c[2]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC0FCCAA)) 
    \r_c[2]_i_1__8 
       (.I0(\r_c[2]_i_2__8_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [3]),
        .I2(\r_c[3]_i_2__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I4(\r_c[14]_i_4__5_n_0 ),
        .O(\r_c[2]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    \r_c[2]_i_2 
       (.I0(\r_c[17]_i_3_n_0 ),
        .I1(\r_c[20]_i_2__6_n_0 ),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [1]),
        .I3(\r_c[18]_i_3_n_0 ),
        .O(\r_c[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFBF)) 
    \r_c[2]_i_2__0 
       (.I0(\r_c[1]_i_3__6_n_0 ),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [1]),
        .I2(_inferred__1_carry_i_6__7_n_0),
        .I3(_inferred__1_carry_i_7__7_n_0),
        .O(\r_c[2]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFBF)) 
    \r_c[2]_i_2__1 
       (.I0(\r_c[1]_i_3__7_n_0 ),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [1]),
        .I2(_inferred__1_carry_i_6__9_n_0),
        .I3(_inferred__1_carry_i_7__9_n_0),
        .O(\r_c[2]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[2]_i_2__2 
       (.I0(\r_c[1]_i_3_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [1]),
        .I2(_inferred__1_carry_i_6_n_0),
        .I3(_inferred__1_carry_i_7_n_0),
        .O(\r_c[2]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[2]_i_2__3 
       (.I0(\r_c[1]_i_3__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [1]),
        .I2(_inferred__1_carry_i_6__0_n_0),
        .I3(_inferred__1_carry_i_7__0_n_0),
        .O(\r_c[2]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[2]_i_2__4 
       (.I0(\r_c[1]_i_3__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [1]),
        .I2(_inferred__1_carry_i_6__1_n_0),
        .I3(_inferred__1_carry_i_7__1_n_0),
        .O(\r_c[2]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[2]_i_2__5 
       (.I0(\r_c[1]_i_3__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [1]),
        .I2(_inferred__1_carry_i_6__2_n_0),
        .I3(_inferred__1_carry_i_7__2_n_0),
        .O(\r_c[2]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[2]_i_2__6 
       (.I0(\r_c[1]_i_3__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [1]),
        .I2(_inferred__1_carry_i_6__3_n_0),
        .I3(_inferred__1_carry_i_7__3_n_0),
        .O(\r_c[2]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[2]_i_2__7 
       (.I0(\r_c[1]_i_3__4_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [1]),
        .I2(_inferred__1_carry_i_6__4_n_0),
        .I3(_inferred__1_carry_i_7__4_n_0),
        .O(\r_c[2]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \r_c[2]_i_2__8 
       (.I0(\r_c[1]_i_3__5_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [1]),
        .I2(_inferred__1_carry_i_6__5_n_0),
        .I3(_inferred__1_carry_i_7__5_n_0),
        .O(\r_c[2]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT2 #(
    .INIT(4'hD)) 
    \r_c[31]_inv_i_1 
       (.I0(g0_b31_n_0),
        .I1(\u_geo/w_vw_clip [14]),
        .O(\r_c[31]_inv_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[3]_i_1 
       (.I0(\r_c[3]_i_2_n_0 ),
        .I1(\r_c[14]_i_4_n_0 ),
        .I2(\r_c[4]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [4]),
        .O(\r_c[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[3]_i_1__0 
       (.I0(\r_c[3]_i_2__0_n_0 ),
        .I1(\r_c[14]_i_4__0_n_0 ),
        .I2(\r_c[4]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [4]),
        .O(\r_c[3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[3]_i_1__1 
       (.I0(\r_c[3]_i_2__1_n_0 ),
        .I1(\r_c[14]_i_4__1_n_0 ),
        .I2(\r_c[4]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [4]),
        .O(\r_c[3]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[3]_i_1__2 
       (.I0(\r_c[3]_i_2__2_n_0 ),
        .I1(\r_c[14]_i_4__2_n_0 ),
        .I2(\r_c[4]_i_2__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [4]),
        .O(\r_c[3]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[3]_i_1__3 
       (.I0(\r_c[3]_i_2__3_n_0 ),
        .I1(\r_c[14]_i_4__3_n_0 ),
        .I2(\r_c[4]_i_2__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [4]),
        .O(\r_c[3]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[3]_i_1__4 
       (.I0(\r_c[3]_i_2__4_n_0 ),
        .I1(\r_c[14]_i_4__4_n_0 ),
        .I2(\r_c[4]_i_2__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [4]),
        .O(\r_c[3]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[3]_i_1__5 
       (.I0(\r_c[3]_i_2__5_n_0 ),
        .I1(\r_c[14]_i_4__5_n_0 ),
        .I2(\r_c[4]_i_2__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [4]),
        .O(\r_c[3]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[3]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[3]_i_2__6_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[4]_i_2__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[3]_i_1__7 
       (.I0(\r_c[3]_i_2__7_n_0 ),
        .I1(\r_c[14]_i_4__7_n_0 ),
        .I2(\r_c[4]_i_2__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [4]),
        .O(\r_c[3]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[3]_i_1__8 
       (.I0(\r_c[3]_i_2__8_n_0 ),
        .I1(\r_c[14]_i_4__8_n_0 ),
        .I2(\r_c[4]_i_2__8_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [4]),
        .O(\r_c[3]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[3]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [0]),
        .I1(\r_c[1]_i_3_n_0 ),
        .I2(_inferred__1_carry_i_7_n_0),
        .I3(_inferred__1_carry_i_6_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [2]),
        .O(\r_c[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[3]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [0]),
        .I1(\r_c[1]_i_3__0_n_0 ),
        .I2(_inferred__1_carry_i_7__0_n_0),
        .I3(_inferred__1_carry_i_6__0_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [2]),
        .O(\r_c[3]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[3]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [0]),
        .I1(\r_c[1]_i_3__1_n_0 ),
        .I2(_inferred__1_carry_i_7__1_n_0),
        .I3(_inferred__1_carry_i_6__1_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [2]),
        .O(\r_c[3]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[3]_i_2__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [0]),
        .I1(\r_c[1]_i_3__2_n_0 ),
        .I2(_inferred__1_carry_i_7__2_n_0),
        .I3(_inferred__1_carry_i_6__2_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [2]),
        .O(\r_c[3]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[3]_i_2__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [0]),
        .I1(\r_c[1]_i_3__3_n_0 ),
        .I2(_inferred__1_carry_i_7__3_n_0),
        .I3(_inferred__1_carry_i_6__3_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [2]),
        .O(\r_c[3]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[3]_i_2__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [0]),
        .I1(\r_c[1]_i_3__4_n_0 ),
        .I2(_inferred__1_carry_i_7__4_n_0),
        .I3(_inferred__1_carry_i_6__4_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [2]),
        .O(\r_c[3]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[3]_i_2__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [0]),
        .I1(\r_c[1]_i_3__5_n_0 ),
        .I2(_inferred__1_carry_i_7__5_n_0),
        .I3(_inferred__1_carry_i_6__5_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [2]),
        .O(\r_c[3]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \r_c[3]_i_2__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [0]),
        .I1(\r_c[17]_i_3_n_0 ),
        .I2(\r_c[18]_i_3_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [2]),
        .I4(\r_c[20]_i_2__6_n_0 ),
        .O(\r_c[3]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[3]_i_2__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [0]),
        .I1(\r_c[1]_i_3__6_n_0 ),
        .I2(_inferred__1_carry_i_7__7_n_0),
        .I3(_inferred__1_carry_i_6__7_n_0),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [2]),
        .O(\r_c[3]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[3]_i_2__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [0]),
        .I1(\r_c[1]_i_3__7_n_0 ),
        .I2(_inferred__1_carry_i_7__9_n_0),
        .I3(_inferred__1_carry_i_6__9_n_0),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [2]),
        .O(\r_c[3]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[4]_i_1 
       (.I0(\r_c[4]_i_2_n_0 ),
        .I1(\r_c[14]_i_4_n_0 ),
        .I2(\r_c[5]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [5]),
        .O(\r_c[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[4]_i_1__0 
       (.I0(\r_c[4]_i_2__0_n_0 ),
        .I1(\r_c[14]_i_4__0_n_0 ),
        .I2(\r_c[5]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [5]),
        .O(\r_c[4]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[4]_i_1__1 
       (.I0(\r_c[4]_i_2__1_n_0 ),
        .I1(\r_c[14]_i_4__1_n_0 ),
        .I2(\r_c[5]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [5]),
        .O(\r_c[4]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[4]_i_1__2 
       (.I0(\r_c[4]_i_2__2_n_0 ),
        .I1(\r_c[14]_i_4__2_n_0 ),
        .I2(\r_c[5]_i_2__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [5]),
        .O(\r_c[4]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[4]_i_1__3 
       (.I0(\r_c[4]_i_2__3_n_0 ),
        .I1(\r_c[14]_i_4__3_n_0 ),
        .I2(\r_c[5]_i_2__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [5]),
        .O(\r_c[4]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[4]_i_1__4 
       (.I0(\r_c[4]_i_2__4_n_0 ),
        .I1(\r_c[14]_i_4__4_n_0 ),
        .I2(\r_c[5]_i_2__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [5]),
        .O(\r_c[4]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[4]_i_1__5 
       (.I0(\r_c[4]_i_2__5_n_0 ),
        .I1(\r_c[14]_i_4__5_n_0 ),
        .I2(\r_c[5]_i_2__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [5]),
        .O(\r_c[4]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[4]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[4]_i_2__6_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[5]_i_2__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[4]_i_1__7 
       (.I0(\r_c[4]_i_2__7_n_0 ),
        .I1(\r_c[14]_i_4__7_n_0 ),
        .I2(\r_c[5]_i_2__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [5]),
        .O(\r_c[4]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[4]_i_1__8 
       (.I0(\r_c[4]_i_2__8_n_0 ),
        .I1(\r_c[14]_i_4__8_n_0 ),
        .I2(\r_c[5]_i_2__8_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [5]),
        .O(\r_c[4]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[4]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [1]),
        .I1(\r_c[1]_i_3_n_0 ),
        .I2(_inferred__1_carry_i_7_n_0),
        .I3(_inferred__1_carry_i_6_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [3]),
        .O(\r_c[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[4]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [1]),
        .I1(\r_c[1]_i_3__0_n_0 ),
        .I2(_inferred__1_carry_i_7__0_n_0),
        .I3(_inferred__1_carry_i_6__0_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [3]),
        .O(\r_c[4]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[4]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [1]),
        .I1(\r_c[1]_i_3__1_n_0 ),
        .I2(_inferred__1_carry_i_7__1_n_0),
        .I3(_inferred__1_carry_i_6__1_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [3]),
        .O(\r_c[4]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[4]_i_2__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [1]),
        .I1(\r_c[1]_i_3__2_n_0 ),
        .I2(_inferred__1_carry_i_7__2_n_0),
        .I3(_inferred__1_carry_i_6__2_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [3]),
        .O(\r_c[4]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[4]_i_2__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [1]),
        .I1(\r_c[1]_i_3__3_n_0 ),
        .I2(_inferred__1_carry_i_7__3_n_0),
        .I3(_inferred__1_carry_i_6__3_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [3]),
        .O(\r_c[4]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[4]_i_2__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [1]),
        .I1(\r_c[1]_i_3__4_n_0 ),
        .I2(_inferred__1_carry_i_7__4_n_0),
        .I3(_inferred__1_carry_i_6__4_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [3]),
        .O(\r_c[4]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[4]_i_2__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [1]),
        .I1(\r_c[1]_i_3__5_n_0 ),
        .I2(_inferred__1_carry_i_7__5_n_0),
        .I3(_inferred__1_carry_i_6__5_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [3]),
        .O(\r_c[4]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \r_c[4]_i_2__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [1]),
        .I1(\r_c[17]_i_3_n_0 ),
        .I2(\r_c[18]_i_3_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [3]),
        .I4(\r_c[20]_i_2__6_n_0 ),
        .O(\r_c[4]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[4]_i_2__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [1]),
        .I1(\r_c[1]_i_3__6_n_0 ),
        .I2(_inferred__1_carry_i_7__7_n_0),
        .I3(_inferred__1_carry_i_6__7_n_0),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [3]),
        .O(\r_c[4]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    \r_c[4]_i_2__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [1]),
        .I1(\r_c[1]_i_3__7_n_0 ),
        .I2(_inferred__1_carry_i_7__9_n_0),
        .I3(_inferred__1_carry_i_6__9_n_0),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [3]),
        .O(\r_c[4]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[5]_i_1 
       (.I0(\r_c[5]_i_2_n_0 ),
        .I1(\r_c[14]_i_4_n_0 ),
        .I2(\r_c[6]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [6]),
        .O(\r_c[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[5]_i_1__0 
       (.I0(\r_c[5]_i_2__0_n_0 ),
        .I1(\r_c[14]_i_4__0_n_0 ),
        .I2(\r_c[6]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [6]),
        .O(\r_c[5]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[5]_i_1__1 
       (.I0(\r_c[5]_i_2__1_n_0 ),
        .I1(\r_c[14]_i_4__1_n_0 ),
        .I2(\r_c[6]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [6]),
        .O(\r_c[5]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[5]_i_1__2 
       (.I0(\r_c[5]_i_2__2_n_0 ),
        .I1(\r_c[14]_i_4__2_n_0 ),
        .I2(\r_c[6]_i_2__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [6]),
        .O(\r_c[5]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[5]_i_1__3 
       (.I0(\r_c[5]_i_2__3_n_0 ),
        .I1(\r_c[14]_i_4__3_n_0 ),
        .I2(\r_c[6]_i_2__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [6]),
        .O(\r_c[5]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[5]_i_1__4 
       (.I0(\r_c[5]_i_2__4_n_0 ),
        .I1(\r_c[14]_i_4__4_n_0 ),
        .I2(\r_c[6]_i_2__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [6]),
        .O(\r_c[5]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[5]_i_1__5 
       (.I0(\r_c[5]_i_2__5_n_0 ),
        .I1(\r_c[14]_i_4__5_n_0 ),
        .I2(\r_c[6]_i_2__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [6]),
        .O(\r_c[5]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[5]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[5]_i_2__6_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[6]_i_2__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[5]_i_1__7 
       (.I0(\r_c[5]_i_2__7_n_0 ),
        .I1(\r_c[14]_i_4__7_n_0 ),
        .I2(\r_c[6]_i_2__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [6]),
        .O(\r_c[5]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[5]_i_1__8 
       (.I0(\r_c[5]_i_2__8_n_0 ),
        .I1(\r_c[14]_i_4__8_n_0 ),
        .I2(\r_c[6]_i_2__8_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [6]),
        .O(\r_c[5]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[5]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [2]),
        .I1(\r_c[1]_i_3_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [0]),
        .I3(_inferred__1_carry_i_7_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [4]),
        .I5(_inferred__1_carry_i_6_n_0),
        .O(\r_c[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[5]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [2]),
        .I1(\r_c[1]_i_3__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [0]),
        .I3(_inferred__1_carry_i_7__0_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [4]),
        .I5(_inferred__1_carry_i_6__0_n_0),
        .O(\r_c[5]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[5]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [2]),
        .I1(\r_c[1]_i_3__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [0]),
        .I3(_inferred__1_carry_i_7__1_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [4]),
        .I5(_inferred__1_carry_i_6__1_n_0),
        .O(\r_c[5]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[5]_i_2__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [2]),
        .I1(\r_c[1]_i_3__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [0]),
        .I3(_inferred__1_carry_i_7__2_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [4]),
        .I5(_inferred__1_carry_i_6__2_n_0),
        .O(\r_c[5]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[5]_i_2__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [2]),
        .I1(\r_c[1]_i_3__3_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [0]),
        .I3(_inferred__1_carry_i_7__3_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [4]),
        .I5(_inferred__1_carry_i_6__3_n_0),
        .O(\r_c[5]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[5]_i_2__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [2]),
        .I1(\r_c[1]_i_3__4_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [0]),
        .I3(_inferred__1_carry_i_7__4_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [4]),
        .I5(_inferred__1_carry_i_6__4_n_0),
        .O(\r_c[5]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[5]_i_2__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [2]),
        .I1(\r_c[1]_i_3__5_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [0]),
        .I3(_inferred__1_carry_i_7__5_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [4]),
        .I5(_inferred__1_carry_i_6__5_n_0),
        .O(\r_c[5]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFCF44FFFFCF77)) 
    \r_c[5]_i_2__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [2]),
        .I1(\r_c[17]_i_3_n_0 ),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [0]),
        .I3(\r_c[18]_i_3_n_0 ),
        .I4(\r_c[20]_i_2__6_n_0 ),
        .I5(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [4]),
        .O(\r_c[5]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[5]_i_2__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [2]),
        .I1(\r_c[1]_i_3__6_n_0 ),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [0]),
        .I3(_inferred__1_carry_i_7__7_n_0),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [4]),
        .I5(_inferred__1_carry_i_6__7_n_0),
        .O(\r_c[5]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[5]_i_2__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [2]),
        .I1(\r_c[1]_i_3__7_n_0 ),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [0]),
        .I3(_inferred__1_carry_i_7__9_n_0),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [4]),
        .I5(_inferred__1_carry_i_6__9_n_0),
        .O(\r_c[5]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[6]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[6]_i_2__6_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[7]_i_2__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC5C0C5CF)) 
    \r_c[6]_i_1__0 
       (.I0(\r_c[7]_i_2_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [7]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I3(\r_c[14]_i_4_n_0 ),
        .I4(\r_c[6]_i_2_n_0 ),
        .O(\r_c[6]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC5C0C5CF)) 
    \r_c[6]_i_1__1 
       (.I0(\r_c[7]_i_2__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [7]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I3(\r_c[14]_i_4__0_n_0 ),
        .I4(\r_c[6]_i_2__0_n_0 ),
        .O(\r_c[6]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC5C0C5CF)) 
    \r_c[6]_i_1__2 
       (.I0(\r_c[7]_i_2__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [7]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I3(\r_c[14]_i_4__1_n_0 ),
        .I4(\r_c[6]_i_2__1_n_0 ),
        .O(\r_c[6]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC5C0C5CF)) 
    \r_c[6]_i_1__3 
       (.I0(\r_c[7]_i_2__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [7]),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I3(\r_c[14]_i_4__2_n_0 ),
        .I4(\r_c[6]_i_2__2_n_0 ),
        .O(\r_c[6]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC5C0C5CF)) 
    \r_c[6]_i_1__4 
       (.I0(\r_c[7]_i_2__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [7]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I3(\r_c[14]_i_4__3_n_0 ),
        .I4(\r_c[6]_i_2__3_n_0 ),
        .O(\r_c[6]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC5C0C5CF)) 
    \r_c[6]_i_1__5 
       (.I0(\r_c[7]_i_2__4_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [7]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I3(\r_c[14]_i_4__4_n_0 ),
        .I4(\r_c[6]_i_2__4_n_0 ),
        .O(\r_c[6]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC5C0C5CF)) 
    \r_c[6]_i_1__6 
       (.I0(\r_c[7]_i_2__5_n_0 ),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [7]),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I3(\r_c[14]_i_4__5_n_0 ),
        .I4(\r_c[6]_i_2__5_n_0 ),
        .O(\r_c[6]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC5C0C5CF)) 
    \r_c[6]_i_1__7 
       (.I0(\r_c[7]_i_2__7_n_0 ),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [7]),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I3(\r_c[14]_i_4__7_n_0 ),
        .I4(\r_c[6]_i_2__7_n_0 ),
        .O(\r_c[6]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC5C0C5CF)) 
    \r_c[6]_i_1__8 
       (.I0(\r_c[7]_i_2__8_n_0 ),
        .I1(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [7]),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I3(\r_c[14]_i_4__8_n_0 ),
        .I4(\r_c[6]_i_2__8_n_0 ),
        .O(\r_c[6]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[6]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [3]),
        .I1(\r_c[1]_i_3_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [1]),
        .I3(_inferred__1_carry_i_7_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [5]),
        .I5(_inferred__1_carry_i_6_n_0),
        .O(\r_c[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[6]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [3]),
        .I1(\r_c[1]_i_3__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [1]),
        .I3(_inferred__1_carry_i_7__0_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [5]),
        .I5(_inferred__1_carry_i_6__0_n_0),
        .O(\r_c[6]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[6]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [3]),
        .I1(\r_c[1]_i_3__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [1]),
        .I3(_inferred__1_carry_i_7__1_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [5]),
        .I5(_inferred__1_carry_i_6__1_n_0),
        .O(\r_c[6]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[6]_i_2__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [3]),
        .I1(\r_c[1]_i_3__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [1]),
        .I3(_inferred__1_carry_i_7__2_n_0),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [5]),
        .I5(_inferred__1_carry_i_6__2_n_0),
        .O(\r_c[6]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[6]_i_2__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [3]),
        .I1(\r_c[1]_i_3__3_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [1]),
        .I3(_inferred__1_carry_i_7__3_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [5]),
        .I5(_inferred__1_carry_i_6__3_n_0),
        .O(\r_c[6]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[6]_i_2__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [3]),
        .I1(\r_c[1]_i_3__4_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [1]),
        .I3(_inferred__1_carry_i_7__4_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [5]),
        .I5(_inferred__1_carry_i_6__4_n_0),
        .O(\r_c[6]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[6]_i_2__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [3]),
        .I1(\r_c[1]_i_3__5_n_0 ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [1]),
        .I3(_inferred__1_carry_i_7__5_n_0),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [5]),
        .I5(_inferred__1_carry_i_6__5_n_0),
        .O(\r_c[6]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFCF44FFFFCF77)) 
    \r_c[6]_i_2__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [3]),
        .I1(\r_c[17]_i_3_n_0 ),
        .I2(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [1]),
        .I3(\r_c[18]_i_3_n_0 ),
        .I4(\r_c[20]_i_2__6_n_0 ),
        .I5(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [5]),
        .O(\r_c[6]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[6]_i_2__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [3]),
        .I1(\r_c[1]_i_3__6_n_0 ),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [1]),
        .I3(_inferred__1_carry_i_7__7_n_0),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [5]),
        .I5(_inferred__1_carry_i_6__7_n_0),
        .O(\r_c[6]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \r_c[6]_i_2__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [3]),
        .I1(\r_c[1]_i_3__7_n_0 ),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [1]),
        .I3(_inferred__1_carry_i_7__9_n_0),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [5]),
        .I5(_inferred__1_carry_i_6__9_n_0),
        .O(\r_c[6]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[7]_i_1 
       (.I0(\r_c[7]_i_2_n_0 ),
        .I1(\r_c[14]_i_4_n_0 ),
        .I2(\r_c[8]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [8]),
        .O(\r_c[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[7]_i_1__0 
       (.I0(\r_c[7]_i_2__0_n_0 ),
        .I1(\r_c[14]_i_4__0_n_0 ),
        .I2(\r_c[8]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [8]),
        .O(\r_c[7]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[7]_i_1__1 
       (.I0(\r_c[7]_i_2__1_n_0 ),
        .I1(\r_c[14]_i_4__1_n_0 ),
        .I2(\r_c[8]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [8]),
        .O(\r_c[7]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[7]_i_1__2 
       (.I0(\r_c[7]_i_2__2_n_0 ),
        .I1(\r_c[14]_i_4__2_n_0 ),
        .I2(\r_c[8]_i_2__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [8]),
        .O(\r_c[7]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[7]_i_1__3 
       (.I0(\r_c[7]_i_2__3_n_0 ),
        .I1(\r_c[14]_i_4__3_n_0 ),
        .I2(\r_c[8]_i_2__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [8]),
        .O(\r_c[7]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[7]_i_1__4 
       (.I0(\r_c[7]_i_2__4_n_0 ),
        .I1(\r_c[14]_i_4__4_n_0 ),
        .I2(\r_c[8]_i_2__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [8]),
        .O(\r_c[7]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[7]_i_1__5 
       (.I0(\r_c[7]_i_2__5_n_0 ),
        .I1(\r_c[14]_i_4__5_n_0 ),
        .I2(\r_c[8]_i_2__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [8]),
        .O(\r_c[7]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[7]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[7]_i_2__6_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[8]_i_2__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[7]_i_1__7 
       (.I0(\r_c[7]_i_2__7_n_0 ),
        .I1(\r_c[14]_i_4__7_n_0 ),
        .I2(\r_c[8]_i_2__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [8]),
        .O(\r_c[7]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[7]_i_1__8 
       (.I0(\r_c[7]_i_2__8_n_0 ),
        .I1(\r_c[14]_i_4__8_n_0 ),
        .I2(\r_c[8]_i_2__8_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [8]),
        .O(\r_c[7]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[7]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [0]),
        .I1(_inferred__1_carry_i_7_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [4]),
        .I3(_inferred__1_carry_i_6_n_0),
        .I4(\r_c[1]_i_3_n_0 ),
        .I5(\r_c[7]_i_3_n_0 ),
        .O(\r_c[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[7]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [0]),
        .I1(_inferred__1_carry_i_7__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [4]),
        .I3(_inferred__1_carry_i_6__0_n_0),
        .I4(\r_c[1]_i_3__0_n_0 ),
        .I5(\r_c[7]_i_3__0_n_0 ),
        .O(\r_c[7]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[7]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [0]),
        .I1(_inferred__1_carry_i_7__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [4]),
        .I3(_inferred__1_carry_i_6__1_n_0),
        .I4(\r_c[1]_i_3__1_n_0 ),
        .I5(\r_c[7]_i_3__1_n_0 ),
        .O(\r_c[7]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[7]_i_2__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [0]),
        .I1(_inferred__1_carry_i_7__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [4]),
        .I3(_inferred__1_carry_i_6__2_n_0),
        .I4(\r_c[1]_i_3__2_n_0 ),
        .I5(\r_c[7]_i_3__2_n_0 ),
        .O(\r_c[7]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[7]_i_2__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [0]),
        .I1(_inferred__1_carry_i_7__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [4]),
        .I3(_inferred__1_carry_i_6__3_n_0),
        .I4(\r_c[1]_i_3__3_n_0 ),
        .I5(\r_c[7]_i_3__3_n_0 ),
        .O(\r_c[7]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[7]_i_2__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [0]),
        .I1(_inferred__1_carry_i_7__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [4]),
        .I3(_inferred__1_carry_i_6__4_n_0),
        .I4(\r_c[1]_i_3__4_n_0 ),
        .I5(\r_c[7]_i_3__4_n_0 ),
        .O(\r_c[7]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[7]_i_2__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [0]),
        .I1(_inferred__1_carry_i_7__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [4]),
        .I3(_inferred__1_carry_i_6__5_n_0),
        .I4(\r_c[1]_i_3__5_n_0 ),
        .I5(\r_c[7]_i_3__5_n_0 ),
        .O(\r_c[7]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \r_c[7]_i_2__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [0]),
        .I1(\r_c[18]_i_3_n_0 ),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [4]),
        .I4(\r_c[17]_i_3_n_0 ),
        .I5(\r_c[7]_i_3__6_n_0 ),
        .O(\r_c[7]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[7]_i_2__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [0]),
        .I1(_inferred__1_carry_i_7__7_n_0),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [4]),
        .I3(_inferred__1_carry_i_6__7_n_0),
        .I4(\r_c[1]_i_3__6_n_0 ),
        .I5(\r_c[7]_i_3__7_n_0 ),
        .O(\r_c[7]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[7]_i_2__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [0]),
        .I1(_inferred__1_carry_i_7__9_n_0),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [4]),
        .I3(_inferred__1_carry_i_6__9_n_0),
        .I4(\r_c[1]_i_3__7_n_0 ),
        .I5(\r_c[7]_i_3__8_n_0 ),
        .O(\r_c[7]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[7]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [2]),
        .I1(_inferred__1_carry_i_7_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [6]),
        .I3(_inferred__1_carry_i_6_n_0),
        .O(\r_c[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[7]_i_3__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [2]),
        .I1(_inferred__1_carry_i_7__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [6]),
        .I3(_inferred__1_carry_i_6__0_n_0),
        .O(\r_c[7]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[7]_i_3__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [2]),
        .I1(_inferred__1_carry_i_7__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [6]),
        .I3(_inferred__1_carry_i_6__1_n_0),
        .O(\r_c[7]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[7]_i_3__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [2]),
        .I1(_inferred__1_carry_i_7__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [6]),
        .I3(_inferred__1_carry_i_6__2_n_0),
        .O(\r_c[7]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[7]_i_3__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [2]),
        .I1(_inferred__1_carry_i_7__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [6]),
        .I3(_inferred__1_carry_i_6__3_n_0),
        .O(\r_c[7]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[7]_i_3__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [2]),
        .I1(_inferred__1_carry_i_7__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [6]),
        .I3(_inferred__1_carry_i_6__4_n_0),
        .O(\r_c[7]_i_3__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[7]_i_3__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [2]),
        .I1(_inferred__1_carry_i_7__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [6]),
        .I3(_inferred__1_carry_i_6__5_n_0),
        .O(\r_c[7]_i_3__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \r_c[7]_i_3__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [2]),
        .I1(\r_c[18]_i_3_n_0 ),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [6]),
        .O(\r_c[7]_i_3__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[7]_i_3__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [2]),
        .I1(_inferred__1_carry_i_7__7_n_0),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [6]),
        .I3(_inferred__1_carry_i_6__7_n_0),
        .O(\r_c[7]_i_3__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[7]_i_3__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [2]),
        .I1(_inferred__1_carry_i_7__9_n_0),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [6]),
        .I3(_inferred__1_carry_i_6__9_n_0),
        .O(\r_c[7]_i_3__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[8]_i_1 
       (.I0(\r_c[8]_i_2_n_0 ),
        .I1(\r_c[14]_i_4_n_0 ),
        .I2(\r_c[9]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [9]),
        .O(\r_c[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[8]_i_1__0 
       (.I0(\r_c[8]_i_2__0_n_0 ),
        .I1(\r_c[14]_i_4__0_n_0 ),
        .I2(\r_c[9]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [9]),
        .O(\r_c[8]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[8]_i_1__1 
       (.I0(\r_c[8]_i_2__1_n_0 ),
        .I1(\r_c[14]_i_4__1_n_0 ),
        .I2(\r_c[9]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [9]),
        .O(\r_c[8]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[8]_i_1__2 
       (.I0(\r_c[8]_i_2__2_n_0 ),
        .I1(\r_c[14]_i_4__2_n_0 ),
        .I2(\r_c[9]_i_2__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [9]),
        .O(\r_c[8]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[8]_i_1__3 
       (.I0(\r_c[8]_i_2__3_n_0 ),
        .I1(\r_c[14]_i_4__3_n_0 ),
        .I2(\r_c[9]_i_2__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [9]),
        .O(\r_c[8]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[8]_i_1__4 
       (.I0(\r_c[8]_i_2__4_n_0 ),
        .I1(\r_c[14]_i_4__4_n_0 ),
        .I2(\r_c[9]_i_2__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [9]),
        .O(\r_c[8]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[8]_i_1__5 
       (.I0(\r_c[8]_i_2__5_n_0 ),
        .I1(\r_c[14]_i_4__5_n_0 ),
        .I2(\r_c[9]_i_2__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [9]),
        .O(\r_c[8]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[8]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[8]_i_2__6_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[9]_i_2__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[8]_i_1__7 
       (.I0(\r_c[8]_i_2__7_n_0 ),
        .I1(\r_c[14]_i_4__7_n_0 ),
        .I2(\r_c[9]_i_2__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [9]),
        .O(\r_c[8]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[8]_i_1__8 
       (.I0(\r_c[8]_i_2__8_n_0 ),
        .I1(\r_c[14]_i_4__8_n_0 ),
        .I2(\r_c[9]_i_2__8_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [9]),
        .O(\r_c[8]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[8]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [1]),
        .I1(_inferred__1_carry_i_7_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [5]),
        .I3(_inferred__1_carry_i_6_n_0),
        .I4(\r_c[1]_i_3_n_0 ),
        .I5(\r_c[8]_i_3_n_0 ),
        .O(\r_c[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[8]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [1]),
        .I1(_inferred__1_carry_i_7__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [5]),
        .I3(_inferred__1_carry_i_6__0_n_0),
        .I4(\r_c[1]_i_3__0_n_0 ),
        .I5(\r_c[8]_i_3__0_n_0 ),
        .O(\r_c[8]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[8]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [1]),
        .I1(_inferred__1_carry_i_7__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [5]),
        .I3(_inferred__1_carry_i_6__1_n_0),
        .I4(\r_c[1]_i_3__1_n_0 ),
        .I5(\r_c[8]_i_3__1_n_0 ),
        .O(\r_c[8]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[8]_i_2__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [1]),
        .I1(_inferred__1_carry_i_7__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [5]),
        .I3(_inferred__1_carry_i_6__2_n_0),
        .I4(\r_c[1]_i_3__2_n_0 ),
        .I5(\r_c[8]_i_3__2_n_0 ),
        .O(\r_c[8]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[8]_i_2__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [1]),
        .I1(_inferred__1_carry_i_7__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [5]),
        .I3(_inferred__1_carry_i_6__3_n_0),
        .I4(\r_c[1]_i_3__3_n_0 ),
        .I5(\r_c[8]_i_3__3_n_0 ),
        .O(\r_c[8]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[8]_i_2__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [1]),
        .I1(_inferred__1_carry_i_7__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [5]),
        .I3(_inferred__1_carry_i_6__4_n_0),
        .I4(\r_c[1]_i_3__4_n_0 ),
        .I5(\r_c[8]_i_3__4_n_0 ),
        .O(\r_c[8]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[8]_i_2__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [1]),
        .I1(_inferred__1_carry_i_7__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [5]),
        .I3(_inferred__1_carry_i_6__5_n_0),
        .I4(\r_c[1]_i_3__5_n_0 ),
        .I5(\r_c[8]_i_3__5_n_0 ),
        .O(\r_c[8]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \r_c[8]_i_2__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [1]),
        .I1(\r_c[18]_i_3_n_0 ),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [5]),
        .I4(\r_c[17]_i_3_n_0 ),
        .I5(\r_c[8]_i_3__6_n_0 ),
        .O(\r_c[8]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[8]_i_2__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [1]),
        .I1(_inferred__1_carry_i_7__7_n_0),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [5]),
        .I3(_inferred__1_carry_i_6__7_n_0),
        .I4(\r_c[1]_i_3__6_n_0 ),
        .I5(\r_c[8]_i_3__7_n_0 ),
        .O(\r_c[8]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[8]_i_2__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [1]),
        .I1(_inferred__1_carry_i_7__9_n_0),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [5]),
        .I3(_inferred__1_carry_i_6__9_n_0),
        .I4(\r_c[1]_i_3__7_n_0 ),
        .I5(\r_c[8]_i_3__8_n_0 ),
        .O(\r_c[8]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[8]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [3]),
        .I1(_inferred__1_carry_i_7_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [7]),
        .I3(_inferred__1_carry_i_6_n_0),
        .O(\r_c[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[8]_i_3__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [3]),
        .I1(_inferred__1_carry_i_7__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [7]),
        .I3(_inferred__1_carry_i_6__0_n_0),
        .O(\r_c[8]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[8]_i_3__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [3]),
        .I1(_inferred__1_carry_i_7__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [7]),
        .I3(_inferred__1_carry_i_6__1_n_0),
        .O(\r_c[8]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[8]_i_3__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [3]),
        .I1(_inferred__1_carry_i_7__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [7]),
        .I3(_inferred__1_carry_i_6__2_n_0),
        .O(\r_c[8]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[8]_i_3__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [3]),
        .I1(_inferred__1_carry_i_7__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [7]),
        .I3(_inferred__1_carry_i_6__3_n_0),
        .O(\r_c[8]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[8]_i_3__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [3]),
        .I1(_inferred__1_carry_i_7__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [7]),
        .I3(_inferred__1_carry_i_6__4_n_0),
        .O(\r_c[8]_i_3__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[8]_i_3__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [3]),
        .I1(_inferred__1_carry_i_7__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [7]),
        .I3(_inferred__1_carry_i_6__5_n_0),
        .O(\r_c[8]_i_3__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \r_c[8]_i_3__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [3]),
        .I1(\r_c[18]_i_3_n_0 ),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [7]),
        .O(\r_c[8]_i_3__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[8]_i_3__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [3]),
        .I1(_inferred__1_carry_i_7__7_n_0),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [7]),
        .I3(_inferred__1_carry_i_6__7_n_0),
        .O(\r_c[8]_i_3__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    \r_c[8]_i_3__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [3]),
        .I1(_inferred__1_carry_i_7__9_n_0),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [7]),
        .I3(_inferred__1_carry_i_6__9_n_0),
        .O(\r_c[8]_i_3__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[9]_i_1 
       (.I0(\r_c[9]_i_2_n_0 ),
        .I1(\r_c[14]_i_4_n_0 ),
        .I2(\r_c[10]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [10]),
        .O(\r_c[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[9]_i_1__0 
       (.I0(\r_c[9]_i_2__0_n_0 ),
        .I1(\r_c[14]_i_4__0_n_0 ),
        .I2(\r_c[10]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [10]),
        .O(\r_c[9]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[9]_i_1__1 
       (.I0(\r_c[9]_i_2__1_n_0 ),
        .I1(\r_c[14]_i_4__1_n_0 ),
        .I2(\r_c[10]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [10]),
        .O(\r_c[9]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[9]_i_1__2 
       (.I0(\r_c[9]_i_2__2_n_0 ),
        .I1(\r_c[14]_i_4__2_n_0 ),
        .I2(\r_c[10]_i_2__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [10]),
        .O(\r_c[9]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[9]_i_1__3 
       (.I0(\r_c[9]_i_2__3_n_0 ),
        .I1(\r_c[14]_i_4__3_n_0 ),
        .I2(\r_c[10]_i_2__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [10]),
        .O(\r_c[9]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[9]_i_1__4 
       (.I0(\r_c[9]_i_2__4_n_0 ),
        .I1(\r_c[14]_i_4__4_n_0 ),
        .I2(\r_c[10]_i_2__4_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [10]),
        .O(\r_c[9]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[9]_i_1__5 
       (.I0(\r_c[9]_i_2__5_n_0 ),
        .I1(\r_c[14]_i_4__5_n_0 ),
        .I2(\r_c[10]_i_2__5_n_0 ),
        .I3(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .I4(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [10]),
        .O(\r_c[9]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FEFEFE00FE)) 
    \r_c[9]_i_1__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .I2(\r_c[14]_i_2__6_n_0 ),
        .I3(\r_c[9]_i_2__6_n_0 ),
        .I4(\r_c[17]_i_2_n_0 ),
        .I5(\r_c[10]_i_2__6_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_c [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[9]_i_1__7 
       (.I0(\r_c[9]_i_2__7_n_0 ),
        .I1(\r_c[14]_i_4__7_n_0 ),
        .I2(\r_c[10]_i_2__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [10]),
        .O(\r_c[9]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF1D001D)) 
    \r_c[9]_i_1__8 
       (.I0(\r_c[9]_i_2__8_n_0 ),
        .I1(\r_c[14]_i_4__8_n_0 ),
        .I2(\r_c[10]_i_2__8_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .I4(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [10]),
        .O(\r_c[9]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[9]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [2]),
        .I1(_inferred__1_carry_i_7_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [6]),
        .I3(_inferred__1_carry_i_6_n_0),
        .I4(\r_c[1]_i_3_n_0 ),
        .I5(\r_c[11]_i_3_n_0 ),
        .O(\r_c[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[9]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [2]),
        .I1(_inferred__1_carry_i_7__0_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [6]),
        .I3(_inferred__1_carry_i_6__0_n_0),
        .I4(\r_c[1]_i_3__0_n_0 ),
        .I5(\r_c[11]_i_3__0_n_0 ),
        .O(\r_c[9]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[9]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [2]),
        .I1(_inferred__1_carry_i_7__1_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [6]),
        .I3(_inferred__1_carry_i_6__1_n_0),
        .I4(\r_c[1]_i_3__1_n_0 ),
        .I5(\r_c[11]_i_3__1_n_0 ),
        .O(\r_c[9]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[9]_i_2__2 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [2]),
        .I1(_inferred__1_carry_i_7__2_n_0),
        .I2(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [6]),
        .I3(_inferred__1_carry_i_6__2_n_0),
        .I4(\r_c[1]_i_3__2_n_0 ),
        .I5(\r_c[11]_i_3__2_n_0 ),
        .O(\r_c[9]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[9]_i_2__3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [2]),
        .I1(_inferred__1_carry_i_7__3_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [6]),
        .I3(_inferred__1_carry_i_6__3_n_0),
        .I4(\r_c[1]_i_3__3_n_0 ),
        .I5(\r_c[11]_i_3__3_n_0 ),
        .O(\r_c[9]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[9]_i_2__4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [2]),
        .I1(_inferred__1_carry_i_7__4_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [6]),
        .I3(_inferred__1_carry_i_6__4_n_0),
        .I4(\r_c[1]_i_3__4_n_0 ),
        .I5(\r_c[11]_i_3__4_n_0 ),
        .O(\r_c[9]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[9]_i_2__5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [2]),
        .I1(_inferred__1_carry_i_7__5_n_0),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [6]),
        .I3(_inferred__1_carry_i_6__5_n_0),
        .I4(\r_c[1]_i_3__5_n_0 ),
        .I5(\r_c[11]_i_3__5_n_0 ),
        .O(\r_c[9]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \r_c[9]_i_2__6 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [2]),
        .I1(\r_c[18]_i_3_n_0 ),
        .I2(\r_c[20]_i_2__6_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [6]),
        .I4(\r_c[17]_i_3_n_0 ),
        .I5(\r_c[11]_i_3__6_n_0 ),
        .O(\r_c[9]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[9]_i_2__7 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [2]),
        .I1(_inferred__1_carry_i_7__7_n_0),
        .I2(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [6]),
        .I3(_inferred__1_carry_i_6__7_n_0),
        .I4(\r_c[1]_i_3__6_n_0 ),
        .I5(\r_c[11]_i_3__7_n_0 ),
        .O(\r_c[9]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    \r_c[9]_i_2__8 
       (.I0(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [2]),
        .I1(_inferred__1_carry_i_7__9_n_0),
        .I2(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [6]),
        .I3(_inferred__1_carry_i_6__9_n_0),
        .I4(\r_c[1]_i_3__7_n_0 ),
        .I5(\r_c[11]_i_3__8_n_0 ),
        .O(\r_c[9]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBF80)) 
    r_ccw_i_1
       (.I0(s_wb_dat_i[16]),
        .I1(r_dma_start_i_2_n_0),
        .I2(s_wb_sel_i[2]),
        .I3(w_ccw),
        .O(r_ccw_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r_ce_tmp[1]_i_1 
       (.I0(\u_geo/w_vw_clip [16]),
        .I1(\u_geo/w_vw_clip [17]),
        .O(r_ce_tmp));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT3 #(
    .INIT(8'h87)) 
    \r_ce_tmp[2]_i_1 
       (.I0(\u_geo/w_vw_clip [17]),
        .I1(\u_geo/w_vw_clip [16]),
        .I2(\u_geo/w_vw_clip [18]),
        .O(\r_ce_tmp[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT4 #(
    .INIT(16'h807F)) 
    \r_ce_tmp[3]_i_1 
       (.I0(\u_geo/w_vw_clip [18]),
        .I1(\u_geo/w_vw_clip [16]),
        .I2(\u_geo/w_vw_clip [17]),
        .I3(\u_geo/w_vw_clip [19]),
        .O(\r_ce_tmp[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT5 #(
    .INIT(32'h80007FFF)) 
    \r_ce_tmp[4]_i_1 
       (.I0(\u_geo/w_vw_clip [19]),
        .I1(\u_geo/w_vw_clip [17]),
        .I2(\u_geo/w_vw_clip [16]),
        .I3(\u_geo/w_vw_clip [18]),
        .I4(\u_geo/w_vw_clip [20]),
        .O(\r_ce_tmp[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFA959)) 
    \r_ce_tmp_1z[0]_i_1 
       (.I0(\r_ce_tmp_1z[0]_i_2_n_0 ),
        .I1(\u_geo/u_geo_matrix/r_vx_in [16]),
        .I2(\u_geo/w_state_mat ),
        .I3(\u_geo/w_vx_dma [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m0/w_adder_out ),
        .O(\r_ce_tmp_1z[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFA959)) 
    \r_ce_tmp_1z[0]_i_1__0 
       (.I0(\r_ce_tmp_1z[0]_i_2__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/r_vy_in [16]),
        .I2(\u_geo/w_state_mat ),
        .I3(\u_geo/w_vy_dma [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m1/w_adder_out ),
        .O(r_ce_tmp_1z));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFA959)) 
    \r_ce_tmp_1z[0]_i_1__1 
       (.I0(\r_ce_tmp_1z[0]_i_2__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/r_vz_in [16]),
        .I2(\u_geo/w_state_mat ),
        .I3(\u_geo/w_vz_dma [16]),
        .I4(\u_geo/u_geo_matrix/u_fmul_m2/w_adder_out ),
        .O(\r_ce_tmp_1z[0]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[0]_i_1__2 
       (.I0(w_m13[16]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[0]_i_2__2_n_0 ),
        .O(\r_ce_tmp_1z[0]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[0]_i_2 
       (.I0(w_m10[16]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[1]_i_5_n_0 ),
        .O(\r_ce_tmp_1z[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[0]_i_2__0 
       (.I0(w_m11[16]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[1]_i_5__0_n_0 ),
        .O(\r_ce_tmp_1z[0]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[0]_i_2__1 
       (.I0(w_m12[16]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[1]_i_5__1_n_0 ),
        .O(\r_ce_tmp_1z[0]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[0]_i_2__2 
       (.I0(w_m23[16]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[16]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[16]),
        .O(\r_ce_tmp_1z[0]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF47B8B847)) 
    \r_ce_tmp_1z[1]_i_1 
       (.I0(\u_geo/w_vx_dma [17]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [17]),
        .I3(\r_ce_tmp_1z[1]_i_2_n_0 ),
        .I4(\r_ce_tmp_1z[1]_i_3_n_0 ),
        .I5(\u_geo/u_geo_matrix/u_fmul_m0/w_adder_out ),
        .O(\r_ce_tmp_1z[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF47B8B847)) 
    \r_ce_tmp_1z[1]_i_1__0 
       (.I0(\u_geo/w_vy_dma [17]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [17]),
        .I3(\r_ce_tmp_1z[1]_i_2__0_n_0 ),
        .I4(\r_ce_tmp_1z[1]_i_3__0_n_0 ),
        .I5(\u_geo/u_geo_matrix/u_fmul_m1/w_adder_out ),
        .O(\r_ce_tmp_1z[1]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF47B8B847)) 
    \r_ce_tmp_1z[1]_i_1__1 
       (.I0(\u_geo/w_vz_dma [17]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [17]),
        .I3(\r_ce_tmp_1z[1]_i_2__1_n_0 ),
        .I4(\r_ce_tmp_1z[1]_i_3__1_n_0 ),
        .I5(\u_geo/u_geo_matrix/u_fmul_m2/w_adder_out ),
        .O(\r_ce_tmp_1z[1]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[1]_i_1__2 
       (.I0(w_m13[17]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[1]_i_2__2_n_0 ),
        .O(\r_ce_tmp_1z[1]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[1]_i_2 
       (.I0(w_m10[17]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[1]_i_4_n_0 ),
        .O(\r_ce_tmp_1z[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[1]_i_2__0 
       (.I0(w_m11[17]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[1]_i_4__0_n_0 ),
        .O(\r_ce_tmp_1z[1]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[1]_i_2__1 
       (.I0(w_m12[17]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[1]_i_4__1_n_0 ),
        .O(\r_ce_tmp_1z[1]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[1]_i_2__2 
       (.I0(w_m23[17]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[17]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[17]),
        .O(\r_ce_tmp_1z[1]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFB8B8B8FFB8)) 
    \r_ce_tmp_1z[1]_i_2__3 
       (.I0(\u_geo/w_vx_pdiv [16]),
        .I1(\r_ce_tmp_1z[4]_i_3__2_n_0 ),
        .I2(\u_geo/w_vy_pdiv [16]),
        .I3(\u_geo/u_geo_persdiv/r_ivw [16]),
        .I4(r_ivw),
        .I5(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[16] ),
        .O(\r_ce_tmp_1z[1]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h001B)) 
    \r_ce_tmp_1z[1]_i_2__4 
       (.I0(\r_ce_tmp_1z[4]_i_3__3_n_0 ),
        .I1(w_vh[16]),
        .I2(w_vw[16]),
        .I3(\u_geo/u_geo_viewport/w_a_exp [0]),
        .O(\r_ce_tmp_1z[1]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000001D1D1D001D)) 
    \r_ce_tmp_1z[1]_i_3 
       (.I0(\r_ce_tmp_1z[1]_i_5_n_0 ),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_m10[16]),
        .I3(\u_geo/u_geo_matrix/r_vx_in [16]),
        .I4(\u_geo/w_state_mat ),
        .I5(\u_geo/w_vx_dma [16]),
        .O(\r_ce_tmp_1z[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000001D1D1D001D)) 
    \r_ce_tmp_1z[1]_i_3__0 
       (.I0(\r_ce_tmp_1z[1]_i_5__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_m11[16]),
        .I3(\u_geo/u_geo_matrix/r_vy_in [16]),
        .I4(\u_geo/w_state_mat ),
        .I5(\u_geo/w_vy_dma [16]),
        .O(\r_ce_tmp_1z[1]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000001D1D1D001D)) 
    \r_ce_tmp_1z[1]_i_3__1 
       (.I0(\r_ce_tmp_1z[1]_i_5__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_m12[16]),
        .I3(\u_geo/u_geo_matrix/r_vz_in [16]),
        .I4(\u_geo/w_state_mat ),
        .I5(\u_geo/w_vz_dma [16]),
        .O(\r_ce_tmp_1z[1]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[1]_i_4 
       (.I0(w_m20[17]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[17]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[17]),
        .O(\r_ce_tmp_1z[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[1]_i_4__0 
       (.I0(w_m21[17]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[17]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[17]),
        .O(\r_ce_tmp_1z[1]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[1]_i_4__1 
       (.I0(w_m22[17]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[17]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[17]),
        .O(\r_ce_tmp_1z[1]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[1]_i_5 
       (.I0(w_m20[16]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[16]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[16]),
        .O(\r_ce_tmp_1z[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[1]_i_5__0 
       (.I0(w_m21[16]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[16]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[16]),
        .O(\r_ce_tmp_1z[1]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[1]_i_5__1 
       (.I0(w_m22[16]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[16]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[16]),
        .O(\r_ce_tmp_1z[1]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFA95956A6)) 
    \r_ce_tmp_1z[2]_i_1 
       (.I0(\r_ce_tmp_1z[2]_i_2_n_0 ),
        .I1(\u_geo/u_geo_matrix/r_vx_in [18]),
        .I2(\u_geo/w_state_mat ),
        .I3(\u_geo/w_vx_dma [18]),
        .I4(\r_ce_tmp_1z[2]_i_3_n_0 ),
        .I5(\u_geo/u_geo_matrix/u_fmul_m0/w_adder_out ),
        .O(\r_ce_tmp_1z[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFA95956A6)) 
    \r_ce_tmp_1z[2]_i_1__0 
       (.I0(\r_ce_tmp_1z[2]_i_2__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/r_vy_in [18]),
        .I2(\u_geo/w_state_mat ),
        .I3(\u_geo/w_vy_dma [18]),
        .I4(\r_ce_tmp_1z[2]_i_3__0_n_0 ),
        .I5(\u_geo/u_geo_matrix/u_fmul_m1/w_adder_out ),
        .O(\r_ce_tmp_1z[2]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFA95956A6)) 
    \r_ce_tmp_1z[2]_i_1__1 
       (.I0(\r_ce_tmp_1z[2]_i_2__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/r_vz_in [18]),
        .I2(\u_geo/w_state_mat ),
        .I3(\u_geo/w_vz_dma [18]),
        .I4(\r_ce_tmp_1z[2]_i_3__1_n_0 ),
        .I5(\u_geo/u_geo_matrix/u_fmul_m2/w_adder_out ),
        .O(\r_ce_tmp_1z[2]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[2]_i_1__2 
       (.I0(w_m13[18]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[2]_i_2__2_n_0 ),
        .O(\r_ce_tmp_1z[2]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDDD444D4)) 
    \r_ce_tmp_1z[2]_i_2 
       (.I0(\r_ce_tmp_1z[1]_i_3_n_0 ),
        .I1(\r_ce_tmp_1z[1]_i_2_n_0 ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [17]),
        .I3(\u_geo/w_state_mat ),
        .I4(\u_geo/w_vx_dma [17]),
        .O(\r_ce_tmp_1z[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDDD444D4)) 
    \r_ce_tmp_1z[2]_i_2__0 
       (.I0(\r_ce_tmp_1z[1]_i_3__0_n_0 ),
        .I1(\r_ce_tmp_1z[1]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [17]),
        .I3(\u_geo/w_state_mat ),
        .I4(\u_geo/w_vy_dma [17]),
        .O(\r_ce_tmp_1z[2]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDDD444D4)) 
    \r_ce_tmp_1z[2]_i_2__1 
       (.I0(\r_ce_tmp_1z[1]_i_3__1_n_0 ),
        .I1(\r_ce_tmp_1z[1]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [17]),
        .I3(\u_geo/w_state_mat ),
        .I4(\u_geo/w_vz_dma [17]),
        .O(\r_ce_tmp_1z[2]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[2]_i_2__2 
       (.I0(w_m23[18]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[18]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[18]),
        .O(\r_ce_tmp_1z[2]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h1015757F)) 
    \r_ce_tmp_1z[2]_i_2__3 
       (.I0(\r_ce_tmp_1z[1]_i_2__3_n_0 ),
        .I1(\u_geo/w_vx_pdiv [17]),
        .I2(\r_ce_tmp_1z[4]_i_3__2_n_0 ),
        .I3(\u_geo/w_vy_pdiv [17]),
        .I4(\u_geo/u_geo_persdiv/w_b_exp [1]),
        .O(\r_ce_tmp_1z[2]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFD755410)) 
    \r_ce_tmp_1z[2]_i_2__4 
       (.I0(\r_ce_tmp_1z[1]_i_2__4_n_0 ),
        .I1(\r_ce_tmp_1z[4]_i_3__3_n_0 ),
        .I2(w_vh[17]),
        .I3(w_vw[17]),
        .I4(\u_geo/u_geo_viewport/w_a_exp [1]),
        .O(\r_ce_tmp_1z[2]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[2]_i_3 
       (.I0(w_m10[18]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[2]_i_4_n_0 ),
        .O(\r_ce_tmp_1z[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[2]_i_3__0 
       (.I0(w_m11[18]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[2]_i_4__0_n_0 ),
        .O(\r_ce_tmp_1z[2]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[2]_i_3__1 
       (.I0(w_m12[18]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[2]_i_4__1_n_0 ),
        .O(\r_ce_tmp_1z[2]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[2]_i_4 
       (.I0(w_m20[18]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[18]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[18]),
        .O(\r_ce_tmp_1z[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[2]_i_4__0 
       (.I0(w_m21[18]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[18]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[18]),
        .O(\r_ce_tmp_1z[2]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[2]_i_4__1 
       (.I0(w_m22[18]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[18]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[18]),
        .O(\r_ce_tmp_1z[2]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF99966696)) 
    \r_ce_tmp_1z[3]_i_1 
       (.I0(\r_ce_tmp_1z[3]_i_2_n_0 ),
        .I1(\r_ce_tmp_1z[3]_i_3_n_0 ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [19]),
        .I3(\u_geo/w_state_mat ),
        .I4(\u_geo/w_vx_dma [19]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m0/w_adder_out ),
        .O(\r_ce_tmp_1z[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF99966696)) 
    \r_ce_tmp_1z[3]_i_1__0 
       (.I0(\r_ce_tmp_1z[3]_i_2__0_n_0 ),
        .I1(\r_ce_tmp_1z[3]_i_3__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [19]),
        .I3(\u_geo/w_state_mat ),
        .I4(\u_geo/w_vy_dma [19]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m1/w_adder_out ),
        .O(\r_ce_tmp_1z[3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF99966696)) 
    \r_ce_tmp_1z[3]_i_1__1 
       (.I0(\r_ce_tmp_1z[3]_i_2__1_n_0 ),
        .I1(\r_ce_tmp_1z[3]_i_3__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [19]),
        .I3(\u_geo/w_state_mat ),
        .I4(\u_geo/w_vz_dma [19]),
        .I5(\u_geo/u_geo_matrix/u_fmul_m2/w_adder_out ),
        .O(\r_ce_tmp_1z[3]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[3]_i_1__2 
       (.I0(w_m13[19]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[3]_i_2__2_n_0 ),
        .O(\r_ce_tmp_1z[3]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFEAEA808)) 
    \r_ce_tmp_1z[3]_i_2 
       (.I0(\r_ce_tmp_1z[2]_i_2_n_0 ),
        .I1(\u_geo/u_geo_matrix/r_vx_in [18]),
        .I2(\u_geo/w_state_mat ),
        .I3(\u_geo/w_vx_dma [18]),
        .I4(\r_ce_tmp_1z[2]_i_3_n_0 ),
        .O(\r_ce_tmp_1z[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFEAEA808)) 
    \r_ce_tmp_1z[3]_i_2__0 
       (.I0(\r_ce_tmp_1z[2]_i_2__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/r_vy_in [18]),
        .I2(\u_geo/w_state_mat ),
        .I3(\u_geo/w_vy_dma [18]),
        .I4(\r_ce_tmp_1z[2]_i_3__0_n_0 ),
        .O(\r_ce_tmp_1z[3]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFEAEA808)) 
    \r_ce_tmp_1z[3]_i_2__1 
       (.I0(\r_ce_tmp_1z[2]_i_2__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/r_vz_in [18]),
        .I2(\u_geo/w_state_mat ),
        .I3(\u_geo/w_vz_dma [18]),
        .I4(\r_ce_tmp_1z[2]_i_3__1_n_0 ),
        .O(\r_ce_tmp_1z[3]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[3]_i_2__2 
       (.I0(w_m23[19]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[19]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[19]),
        .O(\r_ce_tmp_1z[3]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h202ABABF)) 
    \r_ce_tmp_1z[3]_i_2__3 
       (.I0(\r_ce_tmp_1z[2]_i_2__3_n_0 ),
        .I1(\u_geo/w_vx_pdiv [18]),
        .I2(\r_ce_tmp_1z[4]_i_3__2_n_0 ),
        .I3(\u_geo/w_vy_pdiv [18]),
        .I4(\u_geo/u_geo_persdiv/w_b_exp [2]),
        .O(\r_ce_tmp_1z[3]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEE88E88)) 
    \r_ce_tmp_1z[3]_i_2__4 
       (.I0(\r_ce_tmp_1z[2]_i_2__4_n_0 ),
        .I1(\u_geo/u_geo_viewport/w_a_exp [2]),
        .I2(\r_ce_tmp_1z[4]_i_3__3_n_0 ),
        .I3(w_vh[18]),
        .I4(w_vw[18]),
        .O(\r_ce_tmp_1z[3]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[3]_i_3 
       (.I0(w_m10[19]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[3]_i_5_n_0 ),
        .O(\r_ce_tmp_1z[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[3]_i_3__0 
       (.I0(w_m11[19]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[3]_i_5__0_n_0 ),
        .O(\r_ce_tmp_1z[3]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[3]_i_3__1 
       (.I0(w_m12[19]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[3]_i_5__1_n_0 ),
        .O(\r_ce_tmp_1z[3]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h42444222)) 
    \r_ce_tmp_1z[3]_i_3__2 
       (.I0(\r_ce_tmp_1z[4]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_persdiv/w_b_exp [4]),
        .I2(\u_geo/w_vx_pdiv [20]),
        .I3(\r_ce_tmp_1z[4]_i_3__2_n_0 ),
        .I4(\u_geo/w_vy_pdiv [20]),
        .O(\u_geo/u_geo_persdiv/u_fmul/w_adder_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h5410028A)) 
    \r_ce_tmp_1z[3]_i_3__3 
       (.I0(\r_ce_tmp_1z[4]_i_4__3_n_0 ),
        .I1(\r_ce_tmp_1z[4]_i_3__3_n_0 ),
        .I2(w_vh[20]),
        .I3(w_vw[20]),
        .I4(\u_geo/u_geo_viewport/w_a_exp [4]),
        .O(\u_geo/u_geo_viewport/u_fmul/w_adder_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44422242)) 
    \r_ce_tmp_1z[3]_i_4 
       (.I0(\r_ce_tmp_1z[4]_i_4_n_0 ),
        .I1(\r_ce_tmp_1z[4]_i_3_n_0 ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [20]),
        .I3(\u_geo/w_state_mat ),
        .I4(\u_geo/w_vx_dma [20]),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/w_adder_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44422242)) 
    \r_ce_tmp_1z[3]_i_4__0 
       (.I0(\r_ce_tmp_1z[4]_i_4__0_n_0 ),
        .I1(\r_ce_tmp_1z[4]_i_3__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [20]),
        .I3(\u_geo/w_state_mat ),
        .I4(\u_geo/w_vy_dma [20]),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/w_adder_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44422242)) 
    \r_ce_tmp_1z[3]_i_4__1 
       (.I0(\r_ce_tmp_1z[4]_i_4__1_n_0 ),
        .I1(\r_ce_tmp_1z[4]_i_3__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [20]),
        .I3(\u_geo/w_state_mat ),
        .I4(\u_geo/w_vz_dma [20]),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/w_adder_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[3]_i_5 
       (.I0(w_m20[19]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[19]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[19]),
        .O(\r_ce_tmp_1z[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[3]_i_5__0 
       (.I0(w_m21[19]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[19]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[19]),
        .O(\r_ce_tmp_1z[3]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[3]_i_5__1 
       (.I0(w_m22[19]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[19]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[19]),
        .O(\r_ce_tmp_1z[3]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00470000)) 
    \r_ce_tmp_1z[4]_i_1 
       (.I0(\u_geo/w_vx_dma [20]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [20]),
        .I3(\r_ce_tmp_1z[4]_i_3_n_0 ),
        .I4(\r_ce_tmp_1z[4]_i_4_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00470000)) 
    \r_ce_tmp_1z[4]_i_1__0 
       (.I0(\u_geo/w_vy_dma [20]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [20]),
        .I3(\r_ce_tmp_1z[4]_i_3__0_n_0 ),
        .I4(\r_ce_tmp_1z[4]_i_4__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00470000)) 
    \r_ce_tmp_1z[4]_i_1__1 
       (.I0(\u_geo/w_vz_dma [20]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [20]),
        .I3(\r_ce_tmp_1z[4]_i_3__1_n_0 ),
        .I4(\r_ce_tmp_1z[4]_i_4__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[4]_i_1__2 
       (.I0(w_m13[20]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[4]_i_2__2_n_0 ),
        .O(\r_ce_tmp_1z[4]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h01510000)) 
    \r_ce_tmp_1z[4]_i_1__3 
       (.I0(\u_geo/u_geo_persdiv/w_b_exp [4]),
        .I1(\u_geo/w_vy_pdiv [20]),
        .I2(\r_ce_tmp_1z[4]_i_3__2_n_0 ),
        .I3(\u_geo/w_vx_pdiv [20]),
        .I4(\r_ce_tmp_1z[4]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h11050000)) 
    \r_ce_tmp_1z[4]_i_1__4 
       (.I0(\u_geo/u_geo_viewport/w_a_exp [4]),
        .I1(w_vw[20]),
        .I2(w_vh[20]),
        .I3(\r_ce_tmp_1z[4]_i_3__3_n_0 ),
        .I4(\r_ce_tmp_1z[4]_i_4__3_n_0 ),
        .O(\u_geo/u_geo_viewport/u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB847FFB8)) 
    \r_ce_tmp_1z[4]_i_2 
       (.I0(\u_geo/w_vx_dma [20]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [20]),
        .I3(\r_ce_tmp_1z[4]_i_3_n_0 ),
        .I4(\r_ce_tmp_1z[4]_i_4_n_0 ),
        .O(\r_ce_tmp_1z[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB847FFB8)) 
    \r_ce_tmp_1z[4]_i_2__0 
       (.I0(\u_geo/w_vy_dma [20]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [20]),
        .I3(\r_ce_tmp_1z[4]_i_3__0_n_0 ),
        .I4(\r_ce_tmp_1z[4]_i_4__0_n_0 ),
        .O(\r_ce_tmp_1z[4]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB847FFB8)) 
    \r_ce_tmp_1z[4]_i_2__1 
       (.I0(\u_geo/w_vz_dma [20]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [20]),
        .I3(\r_ce_tmp_1z[4]_i_3__1_n_0 ),
        .I4(\r_ce_tmp_1z[4]_i_4__1_n_0 ),
        .O(\r_ce_tmp_1z[4]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[4]_i_2__2 
       (.I0(w_m23[20]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[20]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[20]),
        .O(\r_ce_tmp_1z[4]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[4]_i_3 
       (.I0(w_m10[20]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[4]_i_5_n_0 ),
        .O(\r_ce_tmp_1z[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[4]_i_3__0 
       (.I0(w_m11[20]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[4]_i_5__0_n_0 ),
        .O(\r_ce_tmp_1z[4]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_ce_tmp_1z[4]_i_3__1 
       (.I0(w_m12[20]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_ce_tmp_1z[4]_i_5__1_n_0 ),
        .O(\r_ce_tmp_1z[4]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \r_ce_tmp_1z[4]_i_3__2 
       (.I0(\u_geo/u_geo_persdiv/r_state [0]),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_ce_tmp_1z[4]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1000)) 
    \r_ce_tmp_1z[4]_i_3__3 
       (.I0(\u_geo/u_geo_viewport/r_state [2]),
        .I1(\u_geo/u_geo_viewport/r_state [3]),
        .I2(\u_geo/u_geo_viewport/r_state [1]),
        .I3(\u_geo/u_geo_viewport/r_state [0]),
        .O(\r_ce_tmp_1z[4]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h015157F7)) 
    \r_ce_tmp_1z[4]_i_4 
       (.I0(\r_ce_tmp_1z[3]_i_3_n_0 ),
        .I1(\u_geo/u_geo_matrix/r_vx_in [19]),
        .I2(\u_geo/w_state_mat ),
        .I3(\u_geo/w_vx_dma [19]),
        .I4(\r_ce_tmp_1z[3]_i_2_n_0 ),
        .O(\r_ce_tmp_1z[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h015157F7)) 
    \r_ce_tmp_1z[4]_i_4__0 
       (.I0(\r_ce_tmp_1z[3]_i_3__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/r_vy_in [19]),
        .I2(\u_geo/w_state_mat ),
        .I3(\u_geo/w_vy_dma [19]),
        .I4(\r_ce_tmp_1z[3]_i_2__0_n_0 ),
        .O(\r_ce_tmp_1z[4]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h015157F7)) 
    \r_ce_tmp_1z[4]_i_4__1 
       (.I0(\r_ce_tmp_1z[3]_i_3__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/r_vz_in [19]),
        .I2(\u_geo/w_state_mat ),
        .I3(\u_geo/w_vz_dma [19]),
        .I4(\r_ce_tmp_1z[3]_i_2__1_n_0 ),
        .O(\r_ce_tmp_1z[4]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h202ABABF)) 
    \r_ce_tmp_1z[4]_i_4__2 
       (.I0(\r_ce_tmp_1z[3]_i_2__3_n_0 ),
        .I1(\u_geo/w_vx_pdiv [19]),
        .I2(\r_ce_tmp_1z[4]_i_3__2_n_0 ),
        .I3(\u_geo/w_vy_pdiv [19]),
        .I4(\u_geo/u_geo_persdiv/w_b_exp [3]),
        .O(\r_ce_tmp_1z[4]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h001B1BFF)) 
    \r_ce_tmp_1z[4]_i_4__3 
       (.I0(\r_ce_tmp_1z[4]_i_3__3_n_0 ),
        .I1(w_vh[19]),
        .I2(w_vw[19]),
        .I3(\u_geo/u_geo_viewport/w_a_exp [3]),
        .I4(\r_ce_tmp_1z[3]_i_2__4_n_0 ),
        .O(\r_ce_tmp_1z[4]_i_4__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[4]_i_5 
       (.I0(w_m20[20]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[20]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[20]),
        .O(\r_ce_tmp_1z[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[4]_i_5__0 
       (.I0(w_m21[20]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[20]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[20]),
        .O(\r_ce_tmp_1z[4]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_ce_tmp_1z[4]_i_5__1 
       (.I0(w_m22[20]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[20]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[20]),
        .O(\r_ce_tmp_1z[4]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F8F8F8F8F8F8F88)) 
    \r_cur_adrs[0]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[0]),
        .I2(w_adrs_geo[2]),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[10]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[10]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2_n_6 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[11]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[11]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2_n_5 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[12]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[12]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2_n_4 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[13]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[13]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_7 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[14]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[14]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_6 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[15]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[15]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_5 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[16]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[16]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_4 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[17]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[17]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_7 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[18]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[18]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_6 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[19]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[19]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_5 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[1]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[1]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_7 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[20]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[20]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_4 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[21]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[21]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_7 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[22]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[22]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_6 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[23]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[23]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_5 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[24]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[24]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_4 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[25]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[25]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_7 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[26]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[26]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_6 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[27]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[27]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_5 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[28]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[28]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_4 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[29]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[29]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[29]_i_2_n_7 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[2]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[2]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_6 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[3]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[3]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_5 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[4]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[4]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_4 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[5]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[5]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_7 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[6]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[6]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_6 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[7]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[7]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_5 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[8]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[8]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_4 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8F8F8F8F8F8F888)) 
    \r_cur_adrs[9]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_top_address[9]),
        .I2(\u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2_n_7 ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I5(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\u_geo/u_geo_mem/r_cur_adrs [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_dma_size[15]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[1]),
        .O(r_dma_size));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \r_dma_size[15]_i_2 
       (.I0(s_wb_adr_i[2]),
        .I1(s_wb_stb_i),
        .I2(s_wb_we_i),
        .O(\r_dma_size[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_dma_size[7]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[0]),
        .O(\r_dma_size[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0BF8080)) 
    r_dma_start_i_1
       (.I0(s_wb_dat_i[0]),
        .I1(s_wb_sel_i[0]),
        .I2(r_dma_start_i_2_n_0),
        .I3(\u_sys/w_int_set ),
        .I4(w_dma_start),
        .O(r_dma_start_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    r_dma_start_i_2
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[6]),
        .I2(s_wb_adr_i[2]),
        .I3(s_wb_stb_i),
        .I4(s_wb_we_i),
        .I5(\r_m10[21]_i_2_n_0 ),
        .O(r_dma_start_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \r_dma_top_address[13]_i_1 
       (.I0(s_wb_adr_i[2]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[6]),
        .I4(s_wb_adr_i[5]),
        .I5(s_wb_sel_i[1]),
        .O(r_dma_top_address));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \r_dma_top_address[21]_i_1 
       (.I0(s_wb_adr_i[2]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[6]),
        .I4(s_wb_adr_i[5]),
        .I5(s_wb_sel_i[2]),
        .O(\r_dma_top_address[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \r_dma_top_address[29]_i_1 
       (.I0(s_wb_adr_i[2]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[6]),
        .I4(s_wb_adr_i[5]),
        .I5(s_wb_sel_i[3]),
        .O(\r_dma_top_address[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \r_dma_top_address[29]_i_2 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_stb_i),
        .I2(s_wb_we_i),
        .O(\r_dma_top_address[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \r_dma_top_address[5]_i_1 
       (.I0(s_wb_adr_i[2]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[6]),
        .I4(s_wb_adr_i[5]),
        .I5(s_wb_sel_i[0]),
        .O(\r_dma_top_address[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4444444400400000)) 
    \r_e2[11]_i_1 
       (.I0(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .I1(\u_ras/u_ras_line/r_state_reg_n_0_ ),
        .I2(m_wb_ack_i),
        .I3(\u_mem_arb/w_pri__0 ),
        .I4(\u_ras/u_ras_mem/r_state ),
        .I5(\u_ras/u_ras_line/w_reject__2 ),
        .O(r_e2));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r_e2[11]_i_2 
       (.I0(\u_ras/w_y ),
        .I1(\u_ras/u_ras_line/w_reject1__7 ),
        .I2(\u_ras/w_x ),
        .I3(\u_ras/u_ras_line/w_reject0__7 ),
        .O(\u_ras/u_ras_line/w_reject__2 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBF80)) 
    r_en_cull_i_1
       (.I0(s_wb_dat_i[8]),
        .I1(r_dma_start_i_2_n_0),
        .I2(s_wb_sel_i[1]),
        .I3(w_en_cull),
        .O(r_en_cull_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_err[0]_i_1 
       (.I0(\u_ras/r_err [0]),
        .I1(\u_ras/w_err [0]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(r_err));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4440444444444444)) 
    \r_err[10]_i_1 
       (.I0(\u_ras/u_ras_line/r_state_reg_n_0_ ),
        .I1(\r_err[10]_i_3_n_0 ),
        .I2(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I3(\r_err[10]_i_4_n_0 ),
        .I4(\u_ras/u_ras_line/w_dx ),
        .I5(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_err[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair260" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_err[10]_i_2 
       (.I0(\u_ras/r_err [10]),
        .I1(\u_ras/w_err [10]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_err[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF5FFDDFD)) 
    \r_err[10]_i_3 
       (.I0(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .I1(r_x_reg[1]),
        .I2(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I3(\u_ras/u_ras_line/w_dx ),
        .I4(\u_ras/u_ras_line/r_e2 ),
        .I5(\u_ras/u_ras_line/w_dym__22 ),
        .O(\r_err[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r_err[10]_i_4 
       (.I0(\u_ras/u_ras_line/result0_carry__0_n_2 ),
        .I1(\u_ras/u_ras_line/r_e2 ),
        .O(\r_err[10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair256" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_err[1]_i_1 
       (.I0(\u_ras/r_err [1]),
        .I1(\u_ras/w_err [1]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_err[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair256" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_err[2]_i_1 
       (.I0(\u_ras/r_err [2]),
        .I1(\u_ras/w_err [2]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_err[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair257" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_err[3]_i_1 
       (.I0(\u_ras/r_err [3]),
        .I1(\u_ras/w_err [3]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_err[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair257" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_err[4]_i_1 
       (.I0(\u_ras/r_err [4]),
        .I1(\u_ras/w_err [4]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_err[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair258" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_err[5]_i_1 
       (.I0(\u_ras/r_err [5]),
        .I1(\u_ras/w_err [5]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_err[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair258" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_err[6]_i_1 
       (.I0(\u_ras/r_err [6]),
        .I1(\u_ras/w_err [6]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_err[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair259" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_err[7]_i_1 
       (.I0(\u_ras/r_err [7]),
        .I1(\u_ras/w_err [7]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_err[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair259" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_err[8]_i_1 
       (.I0(\u_ras/r_err [8]),
        .I1(\u_ras/w_err [8]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_err[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair260" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_err[9]_i_1 
       (.I0(\u_ras/r_err [9]),
        .I1(\u_ras/w_err [9]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_err[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[0]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [16]),
        .I1(\r_exp_1z[3]_i_2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m0_out [16]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_exp_l [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0002A0A2080AA8AA)) 
    \r_exp_1z[0]_i_10 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [16]),
        .I1(\r_exp_1z[0]_i_8_n_0 ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I3(\r_exp_1z[0]_i_7_n_0 ),
        .I4(\u_geo/w_vx_clip [16]),
        .I5(\u_geo/w_vy_clip [16]),
        .O(r_exp_1z));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[0]_i_11 
       (.I0(\u_geo/w_vw_mvp [18]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [18]),
        .O(\u_geo/u_geo_clip/w_add_in_a [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0002A0A2080AA8AA)) 
    \r_exp_1z[0]_i_12 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [19]),
        .I1(\r_exp_1z[0]_i_8_n_0 ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I3(\r_exp_1z[3]_i_4__2_n_0 ),
        .I4(\u_geo/w_vx_clip [19]),
        .I5(\u_geo/w_vy_clip [19]),
        .O(\r_exp_1z[0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[0]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [16]),
        .I1(\r_exp_1z[3]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m2_out [16]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_exp_l [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[0]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [16]),
        .I1(\r_exp_1z[3]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add01_out [16]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_exp_l [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAEEFAEAEA220A2A2)) 
    \r_exp_1z[0]_i_1__2 
       (.I0(\r_exp_1z[0]_i_2_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [20]),
        .I2(\r_exp_1z[4]_i_2_n_0 ),
        .I3(\r_exp_1z[0]_i_4_n_0 ),
        .I4(\r_exp_1z[0]_i_5_n_0 ),
        .I5(\u_geo/u_geo_clip/w_add_in_a [16]),
        .O(\u_geo/u_geo_clip/u_fadd/w_exp_l [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFCCAFFF)) 
    \r_exp_1z[0]_i_1__3 
       (.I0(\u_geo/w_vx_pdiv [16]),
        .I1(\u_geo/w_vy_pdiv [16]),
        .I2(\u_geo/w_vx_pdiv [20]),
        .I3(\r_f0[15]_i_2_n_0 ),
        .I4(\u_geo/w_vy_pdiv [20]),
        .O(\u_geo/u_geo_viewport/u_fadd/w_exp_l [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_exp_1z[0]_i_2 
       (.I0(\u_geo/w_vy_clip [16]),
        .I1(\u_geo/w_vx_clip [16]),
        .I2(\r_exp_1z[0]_i_7_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_exp_1z[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[0]_i_3 
       (.I0(\u_geo/w_vw_mvp [20]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [20]),
        .O(\u_geo/u_geo_clip/w_add_in_a [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FE32DC10)) 
    \r_exp_1z[0]_i_4 
       (.I0(\r_exp_1z[0]_i_8_n_0 ),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_exp_1z[3]_i_4__2_n_0 ),
        .I3(\u_geo/w_vx_clip [19]),
        .I4(\u_geo/w_vy_clip [19]),
        .I5(\u_geo/u_geo_clip/w_add_in_a [19]),
        .O(\r_exp_1z[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFB200FFB2)) 
    \r_exp_1z[0]_i_5 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [17]),
        .I1(\r_exp_1z[1]_i_2_n_0 ),
        .I2(r_exp_1z),
        .I3(\u_geo/u_geo_clip/w_add_in_a [18]),
        .I4(\r_exp_1z[2]_i_2_n_0 ),
        .I5(\r_exp_1z[0]_i_12_n_0 ),
        .O(\r_exp_1z[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[0]_i_6 
       (.I0(\u_geo/w_vw_mvp [16]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [16]),
        .O(\u_geo/u_geo_clip/w_add_in_a [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_exp_1z[0]_i_7 
       (.I0(\u_geo/u_geo_clip/r_vz [16]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [16]),
        .O(\r_exp_1z[0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_exp_1z[0]_i_8 
       (.I0(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .O(\r_exp_1z[0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[0]_i_9 
       (.I0(\u_geo/w_vw_mvp [17]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [17]),
        .O(\u_geo/u_geo_clip/w_add_in_a [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[1]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [17]),
        .I1(\r_exp_1z[3]_i_2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m0_out [17]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_exp_l [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[1]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [17]),
        .I1(\r_exp_1z[3]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m2_out [17]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_exp_l [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[1]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [17]),
        .I1(\r_exp_1z[3]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add01_out [17]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_exp_l [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_exp_1z[1]_i_1__2 
       (.I0(\r_exp_1z[1]_i_2_n_0 ),
        .I1(\r_exp_1z[3]_i_3__2_n_0 ),
        .I2(\u_geo/w_vw_mvp [17]),
        .I3(\u_geo/w_state_clip ),
        .I4(\u_geo/w_vw_clip [17]),
        .O(\u_geo/u_geo_clip/u_fadd/w_exp_l [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFCCAFFF)) 
    \r_exp_1z[1]_i_1__3 
       (.I0(\u_geo/w_vx_pdiv [17]),
        .I1(\u_geo/w_vy_pdiv [17]),
        .I2(\u_geo/w_vx_pdiv [20]),
        .I3(\r_f0[15]_i_2_n_0 ),
        .I4(\u_geo/w_vy_pdiv [20]),
        .O(\u_geo/u_geo_viewport/u_fadd/w_exp_l [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_exp_1z[1]_i_2 
       (.I0(\u_geo/w_vy_clip [17]),
        .I1(\u_geo/w_vx_clip [17]),
        .I2(\r_exp_1z[1]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_exp_1z[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_exp_1z[1]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [17]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [17]),
        .O(\r_exp_1z[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[2]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [18]),
        .I1(\r_exp_1z[3]_i_2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m0_out [18]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_exp_l [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[2]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [18]),
        .I1(\r_exp_1z[3]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m2_out [18]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_exp_l [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[2]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [18]),
        .I1(\r_exp_1z[3]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add01_out [18]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_exp_l [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_exp_1z[2]_i_1__2 
       (.I0(\r_exp_1z[2]_i_2_n_0 ),
        .I1(\r_exp_1z[3]_i_3__2_n_0 ),
        .I2(\u_geo/w_vw_mvp [18]),
        .I3(\u_geo/w_state_clip ),
        .I4(\u_geo/w_vw_clip [18]),
        .O(\u_geo/u_geo_clip/u_fadd/w_exp_l [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFCCAFFF)) 
    \r_exp_1z[2]_i_1__3 
       (.I0(\u_geo/w_vx_pdiv [18]),
        .I1(\u_geo/w_vy_pdiv [18]),
        .I2(\u_geo/w_vx_pdiv [20]),
        .I3(\r_f0[15]_i_2_n_0 ),
        .I4(\u_geo/w_vy_pdiv [20]),
        .O(\u_geo/u_geo_viewport/u_fadd/w_exp_l [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_exp_1z[2]_i_2 
       (.I0(\u_geo/w_vy_clip [18]),
        .I1(\u_geo/w_vx_clip [18]),
        .I2(\r_exp_1z[2]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_exp_1z[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_exp_1z[2]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [18]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [18]),
        .O(\r_exp_1z[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[3]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [19]),
        .I1(\r_exp_1z[3]_i_2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m0_out [19]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_exp_l [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[3]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [19]),
        .I1(\r_exp_1z[3]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m2_out [19]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_exp_l [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_exp_1z[3]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [19]),
        .I1(\r_exp_1z[3]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add01_out [19]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_exp_l [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \r_exp_1z[3]_i_1__2 
       (.I0(\r_exp_1z[3]_i_2__2_n_0 ),
        .I1(\r_exp_1z[3]_i_3__2_n_0 ),
        .I2(\u_geo/w_vw_mvp [19]),
        .I3(\u_geo/w_state_clip ),
        .I4(\u_geo/w_vw_clip [19]),
        .O(\u_geo/u_geo_clip/u_fadd/w_exp_l [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAFCCAFFF)) 
    \r_exp_1z[3]_i_1__3 
       (.I0(\u_geo/w_vx_pdiv [19]),
        .I1(\u_geo/w_vy_pdiv [19]),
        .I2(\u_geo/w_vx_pdiv [20]),
        .I3(\r_f0[15]_i_2_n_0 ),
        .I4(\u_geo/w_vy_pdiv [20]),
        .O(\u_geo/u_geo_viewport/u_fadd/w_exp_l [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4D444D444D44DD4D)) 
    \r_exp_1z[3]_i_2 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [20]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [20]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [19]),
        .I3(\u_geo/u_geo_matrix/w_m1_out [19]),
        .I4(\r_exp_1z[3]_i_3_n_0 ),
        .I5(\r_exp_1z[3]_i_4_n_0 ),
        .O(\r_exp_1z[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4D444D444D44DD4D)) 
    \r_exp_1z[3]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [20]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [20]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [19]),
        .I3(\u_geo/u_geo_matrix/w_m3_out [19]),
        .I4(\r_exp_1z[3]_i_3__0_n_0 ),
        .I5(\r_exp_1z[3]_i_4__0_n_0 ),
        .O(\r_exp_1z[3]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4D444D444D44DD4D)) 
    \r_exp_1z[3]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [20]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [20]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [19]),
        .I3(\u_geo/u_geo_matrix/w_add23_out [19]),
        .I4(\r_exp_1z[3]_i_3__1_n_0 ),
        .I5(\r_exp_1z[3]_i_4__1_n_0 ),
        .O(\r_exp_1z[3]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_exp_1z[3]_i_2__2 
       (.I0(\u_geo/w_vy_clip [19]),
        .I1(\u_geo/w_vx_clip [19]),
        .I2(\r_exp_1z[3]_i_4__2_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_exp_1z[3]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F022F0200002F02)) 
    \r_exp_1z[3]_i_3 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [16]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [16]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [17]),
        .I3(\u_geo/u_geo_matrix/w_m0_out [17]),
        .I4(\u_geo/u_geo_matrix/w_m1_out [18]),
        .I5(\u_geo/u_geo_matrix/w_m0_out [18]),
        .O(\r_exp_1z[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F022F0200002F02)) 
    \r_exp_1z[3]_i_3__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [16]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [16]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [17]),
        .I3(\u_geo/u_geo_matrix/w_m2_out [17]),
        .I4(\u_geo/u_geo_matrix/w_m3_out [18]),
        .I5(\u_geo/u_geo_matrix/w_m2_out [18]),
        .O(\r_exp_1z[3]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F022F0200002F02)) 
    \r_exp_1z[3]_i_3__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [16]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [16]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [17]),
        .I3(\u_geo/u_geo_matrix/w_add01_out [17]),
        .I4(\u_geo/u_geo_matrix/w_add23_out [18]),
        .I5(\u_geo/u_geo_matrix/w_add01_out [18]),
        .O(\r_exp_1z[3]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4D444D444D44DD4D)) 
    \r_exp_1z[3]_i_3__2 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [20]),
        .I1(\r_exp_1z[4]_i_2_n_0 ),
        .I2(\u_geo/u_geo_clip/w_add_in_a [19]),
        .I3(\r_exp_1z[3]_i_2__2_n_0 ),
        .I4(\r_exp_1z[3]_i_5_n_0 ),
        .I5(\r_exp_1z[3]_i_6_n_0 ),
        .O(\r_exp_1z[3]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_exp_1z[3]_i_4 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [18]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [18]),
        .O(\r_exp_1z[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_exp_1z[3]_i_4__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [18]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [18]),
        .O(\r_exp_1z[3]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_exp_1z[3]_i_4__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [18]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [18]),
        .O(\r_exp_1z[3]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_exp_1z[3]_i_4__2 
       (.I0(\u_geo/u_geo_clip/r_vz [19]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [19]),
        .O(\r_exp_1z[3]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002F02)) 
    \r_exp_1z[3]_i_5 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [16]),
        .I1(\r_exp_1z[0]_i_2_n_0 ),
        .I2(\r_exp_1z[1]_i_2_n_0 ),
        .I3(\u_geo/u_geo_clip/w_add_in_a [17]),
        .I4(\r_exp_1z[3]_i_7_n_0 ),
        .O(\r_exp_1z[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \r_exp_1z[3]_i_6 
       (.I0(\u_geo/w_vw_clip [18]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_mvp [18]),
        .I3(\r_exp_1z[2]_i_2_n_0 ),
        .O(\r_exp_1z[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FE32DC10)) 
    \r_exp_1z[3]_i_7 
       (.I0(\r_exp_1z[0]_i_8_n_0 ),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I2(\r_exp_1z[2]_i_3_n_0 ),
        .I3(\u_geo/w_vx_clip [18]),
        .I4(\u_geo/w_vy_clip [18]),
        .I5(\u_geo/u_geo_clip/w_add_in_a [18]),
        .O(\r_exp_1z[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_exp_1z[4]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [20]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [20]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_exp_l [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_exp_1z[4]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [20]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [20]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_exp_l [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_exp_1z[4]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [20]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [20]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_exp_l [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFE2)) 
    \r_exp_1z[4]_i_1__2 
       (.I0(\u_geo/w_vw_clip [20]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_mvp [20]),
        .I3(\r_exp_1z[4]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/u_fadd/w_exp_l [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_exp_1z[4]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [20]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [20]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_exp_1z[4]_i_2 
       (.I0(\u_geo/w_vy_clip [20]),
        .I1(\u_geo/w_vx_clip [20]),
        .I2(\r_exp_1z[4]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_exp_1z[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_exp_1z[4]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [20]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [20]),
        .O(\r_exp_1z[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair269" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[0]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [0]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [0]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[0]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [0]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [0]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[0]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [0]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [0]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[0]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [0]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [0]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(r_f0),
        .O(\u_geo/u_geo_clip/w_f0 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[0]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [0]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [0]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[0]_i_2 
       (.I0(\u_geo/w_vy_clip [0]),
        .I1(\u_geo/w_vx_clip [0]),
        .I2(\r_f0[0]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(r_f0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[0]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [0]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [0]),
        .O(\r_f0[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[10]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [10]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [10]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair247" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[10]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [10]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [10]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[10]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [10]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [10]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[10]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [10]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [10]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[10]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[10]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [10]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [10]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[10]_i_2 
       (.I0(\u_geo/w_vy_clip [10]),
        .I1(\u_geo/w_vx_clip [10]),
        .I2(\r_f0[10]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[10]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [10]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [10]),
        .O(\r_f0[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[11]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [11]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [11]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair246" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[11]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [11]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [11]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[11]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [11]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [11]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[11]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [11]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [11]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[11]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[11]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [11]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [11]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[11]_i_2 
       (.I0(\u_geo/w_vy_clip [11]),
        .I1(\u_geo/w_vx_clip [11]),
        .I2(\r_f0[11]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[11]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [11]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [11]),
        .O(\r_f0[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[12]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [12]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [12]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair245" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[12]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [12]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [12]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[12]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [12]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [12]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[12]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [12]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [12]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[12]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[12]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [12]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [12]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[12]_i_2 
       (.I0(\u_geo/w_vy_clip [12]),
        .I1(\u_geo/w_vx_clip [12]),
        .I2(\r_f0[12]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[12]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [12]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [12]),
        .O(\r_f0[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[13]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [13]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [13]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair244" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[13]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [13]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [13]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[13]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [13]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [13]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[13]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [13]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [13]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[13]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[13]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [13]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [13]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[13]_i_2 
       (.I0(\u_geo/w_vy_clip [13]),
        .I1(\u_geo/w_vx_clip [13]),
        .I2(\r_f0[13]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[13]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [13]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [13]),
        .O(\r_f0[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[14]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [14]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [14]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010000)) 
    \r_f0[14]_i_10 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [11]),
        .I1(\u_geo/u_geo_viewport/w_fadd_a [12]),
        .I2(\u_geo/u_geo_viewport/w_fadd_a [13]),
        .I3(\u_geo/u_geo_viewport/w_fadd_a [14]),
        .I4(\r_f0[14]_i_14_n_0 ),
        .O(\r_f0[14]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000110C1D)) 
    \r_f0[14]_i_11 
       (.I0(\u_geo/w_vy_pdiv [2]),
        .I1(\r_f0[15]_i_2_n_0 ),
        .I2(\u_geo/w_vx_pdiv [2]),
        .I3(\u_geo/w_vy_pdiv [1]),
        .I4(\u_geo/w_vx_pdiv [1]),
        .I5(\u_geo/u_geo_viewport/w_fadd_a [0]),
        .O(\r_f0[14]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000151)) 
    \r_f0[14]_i_12 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [6]),
        .I1(\u_geo/w_vy_pdiv [5]),
        .I2(\r_f0[15]_i_2_n_0 ),
        .I3(\u_geo/w_vx_pdiv [5]),
        .I4(\u_geo/u_geo_viewport/w_fadd_a [4]),
        .I5(\u_geo/u_geo_viewport/w_fadd_a [3]),
        .O(\r_f0[14]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \r_f0[14]_i_13 
       (.I0(\u_geo/u_geo_viewport/sel0 [1]),
        .I1(\u_geo/u_geo_viewport/sel0 [0]),
        .I2(\u_geo/u_geo_viewport/sel0 [2]),
        .O(\r_f0[14]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000101010001)) 
    \r_f0[14]_i_14 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [10]),
        .I1(\u_geo/u_geo_viewport/w_fadd_a [9]),
        .I2(\u_geo/u_geo_viewport/w_fadd_a [8]),
        .I3(\u_geo/w_vy_pdiv [7]),
        .I4(\r_f0[15]_i_2_n_0 ),
        .I5(\u_geo/w_vx_pdiv [7]),
        .O(\r_f0[14]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair243" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[14]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [14]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [14]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[14]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [14]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [14]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[14]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [14]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [14]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[14]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3333333733333332)) 
    \r_f0[14]_i_1__3 
       (.I0(\u_geo/u_geo_viewport/sel0 [4]),
        .I1(\u_geo/u_geo_viewport/w_fadd_a [20]),
        .I2(\u_geo/u_geo_viewport/sel0 [3]),
        .I3(\u_geo/u_geo_viewport/sel0 [2]),
        .I4(\u_geo/u_geo_viewport/sel0 [1]),
        .I5(\r_f0[14]_i_7_n_0 ),
        .O(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[14]_i_2 
       (.I0(\u_geo/w_vy_clip [14]),
        .I1(\u_geo/w_vx_clip [14]),
        .I2(\r_f0[14]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[14]_i_2__0 
       (.I0(\u_geo/w_vy_pdiv [14]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [14]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[14]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [14]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [14]),
        .O(\r_f0[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC00CA0A0C00C0A0A)) 
    \r_f0[14]_i_3__0 
       (.I0(\u_geo/w_vy_pdiv [19]),
        .I1(\u_geo/w_vx_pdiv [19]),
        .I2(\r_f0[14]_i_8_n_0 ),
        .I3(\u_geo/w_vx_pdiv [20]),
        .I4(\r_f0[15]_i_2_n_0 ),
        .I5(\u_geo/w_vy_pdiv [20]),
        .O(\u_geo/u_geo_viewport/sel0 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h665A)) 
    \r_f0[14]_i_4 
       (.I0(\r_f0[14]_i_8_n_0 ),
        .I1(\u_geo/w_vx_pdiv [19]),
        .I2(\u_geo/w_vy_pdiv [19]),
        .I3(\r_f0[15]_i_2_n_0 ),
        .O(\u_geo/u_geo_viewport/sel0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h665A)) 
    \r_f0[14]_i_5 
       (.I0(\r_f0[14]_i_9_n_0 ),
        .I1(\u_geo/w_vx_pdiv [18]),
        .I2(\u_geo/w_vy_pdiv [18]),
        .I3(\r_f0[15]_i_2_n_0 ),
        .O(\u_geo/u_geo_viewport/sel0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5A335ACC0F000FFF)) 
    \r_f0[14]_i_6 
       (.I0(\u_geo/w_vx_pdiv [16]),
        .I1(\u_geo/w_vy_pdiv [16]),
        .I2(\u_geo/w_vx_pdiv [17]),
        .I3(\r_f0[15]_i_2_n_0 ),
        .I4(\u_geo/w_vy_pdiv [17]),
        .I5(\u_geo/u_geo_viewport/w_fadd_a [20]),
        .O(\u_geo/u_geo_viewport/sel0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FFFFD555D555)) 
    \r_f0[14]_i_7 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [15]),
        .I1(\r_f0[14]_i_10_n_0 ),
        .I2(\r_f0[14]_i_11_n_0 ),
        .I3(\r_f0[14]_i_12_n_0 ),
        .I4(\u_geo/u_geo_viewport/w_fadd_a [20]),
        .I5(\r_f0[14]_i_13_n_0 ),
        .O(\r_f0[14]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBA0A088BBAFAF)) 
    \r_f0[14]_i_8 
       (.I0(\r_f0[14]_i_9_n_0 ),
        .I1(\u_geo/w_vx_pdiv [18]),
        .I2(\u_geo/w_vy_pdiv [18]),
        .I3(\u_geo/w_vx_pdiv [20]),
        .I4(\r_f0[15]_i_2_n_0 ),
        .I5(\u_geo/w_vy_pdiv [20]),
        .O(\r_f0[14]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0CCA000FFFFFFFF)) 
    \r_f0[14]_i_9 
       (.I0(\u_geo/w_vx_pdiv [16]),
        .I1(\u_geo/w_vy_pdiv [16]),
        .I2(\u_geo/w_vx_pdiv [17]),
        .I3(\r_f0[15]_i_2_n_0 ),
        .I4(\u_geo/w_vy_pdiv [17]),
        .I5(\u_geo/u_geo_viewport/w_fadd_a [20]),
        .O(\r_f0[14]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[15]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [15]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [15]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF7788FFFF7588FF)) 
    \r_f0[15]_i_10 
       (.I0(\r_f0[15]_i_15_n_0 ),
        .I1(\r_f0[15]_i_16_n_0 ),
        .I2(\r_exp_1z[3]_i_5_n_0 ),
        .I3(\u_geo/u_geo_clip/w_add_in_a [18]),
        .I4(\r_exp_1z[2]_i_2_n_0 ),
        .I5(\r_exp_1z[0]_i_12_n_0 ),
        .O(\r_f0[15]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9A95)) 
    \r_f0[15]_i_11 
       (.I0(\r_exp_1z[2]_i_2_n_0 ),
        .I1(\u_geo/w_vw_mvp [18]),
        .I2(\u_geo/w_state_clip ),
        .I3(\u_geo/w_vw_clip [18]),
        .O(\r_f0[15]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEAEE7F77FFFFFFFF)) 
    \r_f0[15]_i_12 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [16]),
        .I1(\r_f0[15]_i_15_n_0 ),
        .I2(\r_f0[15]_i_16_n_0 ),
        .I3(\r_exp_1z[0]_i_5_n_0 ),
        .I4(\r_exp_1z[0]_i_2_n_0 ),
        .I5(\r_f1t[15]_i_7__2_n_0 ),
        .O(\r_f0[15]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000D4DD2B220000)) 
    \r_f0[15]_i_13 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [20]),
        .I1(\r_exp_1z[4]_i_2_n_0 ),
        .I2(\r_exp_1z[0]_i_4_n_0 ),
        .I3(\r_exp_1z[0]_i_5_n_0 ),
        .I4(\r_exp_1z[1]_i_2_n_0 ),
        .I5(\u_geo/u_geo_clip/w_add_in_a [17]),
        .O(\r_f0[15]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0240)) 
    \r_f0[15]_i_14 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [20]),
        .I1(\r_exp_1z[4]_i_2_n_0 ),
        .I2(\u_geo/u_geo_clip/w_add_in_a [19]),
        .I3(\r_exp_1z[3]_i_2__2_n_0 ),
        .O(\r_f0[15]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f0[15]_i_15 
       (.I0(\r_exp_1z[4]_i_2_n_0 ),
        .I1(\u_geo/w_vw_clip [20]),
        .I2(\u_geo/w_state_clip ),
        .I3(\u_geo/w_vw_mvp [20]),
        .O(\r_f0[15]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \r_f0[15]_i_16 
       (.I0(\u_geo/w_vw_mvp [20]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [20]),
        .I3(\r_exp_1z[4]_i_2_n_0 ),
        .I4(\r_exp_1z[0]_i_4_n_0 ),
        .O(\r_f0[15]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[15]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [15]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [15]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[15]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [15]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [15]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[15]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [15]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/u_geo_clip/r_vw_reg_n_0_ ),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[15]_i_3__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFB8)) 
    \r_f0[15]_i_1__3 
       (.I0(\u_geo/w_vx_pdiv [15]),
        .I1(\r_f0[15]_i_2_n_0 ),
        .I2(\u_geo/w_vy_pdiv [15]),
        .I3(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ),
        .O(\u_geo/u_geo_viewport/w_f0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \r_f0[15]_i_2 
       (.I0(\u_geo/u_geo_viewport/r_state [2]),
        .I1(\u_geo/u_geo_viewport/r_state [3]),
        .I2(\u_geo/u_geo_viewport/r_state [1]),
        .I3(\u_geo/u_geo_viewport/r_state [0]),
        .O(\r_f0[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000400FFFFFFFF)) 
    \r_f0[15]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/data0 ),
        .I1(\r_f1t[15]_i_6_n_0 ),
        .I2(\r_f1t[15]_i_4_n_0 ),
        .I3(\r_f1t[15]_i_5__0_n_0 ),
        .I4(\r_f0[15]_i_3_n_0 ),
        .I5(\r_exp_1z[3]_i_2_n_0 ),
        .O(\r_f0[15]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000400FFFFFFFF)) 
    \r_f0[15]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/data0 ),
        .I1(\r_f1t[15]_i_6__0_n_0 ),
        .I2(\r_f1t[15]_i_4__0_n_0 ),
        .I3(\r_f1t[15]_i_5__1_n_0 ),
        .I4(\r_f0[15]_i_3__0_n_0 ),
        .I5(\r_exp_1z[3]_i_2__0_n_0 ),
        .O(\r_f0[15]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000400FFFFFFFF)) 
    \r_f0[15]_i_2__2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/data0 ),
        .I1(\r_f1t[15]_i_6__1_n_0 ),
        .I2(\r_f1t[15]_i_4__1_n_0 ),
        .I3(\r_f1t[15]_i_5__2_n_0 ),
        .I4(\r_f0[15]_i_3__1_n_0 ),
        .I5(\r_exp_1z[3]_i_2__1_n_0 ),
        .O(\r_f0[15]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000054FFFFFFFF)) 
    \r_f0[15]_i_2__3 
       (.I0(\u_geo/u_geo_clip/data0 ),
        .I1(\r_f0[15]_i_4_n_0 ),
        .I2(\r_f0[15]_i_5_n_0 ),
        .I3(\r_f0[15]_i_6_n_0 ),
        .I4(\r_f0[15]_i_7_n_0 ),
        .I5(\r_exp_1z[3]_i_3__2_n_0 ),
        .O(\r_f0[15]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_f0[15]_i_3 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\r_f1t[11]_i_5_n_0 ),
        .O(\r_f0[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_f0[15]_i_3__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\r_f1t[11]_i_5__0_n_0 ),
        .O(\r_f0[15]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_f0[15]_i_3__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\r_f1t[11]_i_5__1_n_0 ),
        .O(\r_f0[15]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[15]_i_3__2 
       (.I0(\u_geo/w_vy_clip [15]),
        .I1(\u_geo/w_vx_clip [15]),
        .I2(\r_f0[15]_i_8_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[15]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF88880888)) 
    \r_f0[15]_i_4 
       (.I0(\r_f0[15]_i_9_n_0 ),
        .I1(\r_f0[15]_i_10_n_0 ),
        .I2(\r_f0[15]_i_11_n_0 ),
        .I3(\r_f0[15]_i_12_n_0 ),
        .I4(\r_f0[15]_i_13_n_0 ),
        .I5(\r_f0[15]_i_14_n_0 ),
        .O(\r_f0[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB847)) 
    \r_f0[15]_i_5 
       (.I0(\u_geo/w_vw_mvp [20]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [20]),
        .I3(\r_exp_1z[4]_i_2_n_0 ),
        .O(\r_f0[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF3F99F966F6FF3F)) 
    \r_f0[15]_i_6 
       (.I0(\r_exp_1z[3]_i_3__2_n_0 ),
        .I1(\r_f0[15]_i_9_n_0 ),
        .I2(\r_f0[15]_i_12_n_0 ),
        .I3(\r_f0[15]_i_13_n_0 ),
        .I4(\r_exp_1z[2]_i_2_n_0 ),
        .I5(\u_geo/u_geo_clip/w_add_in_a [18]),
        .O(\r_f0[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7D777DDD)) 
    \r_f0[15]_i_7 
       (.I0(\r_f1t[15]_i_7__2_n_0 ),
        .I1(\r_exp_1z[0]_i_2_n_0 ),
        .I2(\u_geo/w_vw_mvp [16]),
        .I3(\u_geo/w_state_clip ),
        .I4(\u_geo/w_vw_clip [16]),
        .O(\r_f0[15]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[15]_i_8 
       (.I0(\u_geo/u_geo_clip/r_vz [15]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [15]),
        .O(\r_f0[15]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB847)) 
    \r_f0[15]_i_9 
       (.I0(\u_geo/w_vw_mvp [19]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [19]),
        .I3(\r_exp_1z[3]_i_2__2_n_0 ),
        .O(\r_f0[15]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair270" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[1]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [1]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [1]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[1]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [1]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [1]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[1]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [1]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [1]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[1]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [1]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [1]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[1]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[1]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [1]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [1]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[1]_i_2 
       (.I0(\u_geo/w_vy_clip [1]),
        .I1(\u_geo/w_vx_clip [1]),
        .I2(\r_f0[1]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[1]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [1]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [1]),
        .O(\r_f0[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair271" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[2]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [2]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [2]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair243" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[2]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [2]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [2]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[2]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [2]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [2]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[2]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [2]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [2]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[2]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[2]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [2]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [2]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[2]_i_2 
       (.I0(\u_geo/w_vy_clip [2]),
        .I1(\u_geo/w_vx_clip [2]),
        .I2(\r_f0[2]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[2]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [2]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [2]),
        .O(\r_f0[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair272" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[3]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [3]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [3]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair244" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[3]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [3]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [3]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[3]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [3]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [3]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[3]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [3]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [3]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[3]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[3]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [3]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [3]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[3]_i_2 
       (.I0(\u_geo/w_vy_clip [3]),
        .I1(\u_geo/w_vx_clip [3]),
        .I2(\r_f0[3]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[3]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [3]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [3]),
        .O(\r_f0[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[4]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [4]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [4]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair245" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[4]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [4]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [4]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[4]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [4]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [4]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[4]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [4]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [4]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[4]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[4]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [4]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [4]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[4]_i_2 
       (.I0(\u_geo/w_vy_clip [4]),
        .I1(\u_geo/w_vx_clip [4]),
        .I2(\r_f0[4]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[4]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [4]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [4]),
        .O(\r_f0[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair272" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[5]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [5]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [5]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair246" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[5]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [5]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [5]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[5]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [5]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [5]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[5]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [5]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [5]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[5]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[5]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [5]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [5]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[5]_i_2 
       (.I0(\u_geo/w_vy_clip [5]),
        .I1(\u_geo/w_vx_clip [5]),
        .I2(\r_f0[5]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[5]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [5]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [5]),
        .O(\r_f0[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair271" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[6]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [6]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [6]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair247" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[6]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [6]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [6]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[6]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [6]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [6]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[6]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [6]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [6]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[6]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[6]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [6]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [6]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[6]_i_2 
       (.I0(\u_geo/w_vy_clip [6]),
        .I1(\u_geo/w_vx_clip [6]),
        .I2(\r_f0[6]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[6]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [6]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [6]),
        .O(\r_f0[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair270" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[7]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [7]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [7]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair248" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[7]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [7]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [7]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[7]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [7]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [7]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[7]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [7]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [7]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[7]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[7]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [7]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [7]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[7]_i_2 
       (.I0(\u_geo/w_vy_clip [7]),
        .I1(\u_geo/w_vx_clip [7]),
        .I2(\r_f0[7]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[7]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [7]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [7]),
        .O(\r_f0[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair269" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[8]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [8]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [8]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[8]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [8]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [8]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[8]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [8]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [8]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[8]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [8]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [8]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[8]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[8]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [8]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [8]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[8]_i_2 
       (.I0(\u_geo/w_vy_clip [8]),
        .I1(\u_geo/w_vx_clip [8]),
        .I2(\r_f0[8]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[8]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [8]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [8]),
        .O(\r_f0[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[9]_i_1 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [9]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [9]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair248" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[9]_i_1__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [9]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [9]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f0[9]_i_1__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [9]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [9]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \r_f0[9]_i_1__2 
       (.I0(\u_geo/w_vw_mvp [9]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [9]),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f0[9]_i_2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f0 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f0[9]_i_1__3 
       (.I0(\u_geo/w_vy_pdiv [9]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [9]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    \r_f0[9]_i_2 
       (.I0(\u_geo/w_vy_clip [9]),
        .I1(\u_geo/w_vx_clip [9]),
        .I2(\r_f0[9]_i_3_n_0 ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(\r_f0[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \r_f0[9]_i_3 
       (.I0(\u_geo/u_geo_clip/r_vz [9]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [9]),
        .O(\r_f0[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[0]_i_1 
       (.I0(\r_f1t[1]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[0]_i_2_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[0]_i_3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[0]_i_1__0 
       (.I0(\r_f1t[1]_i_2__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(r_f1t),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[0]_i_3__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[0]_i_1__1 
       (.I0(\r_f1t[1]_i_2__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[0]_i_2__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[0]_i_3__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[0]_i_1__2 
       (.I0(\r_f1t[1]_i_2__2_n_0 ),
        .I1(\r_f1t[15]_i_6__2_n_0 ),
        .I2(\r_f1t[0]_i_2__2_n_0 ),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f1t[15]_i_5_n_0 ),
        .I5(\r_f1t[0]_i_3__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF544454445444)) 
    \r_f1t[0]_i_1__3 
       (.I0(\r_f1t[13]_i_4__2_n_0 ),
        .I1(\r_f1t[0]_i_2__3_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[1]_i_2__3_n_0 ),
        .I4(\r_f1t[12]_i_2__3_n_0 ),
        .I5(\r_f1t[3]_i_2__3_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[0]_i_2 
       (.I0(\r_f1t[2]_i_4__0_n_0 ),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[0]_i_4__1_n_0 ),
        .O(\r_f1t[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[0]_i_2__0 
       (.I0(\r_f1t[2]_i_4__1_n_0 ),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[0]_i_4__2_n_0 ),
        .O(r_f1t));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[0]_i_2__1 
       (.I0(\r_f1t[2]_i_4__2_n_0 ),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[0]_i_4__3_n_0 ),
        .O(\r_f1t[0]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[0]_i_2__2 
       (.I0(\r_f1t[2]_i_4_n_0 ),
        .I1(\r_f1t[15]_i_2_n_0 ),
        .I2(\r_f1t[0]_i_4_n_0 ),
        .O(\r_f1t[0]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000AAAAFCCC)) 
    \r_f1t[0]_i_2__3 
       (.I0(\r_f1t[2]_i_3__3_n_0 ),
        .I1(\r_f1t[0]_i_3__3_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [2]),
        .I3(\r_f1t[0]_i_4__0_n_0 ),
        .I4(\u_geo/u_geo_viewport/sel0 [1]),
        .I5(\u_geo/u_geo_viewport/sel0 [0]),
        .O(\r_f1t[0]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[0]_i_3 
       (.I0(\r_f1t[2]_i_6_n_0 ),
        .I1(\r_f1t[0]_i_5__0_n_0 ),
        .I2(\r_f1t[15]_i_5__0_n_0 ),
        .I3(\r_f1t[3]_i_5__0_n_0 ),
        .I4(\r_f1t[15]_i_4_n_0 ),
        .I5(\r_f1t[1]_i_5__0_n_0 ),
        .O(\r_f1t[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[0]_i_3__0 
       (.I0(\r_f1t[2]_i_6__0_n_0 ),
        .I1(\r_f1t[0]_i_5__1_n_0 ),
        .I2(\r_f1t[15]_i_5__1_n_0 ),
        .I3(\r_f1t[3]_i_5__1_n_0 ),
        .I4(\r_f1t[15]_i_4__0_n_0 ),
        .I5(\r_f1t[1]_i_5__1_n_0 ),
        .O(\r_f1t[0]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[0]_i_3__1 
       (.I0(\r_f1t[2]_i_6__1_n_0 ),
        .I1(\r_f1t[0]_i_5__2_n_0 ),
        .I2(\r_f1t[15]_i_5__2_n_0 ),
        .I3(\r_f1t[3]_i_5__2_n_0 ),
        .I4(\r_f1t[15]_i_4__1_n_0 ),
        .I5(\r_f1t[1]_i_5__2_n_0 ),
        .O(\r_f1t[0]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[0]_i_3__2 
       (.I0(\r_f1t[2]_i_5__2_n_0 ),
        .I1(\r_f1t[0]_i_5_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[3]_i_5_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[1]_i_5_n_0 ),
        .O(\r_f1t[0]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000AAAAFC0C)) 
    \r_f1t[0]_i_3__3 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [8]),
        .I1(\u_geo/w_vy_pdiv [0]),
        .I2(\r_f0[15]_i_2_n_0 ),
        .I3(\u_geo/w_vx_pdiv [0]),
        .I4(\u_geo/u_geo_viewport/sel0 [3]),
        .I5(\u_geo/u_geo_viewport/sel0 [2]),
        .O(\r_f1t[0]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3030505F3F3F505F)) 
    \r_f1t[0]_i_4 
       (.I0(\r_f0[4]_i_2_n_0 ),
        .I1(\r_f0[12]_i_2_n_0 ),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(r_f0),
        .I4(\r_f1t[15]_i_9_n_0 ),
        .I5(\r_f0[8]_i_2_n_0 ),
        .O(\r_f1t[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFAFA0C0C0AFA0)) 
    \r_f1t[0]_i_4__0 
       (.I0(\u_geo/w_vy_pdiv [12]),
        .I1(\u_geo/w_vx_pdiv [12]),
        .I2(\u_geo/u_geo_viewport/sel0 [3]),
        .I3(\u_geo/w_vy_pdiv [4]),
        .I4(\r_f0[15]_i_2_n_0 ),
        .I5(\u_geo/w_vx_pdiv [4]),
        .O(\r_f1t[0]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[0]_i_4__1 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [4]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [12]),
        .I3(\r_f1t[11]_i_5_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m1_out [0]),
        .I5(\u_geo/u_geo_matrix/w_m1_out [8]),
        .O(\r_f1t[0]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[0]_i_4__2 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [4]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [12]),
        .I3(\r_f1t[11]_i_5__0_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m3_out [0]),
        .I5(\u_geo/u_geo_matrix/w_m3_out [8]),
        .O(\r_f1t[0]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[0]_i_4__3 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [4]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [12]),
        .I3(\r_f1t[11]_i_5__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add23_out [0]),
        .I5(\u_geo/u_geo_matrix/w_add23_out [8]),
        .O(\r_f1t[0]_i_4__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3030505F3F3F505F)) 
    \r_f1t[0]_i_5 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [4]),
        .I1(\u_geo/u_geo_clip/w_add_in_a [12]),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\u_geo/u_geo_clip/w_add_in_a [0]),
        .I4(\r_f1t[15]_i_9_n_0 ),
        .I5(\u_geo/u_geo_clip/w_add_in_a [8]),
        .O(\r_f1t[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[0]_i_5__0 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [4]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [12]),
        .I3(\r_f1t[11]_i_5_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m0_out [0]),
        .I5(\u_geo/u_geo_matrix/w_m0_out [8]),
        .O(\r_f1t[0]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[0]_i_5__1 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [4]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [12]),
        .I3(\r_f1t[11]_i_5__0_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m2_out [0]),
        .I5(\u_geo/u_geo_matrix/w_m2_out [8]),
        .O(\r_f1t[0]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[0]_i_5__2 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [4]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [12]),
        .I3(\r_f1t[11]_i_5__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add01_out [0]),
        .I5(\u_geo/u_geo_matrix/w_add01_out [8]),
        .O(\r_f1t[0]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[10]_i_1 
       (.I0(\r_f1t[11]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[10]_i_2_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[10]_i_3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[10]_i_1__0 
       (.I0(\r_f1t[11]_i_2__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\r_f1t[10]_i_2__0_n_0 ),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[10]_i_3__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[10]_i_1__1 
       (.I0(\r_f1t[11]_i_2__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[10]_i_2__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[10]_i_3__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h303F000055550000)) 
    \r_f1t[10]_i_1__2 
       (.I0(\r_f1t[11]_i_2__2_n_0 ),
        .I1(\r_f1t[10]_i_2__2_n_0 ),
        .I2(\r_f0[15]_i_2__3_n_0 ),
        .I3(\r_f1t[10]_i_3__2_n_0 ),
        .I4(\r_f1t[15]_i_5_n_0 ),
        .I5(\r_f1t[15]_i_6__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[10]_i_1__3 
       (.I0(\r_f1t[14]_i_2__3_n_0 ),
        .I1(\r_f1t[11]_i_3__2_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[11]_i_4__0_n_0 ),
        .I4(\r_f1t[10]_i_2__3_n_0 ),
        .I5(\r_f1t[13]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[10]_i_2 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [12]),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[11]_i_4__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m1_out [10]),
        .I4(\r_f1t[11]_i_5_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m1_out [14]),
        .O(\r_f1t[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[10]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [12]),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[11]_i_4__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m3_out [10]),
        .I4(\r_f1t[11]_i_5__0_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m3_out [14]),
        .O(\r_f1t[10]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[10]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [12]),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[11]_i_4__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add23_out [10]),
        .I4(\r_f1t[11]_i_5__1_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_add23_out [14]),
        .O(\r_f1t[10]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[10]_i_2__2 
       (.I0(\r_f0[12]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_2_n_0 ),
        .I2(\r_f1t[15]_i_9_n_0 ),
        .I3(\r_f0[10]_i_2_n_0 ),
        .I4(\r_f1t[15]_i_8__2_n_0 ),
        .I5(\r_f0[14]_i_2_n_0 ),
        .O(\r_f1t[10]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB88830003000)) 
    \r_f1t[10]_i_2__3 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [12]),
        .I1(\u_geo/u_geo_viewport/sel0 [1]),
        .I2(\u_geo/u_geo_viewport/w_fadd_a [14]),
        .I3(\r_f1t[11]_i_5__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/w_fadd_a [10]),
        .I5(\r_f1t[15]_i_4__2_n_0 ),
        .O(\r_f1t[10]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \r_f1t[10]_i_3 
       (.I0(\r_f1t[10]_i_4_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [16]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [16]),
        .I3(\r_f1t[11]_i_6_n_0 ),
        .O(\r_f1t[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \r_f1t[10]_i_3__0 
       (.I0(\r_f1t[10]_i_4__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [16]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [16]),
        .I3(\r_f1t[11]_i_6__0_n_0 ),
        .O(\r_f1t[10]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \r_f1t[10]_i_3__1 
       (.I0(\r_f1t[10]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [16]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [16]),
        .I3(\r_f1t[11]_i_6__1_n_0 ),
        .O(\r_f1t[10]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[10]_i_3__2 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [12]),
        .I1(\r_f1t[15]_i_2_n_0 ),
        .I2(\r_f1t[15]_i_9_n_0 ),
        .I3(\u_geo/u_geo_clip/w_add_in_a [10]),
        .I4(\r_f1t[15]_i_8__2_n_0 ),
        .I5(\u_geo/u_geo_clip/w_add_in_a [14]),
        .O(\r_f1t[10]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[10]_i_4 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [12]),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[11]_i_4__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [10]),
        .I4(\r_f1t[11]_i_5_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m0_out [14]),
        .O(\r_f1t[10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[10]_i_4__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [12]),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[11]_i_4__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [10]),
        .I4(\r_f1t[11]_i_5__0_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m2_out [14]),
        .O(\r_f1t[10]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[10]_i_4__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [12]),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[11]_i_4__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [10]),
        .I4(\r_f1t[11]_i_5__1_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_add01_out [14]),
        .O(\r_f1t[10]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[11]_i_1 
       (.I0(\r_f1t[12]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[11]_i_2_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[11]_i_3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[11]_i_1__0 
       (.I0(\r_f1t[12]_i_2__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\r_f1t[11]_i_2__0_n_0 ),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[11]_i_3__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[11]_i_1__1 
       (.I0(\r_f1t[12]_i_2__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[11]_i_2__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[11]_i_3__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5030)) 
    \r_f1t[11]_i_1__2 
       (.I0(\r_f1t[11]_i_2__2_n_0 ),
        .I1(\r_f1t[12]_i_3__2_n_0 ),
        .I2(\r_f1t[15]_i_5_n_0 ),
        .I3(\r_f1t[15]_i_6__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[11]_i_1__3 
       (.I0(\r_f1t[11]_i_2__3_n_0 ),
        .I1(\r_f1t[11]_i_3__2_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[12]_i_4__2_n_0 ),
        .I4(\r_f1t[11]_i_4__0_n_0 ),
        .I5(\r_f1t[13]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[11]_i_2 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [13]),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[11]_i_4__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m1_out [11]),
        .I4(\r_f1t[11]_i_5_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m1_out [15]),
        .O(\r_f1t[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[11]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [13]),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[11]_i_4__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m3_out [11]),
        .I4(\r_f1t[11]_i_5__0_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m3_out [15]),
        .O(\r_f1t[11]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[11]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [13]),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[11]_i_4__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add23_out [11]),
        .I4(\r_f1t[11]_i_5__1_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_add23_out [15]),
        .O(\r_f1t[11]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[11]_i_2__2 
       (.I0(\r_f1t[11]_i_3__3_n_0 ),
        .I1(\r_f1t[11]_i_4_n_0 ),
        .I2(\r_f0[15]_i_2__3_n_0 ),
        .I3(\r_f1t[11]_i_5__3_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[11]_i_6__2_n_0 ),
        .O(\r_f1t[11]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \r_f1t[11]_i_2__3 
       (.I0(\u_geo/u_geo_viewport/sel0 [0]),
        .I1(\u_geo/u_geo_viewport/sel0 [1]),
        .I2(\u_geo/u_geo_viewport/sel0 [4]),
        .O(\r_f1t[11]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBB8B88BBBB8BBB)) 
    \r_f1t[11]_i_3 
       (.I0(\r_f1t[11]_i_6_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m0_out [14]),
        .I3(\r_f1t[15]_i_4_n_0 ),
        .I4(\r_f0[15]_i_3_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m0_out [12]),
        .O(\r_f1t[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBB8B88BBBB8BBB)) 
    \r_f1t[11]_i_3__0 
       (.I0(\r_f1t[11]_i_6__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m2_out [14]),
        .I3(\r_f1t[15]_i_4__0_n_0 ),
        .I4(\r_f0[15]_i_3__0_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m2_out [12]),
        .O(\r_f1t[11]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBB8B88BBBB8BBB)) 
    \r_f1t[11]_i_3__1 
       (.I0(\r_f1t[11]_i_6__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add01_out [14]),
        .I3(\r_f1t[15]_i_4__1_n_0 ),
        .I4(\r_f0[15]_i_3__1_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_add01_out [12]),
        .O(\r_f1t[11]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_f1t[11]_i_3__2 
       (.I0(\r_f1t[11]_i_5__2_n_0 ),
        .I1(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ),
        .O(\r_f1t[11]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \r_f1t[11]_i_3__3 
       (.I0(\r_f1t[15]_i_8__2_n_0 ),
        .I1(\r_f1t[15]_i_9_n_0 ),
        .I2(\r_f0[13]_i_2_n_0 ),
        .O(\r_f1t[11]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[11]_i_4 
       (.I0(\r_f1t[15]_i_9_n_0 ),
        .I1(\r_f0[11]_i_2_n_0 ),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\r_f0[15]_i_3__2_n_0 ),
        .O(\r_f1t[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBB88830003000)) 
    \r_f1t[11]_i_4__0 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [13]),
        .I1(\u_geo/u_geo_viewport/sel0 [1]),
        .I2(\u_geo/u_geo_viewport/w_fadd_a [15]),
        .I3(\r_f1t[11]_i_5__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/w_fadd_a [11]),
        .I5(\r_f1t[15]_i_4__2_n_0 ),
        .O(\r_f1t[11]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6966996969996669)) 
    \r_f1t[11]_i_4__1 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [19]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [19]),
        .I2(\r_f1t[15]_i_8_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [18]),
        .I4(\u_geo/u_geo_matrix/w_m1_out [18]),
        .I5(\r_exp_1z[3]_i_2_n_0 ),
        .O(\r_f1t[11]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6966996969996669)) 
    \r_f1t[11]_i_4__2 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [19]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [19]),
        .I2(\r_f1t[15]_i_8__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [18]),
        .I4(\u_geo/u_geo_matrix/w_m3_out [18]),
        .I5(\r_exp_1z[3]_i_2__0_n_0 ),
        .O(\r_f1t[11]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6966996969996669)) 
    \r_f1t[11]_i_4__3 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [19]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [19]),
        .I2(\r_f1t[15]_i_8__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [18]),
        .I4(\u_geo/u_geo_matrix/w_add23_out [18]),
        .I5(\r_exp_1z[3]_i_2__1_n_0 ),
        .O(\r_f1t[11]_i_4__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \r_f1t[11]_i_5 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [18]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [18]),
        .I2(\r_f1t[15]_i_8_n_0 ),
        .O(\r_f1t[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \r_f1t[11]_i_5__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [18]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [18]),
        .I2(\r_f1t[15]_i_8__0_n_0 ),
        .O(\r_f1t[11]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h69)) 
    \r_f1t[11]_i_5__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [18]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [18]),
        .I2(\r_f1t[15]_i_8__1_n_0 ),
        .O(\r_f1t[11]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_f1t[11]_i_5__2 
       (.I0(\u_geo/u_geo_viewport/sel0 [2]),
        .I1(\u_geo/u_geo_viewport/sel0 [3]),
        .O(\r_f1t[11]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEFFFEF)) 
    \r_f1t[11]_i_5__3 
       (.I0(\r_f1t[15]_i_8__2_n_0 ),
        .I1(\r_f1t[15]_i_9_n_0 ),
        .I2(\u_geo/w_vw_clip [13]),
        .I3(\u_geo/w_state_clip ),
        .I4(\u_geo/w_vw_mvp [13]),
        .O(\r_f1t[11]_i_5__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[11]_i_6 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [13]),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[11]_i_4__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [11]),
        .I4(\r_f1t[11]_i_5_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m0_out [15]),
        .O(\r_f1t[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[11]_i_6__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [13]),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[11]_i_4__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [11]),
        .I4(\r_f1t[11]_i_5__0_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m2_out [15]),
        .O(\r_f1t[11]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFCF4F7FFFFF4F7)) 
    \r_f1t[11]_i_6__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [13]),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[11]_i_4__3_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [11]),
        .I4(\r_f1t[11]_i_5__1_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_add01_out [15]),
        .O(\r_f1t[11]_i_6__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBABABABFBFBFB)) 
    \r_f1t[11]_i_6__2 
       (.I0(\r_f1t[15]_i_9_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [11]),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\u_geo/w_vw_mvp [15]),
        .I4(\u_geo/w_state_clip ),
        .I5(\u_geo/u_geo_clip/r_vw_reg_n_0_ ),
        .O(\r_f1t[11]_i_6__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[12]_i_1 
       (.I0(\r_f1t[13]_i_3_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[12]_i_2_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[12]_i_3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[12]_i_1__0 
       (.I0(\r_f1t[13]_i_3__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\r_f1t[12]_i_2__0_n_0 ),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[12]_i_3__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[12]_i_1__1 
       (.I0(\r_f1t[13]_i_3__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[12]_i_2__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[12]_i_3__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF000047470000)) 
    \r_f1t[12]_i_1__2 
       (.I0(\r_f1t[13]_i_2__2_n_0 ),
        .I1(\r_f0[15]_i_2__3_n_0 ),
        .I2(\r_f1t[12]_i_2__2_n_0 ),
        .I3(\r_f1t[12]_i_3__2_n_0 ),
        .I4(\r_f1t[15]_i_5_n_0 ),
        .I5(\r_f1t[15]_i_6__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[12]_i_1__3 
       (.I0(\r_f1t[12]_i_2__3_n_0 ),
        .I1(\r_f1t[14]_i_3__3_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[12]_i_3__3_n_0 ),
        .I4(\r_f1t[12]_i_4__2_n_0 ),
        .I5(\r_f1t[13]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \r_f1t[12]_i_2 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [14]),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f0[15]_i_3_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m1_out [12]),
        .O(\r_f1t[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \r_f1t[12]_i_2__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [14]),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f0[15]_i_3__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m3_out [12]),
        .O(\r_f1t[12]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \r_f1t[12]_i_2__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [14]),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f0[15]_i_3__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add23_out [12]),
        .O(\r_f1t[12]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF4FFF7)) 
    \r_f1t[12]_i_2__2 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [15]),
        .I1(\r_f1t[15]_i_2_n_0 ),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\r_f1t[15]_i_9_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [13]),
        .O(\r_f1t[12]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \r_f1t[12]_i_2__3 
       (.I0(\u_geo/u_geo_viewport/sel0 [0]),
        .I1(\u_geo/u_geo_viewport/sel0 [1]),
        .I2(\u_geo/u_geo_viewport/sel0 [4]),
        .O(\r_f1t[12]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \r_f1t[12]_i_3 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [14]),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f0[15]_i_3_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [12]),
        .I4(\r_f1t[15]_i_5__0_n_0 ),
        .I5(\r_f1t[12]_i_4_n_0 ),
        .O(\r_f1t[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \r_f1t[12]_i_3__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [14]),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f0[15]_i_3__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [12]),
        .I4(\r_f1t[15]_i_5__1_n_0 ),
        .I5(\r_f1t[12]_i_4__0_n_0 ),
        .O(\r_f1t[12]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \r_f1t[12]_i_3__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [14]),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f0[15]_i_3__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [12]),
        .I4(\r_f1t[15]_i_5__2_n_0 ),
        .I5(\r_f1t[12]_i_4__1_n_0 ),
        .O(\r_f1t[12]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[12]_i_3__2 
       (.I0(\r_f1t[14]_i_4__0_n_0 ),
        .I1(\r_f1t[12]_i_4__3_n_0 ),
        .I2(\r_f0[15]_i_2__3_n_0 ),
        .I3(\r_f1t[13]_i_4__3_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[12]_i_5_n_0 ),
        .O(\r_f1t[12]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FF0000B8000000)) 
    \r_f1t[12]_i_3__3 
       (.I0(\u_geo/w_vx_pdiv [15]),
        .I1(\r_f0[15]_i_2_n_0 ),
        .I2(\u_geo/w_vy_pdiv [15]),
        .I3(\u_geo/u_geo_viewport/sel0 [1]),
        .I4(\r_f1t[15]_i_4__2_n_0 ),
        .I5(\u_geo/u_geo_viewport/w_fadd_a [13]),
        .O(\r_f1t[12]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \r_f1t[12]_i_4 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [15]),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f0[15]_i_3_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [13]),
        .O(\r_f1t[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \r_f1t[12]_i_4__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [15]),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f0[15]_i_3__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [13]),
        .O(\r_f1t[12]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \r_f1t[12]_i_4__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [15]),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f0[15]_i_3__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [13]),
        .O(\r_f1t[12]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FF0000B8000000)) 
    \r_f1t[12]_i_4__2 
       (.I0(\u_geo/w_vx_pdiv [14]),
        .I1(\r_f0[15]_i_2_n_0 ),
        .I2(\u_geo/w_vy_pdiv [14]),
        .I3(\u_geo/u_geo_viewport/sel0 [1]),
        .I4(\r_f1t[15]_i_4__2_n_0 ),
        .I5(\u_geo/u_geo_viewport/w_fadd_a [12]),
        .O(\r_f1t[12]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \r_f1t[12]_i_4__3 
       (.I0(\r_f1t[15]_i_8__2_n_0 ),
        .I1(\r_f1t[15]_i_9_n_0 ),
        .I2(\r_f0[12]_i_2_n_0 ),
        .O(\r_f1t[12]_i_4__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEFFFEF)) 
    \r_f1t[12]_i_5 
       (.I0(\r_f1t[15]_i_8__2_n_0 ),
        .I1(\r_f1t[15]_i_9_n_0 ),
        .I2(\u_geo/w_vw_clip [12]),
        .I3(\u_geo/w_state_clip ),
        .I4(\u_geo/w_vw_mvp [12]),
        .O(\r_f1t[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[13]_i_1 
       (.I0(\r_f1t[13]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[13]_i_3_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[13]_i_4_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[13]_i_1__0 
       (.I0(\r_f1t[13]_i_2__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\r_f1t[13]_i_3__0_n_0 ),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[13]_i_4__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[13]_i_1__1 
       (.I0(\r_f1t[13]_i_2__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[13]_i_3__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[13]_i_4__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[13]_i_1__2 
       (.I0(\r_f1t[14]_i_2__2_n_0 ),
        .I1(\r_f1t[15]_i_6__2_n_0 ),
        .I2(\r_f1t[13]_i_2__2_n_0 ),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f1t[15]_i_5_n_0 ),
        .I5(\r_f1t[13]_i_3__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88F888FF88F888F8)) 
    \r_f1t[13]_i_1__3 
       (.I0(\r_f1t[14]_i_3__3_n_0 ),
        .I1(\r_f1t[13]_i_2__3_n_0 ),
        .I2(\r_f1t[13]_i_3__3_n_0 ),
        .I3(\r_f1t[13]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/sel0 [1]),
        .I5(\r_f1t[13]_i_5_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    \r_f1t[13]_i_2 
       (.I0(\r_f1t[15]_i_4_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [14]),
        .I2(\r_f0[15]_i_3_n_0 ),
        .O(\r_f1t[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    \r_f1t[13]_i_2__0 
       (.I0(\r_f1t[15]_i_4__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [14]),
        .I2(\r_f0[15]_i_3__0_n_0 ),
        .O(\r_f1t[13]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    \r_f1t[13]_i_2__1 
       (.I0(\r_f1t[15]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [14]),
        .I2(\r_f0[15]_i_3__1_n_0 ),
        .O(\r_f1t[13]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF4FFF7)) 
    \r_f1t[13]_i_2__2 
       (.I0(\r_f0[15]_i_3__2_n_0 ),
        .I1(\r_f1t[15]_i_2_n_0 ),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\r_f1t[15]_i_9_n_0 ),
        .I4(\r_f0[13]_i_2_n_0 ),
        .O(\r_f1t[13]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \r_f1t[13]_i_2__3 
       (.I0(\u_geo/u_geo_viewport/sel0 [0]),
        .I1(\u_geo/u_geo_viewport/sel0 [1]),
        .I2(\u_geo/u_geo_viewport/sel0 [4]),
        .O(\r_f1t[13]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \r_f1t[13]_i_3 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [15]),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f0[15]_i_3_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m1_out [13]),
        .O(\r_f1t[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \r_f1t[13]_i_3__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [15]),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f0[15]_i_3__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m3_out [13]),
        .O(\r_f1t[13]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \r_f1t[13]_i_3__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [15]),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f0[15]_i_3__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add23_out [13]),
        .O(\r_f1t[13]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBBB8)) 
    \r_f1t[13]_i_3__2 
       (.I0(\r_f1t[12]_i_2__2_n_0 ),
        .I1(\r_f1t[15]_i_6__2_n_0 ),
        .I2(\r_f1t[15]_i_2_n_0 ),
        .I3(\r_f1t[13]_i_4__3_n_0 ),
        .O(\r_f1t[13]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000C808)) 
    \r_f1t[13]_i_3__3 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [13]),
        .I1(\r_f1t[15]_i_4__2_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [1]),
        .I3(\u_geo/u_geo_viewport/w_fadd_a [15]),
        .I4(\u_geo/u_geo_viewport/sel0 [0]),
        .O(\r_f1t[13]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF5F305F3F)) 
    \r_f1t[13]_i_4 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [15]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [13]),
        .I2(\r_f1t[15]_i_5__0_n_0 ),
        .I3(\r_f1t[15]_i_4_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m0_out [14]),
        .I5(\r_f0[15]_i_3_n_0 ),
        .O(\r_f1t[13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF5F305F3F)) 
    \r_f1t[13]_i_4__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [15]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [13]),
        .I2(\r_f1t[15]_i_5__1_n_0 ),
        .I3(\r_f1t[15]_i_4__0_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m2_out [14]),
        .I5(\r_f0[15]_i_3__0_n_0 ),
        .O(\r_f1t[13]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF5F305F3F)) 
    \r_f1t[13]_i_4__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [15]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [13]),
        .I2(\r_f1t[15]_i_5__2_n_0 ),
        .I3(\r_f1t[15]_i_4__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add01_out [14]),
        .I5(\r_f0[15]_i_3__1_n_0 ),
        .O(\r_f1t[13]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r_f1t[13]_i_4__2 
       (.I0(\u_geo/u_geo_viewport/sel0 [4]),
        .I1(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ),
        .O(\r_f1t[13]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEFFFEF)) 
    \r_f1t[13]_i_4__3 
       (.I0(\r_f1t[15]_i_8__2_n_0 ),
        .I1(\r_f1t[15]_i_9_n_0 ),
        .I2(\u_geo/w_vw_clip [14]),
        .I3(\u_geo/w_state_clip ),
        .I4(\u_geo/w_vw_mvp [14]),
        .O(\r_f1t[13]_i_4__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hE2000000)) 
    \r_f1t[13]_i_5 
       (.I0(\u_geo/w_vy_pdiv [14]),
        .I1(\r_f0[15]_i_2_n_0 ),
        .I2(\u_geo/w_vx_pdiv [14]),
        .I3(\r_f1t[15]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/sel0 [0]),
        .O(\r_f1t[13]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[14]_i_1 
       (.I0(\r_f1t[15]_i_4__3_n_0 ),
        .I1(\r_f1t[15]_i_6__2_n_0 ),
        .I2(\r_f1t[14]_i_2__2_n_0 ),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f1t[15]_i_5_n_0 ),
        .I5(\r_f1t[14]_i_3__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[14]_i_1__0 
       (.I0(\r_f1t[14]_i_2__3_n_0 ),
        .I1(\r_f1t[14]_i_3__3_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[14]_i_4_n_0 ),
        .I4(\r_f1t[14]_i_5_n_0 ),
        .I5(\r_f1t[14]_i_6_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0022002000000020)) 
    \r_f1t[14]_i_2 
       (.I0(\r_f1t[15]_i_6_n_0 ),
        .I1(\r_f0[15]_i_3_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m0_out [15]),
        .I3(\r_f1t[15]_i_4_n_0 ),
        .I4(\r_f1t[15]_i_5__0_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m0_out [14]),
        .O(\r_f1t[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0022002000000020)) 
    \r_f1t[14]_i_2__0 
       (.I0(\r_f1t[15]_i_6__0_n_0 ),
        .I1(\r_f0[15]_i_3__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m2_out [15]),
        .I3(\r_f1t[15]_i_4__0_n_0 ),
        .I4(\r_f1t[15]_i_5__1_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m2_out [14]),
        .O(\r_f1t[14]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0022002000000020)) 
    \r_f1t[14]_i_2__1 
       (.I0(\r_f1t[15]_i_6__1_n_0 ),
        .I1(\r_f0[15]_i_3__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add01_out [15]),
        .I3(\r_f1t[15]_i_4__1_n_0 ),
        .I4(\r_f1t[15]_i_5__2_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_add01_out [14]),
        .O(\r_f1t[14]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_f1t[14]_i_2__2 
       (.I0(\r_f1t[15]_i_2_n_0 ),
        .I1(\r_f1t[14]_i_4__0_n_0 ),
        .O(\r_f1t[14]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \r_f1t[14]_i_2__3 
       (.I0(\u_geo/u_geo_viewport/sel0 [1]),
        .I1(\u_geo/u_geo_viewport/sel0 [0]),
        .I2(\u_geo/u_geo_viewport/sel0 [4]),
        .O(\r_f1t[14]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0022002000000020)) 
    \r_f1t[14]_i_3 
       (.I0(\r_f1t[15]_i_6_n_0 ),
        .I1(\r_f0[15]_i_3_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [15]),
        .I3(\r_f1t[15]_i_4_n_0 ),
        .I4(\r_f1t[15]_i_5__0_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m1_out [14]),
        .O(\r_f1t[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0022002000000020)) 
    \r_f1t[14]_i_3__0 
       (.I0(\r_f1t[15]_i_6__0_n_0 ),
        .I1(\r_f0[15]_i_3__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [15]),
        .I3(\r_f1t[15]_i_4__0_n_0 ),
        .I4(\r_f1t[15]_i_5__1_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_m3_out [14]),
        .O(\r_f1t[14]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0022002000000020)) 
    \r_f1t[14]_i_3__1 
       (.I0(\r_f1t[15]_i_6__1_n_0 ),
        .I1(\r_f0[15]_i_3__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [15]),
        .I3(\r_f1t[15]_i_4__1_n_0 ),
        .I4(\r_f1t[15]_i_5__2_n_0 ),
        .I5(\u_geo/u_geo_matrix/w_add23_out [14]),
        .O(\r_f1t[14]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F7)) 
    \r_f1t[14]_i_3__2 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [14]),
        .I1(\r_f1t[15]_i_6__2_n_0 ),
        .I2(\r_f1t[15]_i_2_n_0 ),
        .I3(\u_geo/u_geo_clip/w_add_in_a [15]),
        .I4(\r_f1t[15]_i_9_n_0 ),
        .I5(\r_f1t[15]_i_8__2_n_0 ),
        .O(\r_f1t[14]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_f1t[14]_i_3__3 
       (.I0(\r_f1t[15]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ),
        .O(\r_f1t[14]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8A80)) 
    \r_f1t[14]_i_4 
       (.I0(\r_f1t[15]_i_4__2_n_0 ),
        .I1(\u_geo/w_vx_pdiv [15]),
        .I2(\r_f0[15]_i_2_n_0 ),
        .I3(\u_geo/w_vy_pdiv [15]),
        .O(\r_f1t[14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \r_f1t[14]_i_4__0 
       (.I0(\r_f1t[15]_i_8__2_n_0 ),
        .I1(\r_f1t[15]_i_9_n_0 ),
        .I2(\r_f0[14]_i_2_n_0 ),
        .O(\r_f1t[14]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8A80)) 
    \r_f1t[14]_i_5 
       (.I0(\r_f1t[15]_i_4__2_n_0 ),
        .I1(\u_geo/w_vx_pdiv [14]),
        .I2(\r_f0[15]_i_2_n_0 ),
        .I3(\u_geo/w_vy_pdiv [14]),
        .O(\r_f1t[14]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFD)) 
    \r_f1t[14]_i_6 
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ),
        .I1(\u_geo/u_geo_viewport/sel0 [4]),
        .I2(\u_geo/u_geo_viewport/sel0 [1]),
        .O(\r_f1t[14]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0047000000000000)) 
    \r_f1t[15]_i_1 
       (.I0(\r_f1t[15]_i_2__1_n_0 ),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\r_f1t[15]_i_3__0_n_0 ),
        .I3(\r_f1t[15]_i_4_n_0 ),
        .I4(\r_f1t[15]_i_5__0_n_0 ),
        .I5(\r_f1t[15]_i_6_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[15]_i_10 
       (.I0(\u_geo/w_vw_mvp [19]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [19]),
        .O(\u_geo/u_geo_clip/w_add_in_a [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4D44DD4D2BBB222B)) 
    \r_f1t[15]_i_11 
       (.I0(\r_exp_1z[2]_i_2_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [18]),
        .I2(\r_f1t[15]_i_12_n_0 ),
        .I3(\u_geo/u_geo_clip/w_add_in_a [17]),
        .I4(\r_exp_1z[1]_i_2_n_0 ),
        .I5(\r_exp_1z[3]_i_3__2_n_0 ),
        .O(\r_f1t[15]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAEFFAAAEF755FFF7)) 
    \r_f1t[15]_i_12 
       (.I0(\r_exp_1z[0]_i_2_n_0 ),
        .I1(\r_exp_1z[0]_i_5_n_0 ),
        .I2(\r_exp_1z[0]_i_4_n_0 ),
        .I3(\r_exp_1z[4]_i_2_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [20]),
        .I5(\u_geo/u_geo_clip/w_add_in_a [16]),
        .O(\r_f1t[15]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0047000000000000)) 
    \r_f1t[15]_i_1__0 
       (.I0(\r_f1t[15]_i_2__2_n_0 ),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\r_f1t[15]_i_3__1_n_0 ),
        .I3(\r_f1t[15]_i_4__0_n_0 ),
        .I4(\r_f1t[15]_i_5__1_n_0 ),
        .I5(\r_f1t[15]_i_6__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0047000000000000)) 
    \r_f1t[15]_i_1__1 
       (.I0(\r_f1t[15]_i_2__3_n_0 ),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\r_f1t[15]_i_3__2_n_0 ),
        .I3(\r_f1t[15]_i_4__1_n_0 ),
        .I4(\r_f1t[15]_i_5__2_n_0 ),
        .I5(\r_f1t[15]_i_6__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0002000000030000)) 
    \r_f1t[15]_i_1__2 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [15]),
        .I1(\u_geo/u_geo_viewport/sel0 [0]),
        .I2(\u_geo/u_geo_viewport/sel0 [1]),
        .I3(\u_geo/u_geo_viewport/sel0 [4]),
        .I4(\r_f1t[15]_i_4__2_n_0 ),
        .I5(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ),
        .O(\u_geo/u_geo_viewport/w_f1t [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F11000000000000)) 
    \r_f1t[15]_i_1__3 
       (.I0(\r_f1t[15]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_3__3_n_0 ),
        .I2(\r_f1t[15]_i_4__3_n_0 ),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f1t[15]_i_5_n_0 ),
        .I5(\r_f1t[15]_i_6__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555656A9A955555)) 
    \r_f1t[15]_i_2 
       (.I0(\r_f1t[15]_i_7__2_n_0 ),
        .I1(\u_geo/w_vw_mvp [16]),
        .I2(\u_geo/w_state_clip ),
        .I3(\u_geo/w_vw_clip [16]),
        .I4(\r_exp_1z[3]_i_3__2_n_0 ),
        .I5(\r_exp_1z[0]_i_2_n_0 ),
        .O(\r_f1t[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    \r_f1t[15]_i_2__0 
       (.I0(\u_geo/w_vy_pdiv [15]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [15]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r_f1t[15]_i_2__1 
       (.I0(\r_f0[15]_i_3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [15]),
        .O(\r_f1t[15]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r_f1t[15]_i_2__2 
       (.I0(\r_f0[15]_i_3__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [15]),
        .O(\r_f1t[15]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r_f1t[15]_i_2__3 
       (.I0(\r_f0[15]_i_3__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [15]),
        .O(\r_f1t[15]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h1B)) 
    \r_f1t[15]_i_3 
       (.I0(\r_f0[15]_i_2_n_0 ),
        .I1(\u_geo/w_vy_pdiv [16]),
        .I2(\u_geo/w_vx_pdiv [16]),
        .O(\u_geo/u_geo_viewport/sel0 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r_f1t[15]_i_3__0 
       (.I0(\r_f0[15]_i_3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [15]),
        .O(\r_f1t[15]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r_f1t[15]_i_3__1 
       (.I0(\r_f0[15]_i_3__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [15]),
        .O(\r_f1t[15]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r_f1t[15]_i_3__2 
       (.I0(\r_f0[15]_i_3__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [15]),
        .O(\r_f1t[15]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEFFFEF)) 
    \r_f1t[15]_i_3__3 
       (.I0(\r_f1t[15]_i_8__2_n_0 ),
        .I1(\r_f1t[15]_i_9_n_0 ),
        .I2(\u_geo/u_geo_clip/r_vw_reg_n_0_ ),
        .I3(\u_geo/w_state_clip ),
        .I4(\u_geo/w_vw_mvp [15]),
        .O(\r_f1t[15]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66699666)) 
    \r_f1t[15]_i_4 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [17]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [17]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [16]),
        .I3(\r_exp_1z[3]_i_2_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m1_out [16]),
        .O(\r_f1t[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66699666)) 
    \r_f1t[15]_i_4__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [17]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [17]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [16]),
        .I3(\r_exp_1z[3]_i_2__0_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m3_out [16]),
        .O(\r_f1t[15]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66699666)) 
    \r_f1t[15]_i_4__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [17]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [17]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [16]),
        .I3(\r_exp_1z[3]_i_2__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add23_out [16]),
        .O(\r_f1t[15]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r_f1t[15]_i_4__2 
       (.I0(\u_geo/u_geo_viewport/sel0 [3]),
        .I1(\u_geo/u_geo_viewport/sel0 [2]),
        .O(\r_f1t[15]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    \r_f1t[15]_i_4__3 
       (.I0(\r_f1t[15]_i_8__2_n_0 ),
        .I1(\r_f1t[15]_i_9_n_0 ),
        .I2(\r_f0[15]_i_3__2_n_0 ),
        .I3(\r_f1t[15]_i_2_n_0 ),
        .O(\r_f1t[15]_i_4__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF99FFF99F99F99)) 
    \r_f1t[15]_i_5 
       (.I0(\r_exp_1z[4]_i_2_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [20]),
        .I2(\r_exp_1z[3]_i_3__2_n_0 ),
        .I3(\r_exp_1z[3]_i_2__2_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [19]),
        .I5(\r_f1t[15]_i_11_n_0 ),
        .O(\r_f1t[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r_f1t[15]_i_5__0 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [16]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [16]),
        .O(\r_f1t[15]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r_f1t[15]_i_5__1 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [16]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [16]),
        .O(\r_f1t[15]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r_f1t[15]_i_5__2 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [16]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [16]),
        .O(\r_f1t[15]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF99FFF99F99F99)) 
    \r_f1t[15]_i_6 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [20]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [20]),
        .I2(\r_exp_1z[3]_i_2_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m1_out [19]),
        .I4(\u_geo/u_geo_matrix/w_m0_out [19]),
        .I5(\r_f1t[15]_i_7_n_0 ),
        .O(\r_f1t[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF99FFF99F99F99)) 
    \r_f1t[15]_i_6__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [20]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [20]),
        .I2(\r_exp_1z[3]_i_2__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m3_out [19]),
        .I4(\u_geo/u_geo_matrix/w_m2_out [19]),
        .I5(\r_f1t[15]_i_7__0_n_0 ),
        .O(\r_f1t[15]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF99FFF99F99F99)) 
    \r_f1t[15]_i_6__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [20]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [20]),
        .I2(\r_exp_1z[3]_i_2__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add23_out [19]),
        .I4(\u_geo/u_geo_matrix/w_add01_out [19]),
        .I5(\r_f1t[15]_i_7__1_n_0 ),
        .O(\r_f1t[15]_i_6__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE21D)) 
    \r_f1t[15]_i_6__2 
       (.I0(\u_geo/w_vw_clip [16]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_mvp [16]),
        .I3(\r_exp_1z[0]_i_2_n_0 ),
        .O(\r_f1t[15]_i_6__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h24E7)) 
    \r_f1t[15]_i_7 
       (.I0(\r_exp_1z[3]_i_2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [18]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [18]),
        .I3(\r_f1t[15]_i_8_n_0 ),
        .O(\r_f1t[15]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h24E7)) 
    \r_f1t[15]_i_7__0 
       (.I0(\r_exp_1z[3]_i_2__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [18]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [18]),
        .I3(\r_f1t[15]_i_8__0_n_0 ),
        .O(\r_f1t[15]_i_7__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h24E7)) 
    \r_f1t[15]_i_7__1 
       (.I0(\r_exp_1z[3]_i_2__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [18]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [18]),
        .I3(\r_f1t[15]_i_8__1_n_0 ),
        .O(\r_f1t[15]_i_7__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB847)) 
    \r_f1t[15]_i_7__2 
       (.I0(\u_geo/w_vw_mvp [17]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [17]),
        .I3(\r_exp_1z[1]_i_2_n_0 ),
        .O(\r_f1t[15]_i_7__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBF0BD0FD)) 
    \r_f1t[15]_i_8 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [16]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [16]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [17]),
        .I3(\u_geo/u_geo_matrix/w_m1_out [17]),
        .I4(\r_exp_1z[3]_i_2_n_0 ),
        .O(\r_f1t[15]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBF0BD0FD)) 
    \r_f1t[15]_i_8__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [16]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [16]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [17]),
        .I3(\u_geo/u_geo_matrix/w_m3_out [17]),
        .I4(\r_exp_1z[3]_i_2__0_n_0 ),
        .O(\r_f1t[15]_i_8__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBF0BD0FD)) 
    \r_f1t[15]_i_8__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [16]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [16]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [17]),
        .I3(\u_geo/u_geo_matrix/w_add23_out [17]),
        .I4(\r_exp_1z[3]_i_2__1_n_0 ),
        .O(\r_f1t[15]_i_8__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5965696699695965)) 
    \r_f1t[15]_i_8__2 
       (.I0(\r_f0[15]_i_11_n_0 ),
        .I1(\r_exp_1z[3]_i_3__2_n_0 ),
        .I2(\r_exp_1z[1]_i_2_n_0 ),
        .I3(\u_geo/u_geo_clip/w_add_in_a [17]),
        .I4(\u_geo/u_geo_clip/w_add_in_a [16]),
        .I5(\r_exp_1z[0]_i_2_n_0 ),
        .O(\r_f1t[15]_i_8__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A55AA9A9AAA559A)) 
    \r_f1t[15]_i_9 
       (.I0(\r_f0[15]_i_9_n_0 ),
        .I1(\r_f0[15]_i_13_n_0 ),
        .I2(\r_f0[15]_i_12_n_0 ),
        .I3(\u_geo/u_geo_clip/w_add_in_a [18]),
        .I4(\r_exp_1z[2]_i_2_n_0 ),
        .I5(\r_exp_1z[3]_i_3__2_n_0 ),
        .O(\r_f1t[15]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[1]_i_1 
       (.I0(\r_f1t[2]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[1]_i_2_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[1]_i_3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[1]_i_1__0 
       (.I0(\r_f1t[2]_i_2__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\r_f1t[1]_i_2__0_n_0 ),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[1]_i_3__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[1]_i_1__1 
       (.I0(\r_f1t[2]_i_2__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[1]_i_2__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[1]_i_3__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[1]_i_1__2 
       (.I0(\r_f1t[2]_i_2__2_n_0 ),
        .I1(\r_f1t[15]_i_6__2_n_0 ),
        .I2(\r_f1t[1]_i_2__2_n_0 ),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f1t[15]_i_5_n_0 ),
        .I5(\r_f1t[1]_i_3__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[1]_i_1__3 
       (.I0(\r_f1t[13]_i_2__3_n_0 ),
        .I1(\r_f1t[3]_i_2__3_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[2]_i_2__3_n_0 ),
        .I4(\r_f1t[1]_i_2__3_n_0 ),
        .I5(\r_f1t[13]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[1]_i_2 
       (.I0(\r_f1t[3]_i_4__1_n_0 ),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[1]_i_4__1_n_0 ),
        .O(\r_f1t[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[1]_i_2__0 
       (.I0(\r_f1t[3]_i_4__2_n_0 ),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[1]_i_4__2_n_0 ),
        .O(\r_f1t[1]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[1]_i_2__1 
       (.I0(\r_f1t[3]_i_4__3_n_0 ),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[1]_i_4__3_n_0 ),
        .O(\r_f1t[1]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[1]_i_2__2 
       (.I0(\r_f1t[3]_i_4_n_0 ),
        .I1(\r_f1t[15]_i_2_n_0 ),
        .I2(\r_f1t[1]_i_4_n_0 ),
        .O(\r_f1t[1]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBB8B8B8)) 
    \r_f1t[1]_i_2__3 
       (.I0(\r_f1t[3]_i_4__0_n_0 ),
        .I1(\u_geo/u_geo_viewport/sel0 [1]),
        .I2(\r_f1t[1]_i_3__3_n_0 ),
        .I3(\u_geo/u_geo_viewport/sel0 [2]),
        .I4(\r_f1t[1]_i_4__0_n_0 ),
        .O(\r_f1t[1]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[1]_i_3 
       (.I0(\r_f1t[3]_i_5__0_n_0 ),
        .I1(\r_f1t[1]_i_5__0_n_0 ),
        .I2(\r_f1t[15]_i_5__0_n_0 ),
        .I3(\r_f1t[2]_i_5_n_0 ),
        .I4(\r_f1t[15]_i_4_n_0 ),
        .I5(\r_f1t[2]_i_6_n_0 ),
        .O(\r_f1t[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[1]_i_3__0 
       (.I0(\r_f1t[3]_i_5__1_n_0 ),
        .I1(\r_f1t[1]_i_5__1_n_0 ),
        .I2(\r_f1t[15]_i_5__1_n_0 ),
        .I3(\r_f1t[2]_i_5__0_n_0 ),
        .I4(\r_f1t[15]_i_4__0_n_0 ),
        .I5(\r_f1t[2]_i_6__0_n_0 ),
        .O(\r_f1t[1]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[1]_i_3__1 
       (.I0(\r_f1t[3]_i_5__2_n_0 ),
        .I1(\r_f1t[1]_i_5__2_n_0 ),
        .I2(\r_f1t[15]_i_5__2_n_0 ),
        .I3(\r_f1t[2]_i_5__1_n_0 ),
        .I4(\r_f1t[15]_i_4__1_n_0 ),
        .I5(\r_f1t[2]_i_6__1_n_0 ),
        .O(\r_f1t[1]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[1]_i_3__2 
       (.I0(\r_f1t[3]_i_5_n_0 ),
        .I1(\r_f1t[1]_i_5_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[4]_i_5__2_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[2]_i_5__2_n_0 ),
        .O(\r_f1t[1]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000AAAAFC0C)) 
    \r_f1t[1]_i_3__3 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [9]),
        .I1(\u_geo/w_vy_pdiv [1]),
        .I2(\r_f0[15]_i_2_n_0 ),
        .I3(\u_geo/w_vx_pdiv [1]),
        .I4(\u_geo/u_geo_viewport/sel0 [3]),
        .I5(\u_geo/u_geo_viewport/sel0 [2]),
        .O(\r_f1t[1]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3030505F3F3F505F)) 
    \r_f1t[1]_i_4 
       (.I0(\r_f0[5]_i_2_n_0 ),
        .I1(\r_f0[13]_i_2_n_0 ),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\r_f0[1]_i_2_n_0 ),
        .I4(\r_f1t[15]_i_9_n_0 ),
        .I5(\r_f0[9]_i_2_n_0 ),
        .O(\r_f1t[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFAFA0C0C0AFA0)) 
    \r_f1t[1]_i_4__0 
       (.I0(\u_geo/w_vy_pdiv [13]),
        .I1(\u_geo/w_vx_pdiv [13]),
        .I2(\u_geo/u_geo_viewport/sel0 [3]),
        .I3(\u_geo/w_vy_pdiv [5]),
        .I4(\r_f0[15]_i_2_n_0 ),
        .I5(\u_geo/w_vx_pdiv [5]),
        .O(\r_f1t[1]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[1]_i_4__1 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [5]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [13]),
        .I3(\r_f1t[11]_i_5_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m1_out [1]),
        .I5(\u_geo/u_geo_matrix/w_m1_out [9]),
        .O(\r_f1t[1]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[1]_i_4__2 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [5]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [13]),
        .I3(\r_f1t[11]_i_5__0_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m3_out [1]),
        .I5(\u_geo/u_geo_matrix/w_m3_out [9]),
        .O(\r_f1t[1]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[1]_i_4__3 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [5]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [13]),
        .I3(\r_f1t[11]_i_5__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add23_out [1]),
        .I5(\u_geo/u_geo_matrix/w_add23_out [9]),
        .O(\r_f1t[1]_i_4__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3030505F3F3F505F)) 
    \r_f1t[1]_i_5 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [5]),
        .I1(\u_geo/u_geo_clip/w_add_in_a [13]),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\u_geo/u_geo_clip/w_add_in_a [1]),
        .I4(\r_f1t[15]_i_9_n_0 ),
        .I5(\u_geo/u_geo_clip/w_add_in_a [9]),
        .O(\r_f1t[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[1]_i_5__0 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [5]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [13]),
        .I3(\r_f1t[11]_i_5_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m0_out [1]),
        .I5(\u_geo/u_geo_matrix/w_m0_out [9]),
        .O(\r_f1t[1]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[1]_i_5__1 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [5]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [13]),
        .I3(\r_f1t[11]_i_5__0_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m2_out [1]),
        .I5(\u_geo/u_geo_matrix/w_m2_out [9]),
        .O(\r_f1t[1]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[1]_i_5__2 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [5]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [13]),
        .I3(\r_f1t[11]_i_5__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add01_out [1]),
        .I5(\u_geo/u_geo_matrix/w_add01_out [9]),
        .O(\r_f1t[1]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[2]_i_1 
       (.I0(\r_f1t[3]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[2]_i_2_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[2]_i_3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[2]_i_1__0 
       (.I0(\r_f1t[3]_i_2__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\r_f1t[2]_i_2__0_n_0 ),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[2]_i_3__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[2]_i_1__1 
       (.I0(\r_f1t[3]_i_2__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[2]_i_2__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[2]_i_3__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[2]_i_1__2 
       (.I0(\r_f1t[3]_i_2__2_n_0 ),
        .I1(\r_f1t[15]_i_6__2_n_0 ),
        .I2(\r_f1t[2]_i_2__2_n_0 ),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f1t[15]_i_5_n_0 ),
        .I5(\r_f1t[2]_i_3__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[2]_i_1__3 
       (.I0(\r_f1t[14]_i_2__3_n_0 ),
        .I1(\r_f1t[3]_i_2__3_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[3]_i_3__3_n_0 ),
        .I4(\r_f1t[2]_i_2__3_n_0 ),
        .I5(\r_f1t[13]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[2]_i_2 
       (.I0(\r_f1t[4]_i_4_n_0 ),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[2]_i_4__0_n_0 ),
        .O(\r_f1t[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[2]_i_2__0 
       (.I0(\r_f1t[4]_i_4__0_n_0 ),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[2]_i_4__1_n_0 ),
        .O(\r_f1t[2]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[2]_i_2__1 
       (.I0(\r_f1t[4]_i_4__1_n_0 ),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[2]_i_4__2_n_0 ),
        .O(\r_f1t[2]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[2]_i_2__2 
       (.I0(\r_f1t[4]_i_4__2_n_0 ),
        .I1(\r_f1t[15]_i_2_n_0 ),
        .I2(\r_f1t[2]_i_4_n_0 ),
        .O(\r_f1t[2]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[2]_i_2__3 
       (.I0(\r_f1t[4]_i_3__0_n_0 ),
        .I1(\u_geo/u_geo_viewport/sel0 [1]),
        .I2(\r_f1t[2]_i_3__3_n_0 ),
        .O(\r_f1t[2]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[2]_i_3 
       (.I0(\r_f1t[2]_i_5_n_0 ),
        .I1(\r_f1t[2]_i_6_n_0 ),
        .I2(\r_f1t[15]_i_5__0_n_0 ),
        .I3(\r_f1t[5]_i_6_n_0 ),
        .I4(\r_f1t[15]_i_4_n_0 ),
        .I5(\r_f1t[3]_i_5__0_n_0 ),
        .O(\r_f1t[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[2]_i_3__0 
       (.I0(\r_f1t[2]_i_5__0_n_0 ),
        .I1(\r_f1t[2]_i_6__0_n_0 ),
        .I2(\r_f1t[15]_i_5__1_n_0 ),
        .I3(\r_f1t[5]_i_6__0_n_0 ),
        .I4(\r_f1t[15]_i_4__0_n_0 ),
        .I5(\r_f1t[3]_i_5__1_n_0 ),
        .O(\r_f1t[2]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[2]_i_3__1 
       (.I0(\r_f1t[2]_i_5__1_n_0 ),
        .I1(\r_f1t[2]_i_6__1_n_0 ),
        .I2(\r_f1t[15]_i_5__2_n_0 ),
        .I3(\r_f1t[5]_i_6__1_n_0 ),
        .I4(\r_f1t[15]_i_4__1_n_0 ),
        .I5(\r_f1t[3]_i_5__2_n_0 ),
        .O(\r_f1t[2]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[2]_i_3__2 
       (.I0(\r_f1t[4]_i_5__2_n_0 ),
        .I1(\r_f1t[2]_i_5__2_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[5]_i_5__2_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[3]_i_5_n_0 ),
        .O(\r_f1t[2]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \r_f1t[2]_i_3__3 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [2]),
        .I1(\u_geo/u_geo_viewport/w_fadd_a [10]),
        .I2(\u_geo/u_geo_viewport/sel0 [2]),
        .I3(\u_geo/u_geo_viewport/w_fadd_a [14]),
        .I4(\u_geo/u_geo_viewport/sel0 [3]),
        .I5(\u_geo/u_geo_viewport/w_fadd_a [6]),
        .O(\r_f1t[2]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3030505F3F3F505F)) 
    \r_f1t[2]_i_4 
       (.I0(\r_f0[6]_i_2_n_0 ),
        .I1(\r_f0[14]_i_2_n_0 ),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\r_f0[2]_i_2_n_0 ),
        .I4(\r_f1t[15]_i_9_n_0 ),
        .I5(\r_f0[10]_i_2_n_0 ),
        .O(\r_f1t[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[2]_i_4__0 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [6]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [14]),
        .I3(\r_f1t[11]_i_5_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m1_out [2]),
        .I5(\u_geo/u_geo_matrix/w_m1_out [10]),
        .O(\r_f1t[2]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[2]_i_4__1 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [6]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [14]),
        .I3(\r_f1t[11]_i_5__0_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m3_out [2]),
        .I5(\u_geo/u_geo_matrix/w_m3_out [10]),
        .O(\r_f1t[2]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[2]_i_4__2 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [6]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [14]),
        .I3(\r_f1t[11]_i_5__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add23_out [2]),
        .I5(\u_geo/u_geo_matrix/w_add23_out [10]),
        .O(\r_f1t[2]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[2]_i_5 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [8]),
        .I1(\r_f1t[11]_i_5_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m0_out [4]),
        .I3(\r_f1t[11]_i_4__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m0_out [12]),
        .O(\r_f1t[2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[2]_i_5__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [8]),
        .I1(\r_f1t[11]_i_5__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m2_out [4]),
        .I3(\r_f1t[11]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m2_out [12]),
        .O(\r_f1t[2]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[2]_i_5__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [8]),
        .I1(\r_f1t[11]_i_5__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add01_out [4]),
        .I3(\r_f1t[11]_i_4__3_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add01_out [12]),
        .O(\r_f1t[2]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3030505F3F3F505F)) 
    \r_f1t[2]_i_5__2 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [6]),
        .I1(\u_geo/u_geo_clip/w_add_in_a [14]),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\u_geo/u_geo_clip/w_add_in_a [2]),
        .I4(\r_f1t[15]_i_9_n_0 ),
        .I5(\u_geo/u_geo_clip/w_add_in_a [10]),
        .O(\r_f1t[2]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[2]_i_6 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [6]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [14]),
        .I3(\r_f1t[11]_i_5_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m0_out [2]),
        .I5(\u_geo/u_geo_matrix/w_m0_out [10]),
        .O(\r_f1t[2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[2]_i_6__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [6]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [14]),
        .I3(\r_f1t[11]_i_5__0_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m2_out [2]),
        .I5(\u_geo/u_geo_matrix/w_m2_out [10]),
        .O(\r_f1t[2]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[2]_i_6__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [6]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [14]),
        .I3(\r_f1t[11]_i_5__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add01_out [2]),
        .I5(\u_geo/u_geo_matrix/w_add01_out [10]),
        .O(\r_f1t[2]_i_6__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[3]_i_1 
       (.I0(\r_f1t[4]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[3]_i_2_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[3]_i_3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[3]_i_1__0 
       (.I0(\r_f1t[4]_i_2__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\r_f1t[3]_i_2__0_n_0 ),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[3]_i_3__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[3]_i_1__1 
       (.I0(\r_f1t[4]_i_2__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[3]_i_2__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[3]_i_3__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[3]_i_1__2 
       (.I0(\r_f1t[4]_i_2__2_n_0 ),
        .I1(\r_f1t[15]_i_6__2_n_0 ),
        .I2(\r_f1t[3]_i_2__2_n_0 ),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f1t[15]_i_5_n_0 ),
        .I5(\r_f1t[3]_i_3__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[3]_i_1__3 
       (.I0(\r_f1t[11]_i_2__3_n_0 ),
        .I1(\r_f1t[3]_i_2__3_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[4]_i_2__3_n_0 ),
        .I4(\r_f1t[3]_i_3__3_n_0 ),
        .I5(\r_f1t[13]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[3]_i_2 
       (.I0(\r_f1t[5]_i_4_n_0 ),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[3]_i_4__1_n_0 ),
        .O(\r_f1t[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[3]_i_2__0 
       (.I0(\r_f1t[5]_i_4__0_n_0 ),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[3]_i_4__2_n_0 ),
        .O(\r_f1t[3]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[3]_i_2__1 
       (.I0(\r_f1t[5]_i_4__1_n_0 ),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[3]_i_4__3_n_0 ),
        .O(\r_f1t[3]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[3]_i_2__2 
       (.I0(\r_f1t[5]_i_4__2_n_0 ),
        .I1(\r_f1t[15]_i_2_n_0 ),
        .I2(\r_f1t[3]_i_4_n_0 ),
        .O(\r_f1t[3]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \r_f1t[3]_i_2__3 
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ),
        .I1(\u_geo/u_geo_viewport/sel0 [3]),
        .I2(\u_geo/u_geo_viewport/sel0 [2]),
        .O(\r_f1t[3]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFFFB8B80000B8)) 
    \r_f1t[3]_i_3 
       (.I0(\r_f1t[5]_i_6_n_0 ),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[3]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [16]),
        .I4(\u_geo/u_geo_matrix/w_m1_out [16]),
        .I5(\r_f1t[4]_i_5_n_0 ),
        .O(\r_f1t[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFFFB8B80000B8)) 
    \r_f1t[3]_i_3__0 
       (.I0(\r_f1t[5]_i_6__0_n_0 ),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[3]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [16]),
        .I4(\u_geo/u_geo_matrix/w_m3_out [16]),
        .I5(\r_f1t[4]_i_5__0_n_0 ),
        .O(\r_f1t[3]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFFFB8B80000B8)) 
    \r_f1t[3]_i_3__1 
       (.I0(\r_f1t[5]_i_6__1_n_0 ),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[3]_i_5__2_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [16]),
        .I4(\u_geo/u_geo_matrix/w_add23_out [16]),
        .I5(\r_f1t[4]_i_5__1_n_0 ),
        .O(\r_f1t[3]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[3]_i_3__2 
       (.I0(\r_f1t[5]_i_5__2_n_0 ),
        .I1(\r_f1t[3]_i_5_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[6]_i_6__2_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[4]_i_5__2_n_0 ),
        .O(\r_f1t[3]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[3]_i_3__3 
       (.I0(\r_f1t[5]_i_3__0_n_0 ),
        .I1(\u_geo/u_geo_viewport/sel0 [1]),
        .I2(\r_f1t[3]_i_4__0_n_0 ),
        .O(\r_f1t[3]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3030505F3F3F505F)) 
    \r_f1t[3]_i_4 
       (.I0(\r_f0[7]_i_2_n_0 ),
        .I1(\r_f0[15]_i_3__2_n_0 ),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\r_f0[3]_i_2_n_0 ),
        .I4(\r_f1t[15]_i_9_n_0 ),
        .I5(\r_f0[11]_i_2_n_0 ),
        .O(\r_f1t[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \r_f1t[3]_i_4__0 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [3]),
        .I1(\u_geo/u_geo_viewport/w_fadd_a [11]),
        .I2(\u_geo/u_geo_viewport/sel0 [2]),
        .I3(\u_geo/u_geo_viewport/w_fadd_a [15]),
        .I4(\u_geo/u_geo_viewport/sel0 [3]),
        .I5(\u_geo/u_geo_viewport/w_fadd_a [7]),
        .O(\r_f1t[3]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[3]_i_4__1 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [7]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [15]),
        .I3(\r_f1t[11]_i_5_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m1_out [3]),
        .I5(\u_geo/u_geo_matrix/w_m1_out [11]),
        .O(\r_f1t[3]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[3]_i_4__2 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [7]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [15]),
        .I3(\r_f1t[11]_i_5__0_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m3_out [3]),
        .I5(\u_geo/u_geo_matrix/w_m3_out [11]),
        .O(\r_f1t[3]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[3]_i_4__3 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [7]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [15]),
        .I3(\r_f1t[11]_i_5__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add23_out [3]),
        .I5(\u_geo/u_geo_matrix/w_add23_out [11]),
        .O(\r_f1t[3]_i_4__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3030505F3F3F505F)) 
    \r_f1t[3]_i_5 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [7]),
        .I1(\u_geo/u_geo_clip/w_add_in_a [15]),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\u_geo/u_geo_clip/w_add_in_a [3]),
        .I4(\r_f1t[15]_i_9_n_0 ),
        .I5(\u_geo/u_geo_clip/w_add_in_a [11]),
        .O(\r_f1t[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[3]_i_5__0 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [7]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [15]),
        .I3(\r_f1t[11]_i_5_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m0_out [3]),
        .I5(\u_geo/u_geo_matrix/w_m0_out [11]),
        .O(\r_f1t[3]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[3]_i_5__1 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [7]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [15]),
        .I3(\r_f1t[11]_i_5__0_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m2_out [3]),
        .I5(\u_geo/u_geo_matrix/w_m2_out [11]),
        .O(\r_f1t[3]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1B001B551BAA1BFF)) 
    \r_f1t[3]_i_5__2 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [7]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [15]),
        .I3(\r_f1t[11]_i_5__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add01_out [3]),
        .I5(\u_geo/u_geo_matrix/w_add01_out [11]),
        .O(\r_f1t[3]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[4]_i_1 
       (.I0(\r_f1t[5]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[4]_i_2_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[4]_i_3__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[4]_i_1__0 
       (.I0(\r_f1t[5]_i_2__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\r_f1t[4]_i_2__0_n_0 ),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[4]_i_3__2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[4]_i_1__1 
       (.I0(\r_f1t[5]_i_2__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[4]_i_2__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[4]_i_3__3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[4]_i_1__2 
       (.I0(\r_f1t[5]_i_2__2_n_0 ),
        .I1(\r_f1t[15]_i_6__2_n_0 ),
        .I2(\r_f1t[4]_i_2__2_n_0 ),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f1t[15]_i_5_n_0 ),
        .I5(\r_f1t[4]_i_3_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[4]_i_1__3 
       (.I0(\r_f1t[12]_i_2__3_n_0 ),
        .I1(\r_f1t[7]_i_2__3_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[5]_i_2__3_n_0 ),
        .I4(\r_f1t[4]_i_2__3_n_0 ),
        .I5(\r_f1t[13]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[4]_i_2 
       (.I0(\r_f1t[6]_i_4_n_0 ),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[4]_i_4_n_0 ),
        .O(\r_f1t[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[4]_i_2__0 
       (.I0(\r_f1t[6]_i_4__0_n_0 ),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[4]_i_4__0_n_0 ),
        .O(\r_f1t[4]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[4]_i_2__1 
       (.I0(\r_f1t[6]_i_4__1_n_0 ),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[4]_i_4__1_n_0 ),
        .O(\r_f1t[4]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[4]_i_2__2 
       (.I0(\r_f1t[6]_i_5__2_n_0 ),
        .I1(\r_f1t[15]_i_2_n_0 ),
        .I2(\r_f1t[4]_i_4__2_n_0 ),
        .O(\r_f1t[4]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[4]_i_2__3 
       (.I0(\r_f1t[6]_i_3__3_n_0 ),
        .I1(\u_geo/u_geo_viewport/sel0 [1]),
        .I2(\r_f1t[4]_i_3__0_n_0 ),
        .O(\r_f1t[4]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[4]_i_3 
       (.I0(\r_f1t[6]_i_6__2_n_0 ),
        .I1(\r_f1t[4]_i_5__2_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[7]_i_5__2_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[5]_i_5__2_n_0 ),
        .O(\r_f1t[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE200FFFFE200E200)) 
    \r_f1t[4]_i_3__0 
       (.I0(\u_geo/w_vy_pdiv [8]),
        .I1(\r_f0[15]_i_2_n_0 ),
        .I2(\u_geo/w_vx_pdiv [8]),
        .I3(\r_f1t[11]_i_5__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/sel0 [2]),
        .I5(\r_f1t[0]_i_4__0_n_0 ),
        .O(\r_f1t[4]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00B8B8B8B8FF00)) 
    \r_f1t[4]_i_3__1 
       (.I0(\r_f1t[5]_i_5_n_0 ),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[5]_i_6_n_0 ),
        .I3(\r_f1t[4]_i_5_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m0_out [16]),
        .I5(\u_geo/u_geo_matrix/w_m1_out [16]),
        .O(\r_f1t[4]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00B8B8B8B8FF00)) 
    \r_f1t[4]_i_3__2 
       (.I0(\r_f1t[5]_i_5__0_n_0 ),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[5]_i_6__0_n_0 ),
        .I3(\r_f1t[4]_i_5__0_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m2_out [16]),
        .I5(\u_geo/u_geo_matrix/w_m3_out [16]),
        .O(\r_f1t[4]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00B8B8B8B8FF00)) 
    \r_f1t[4]_i_3__3 
       (.I0(\r_f1t[5]_i_5__1_n_0 ),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[5]_i_6__1_n_0 ),
        .I3(\r_f1t[4]_i_5__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add01_out [16]),
        .I5(\u_geo/u_geo_matrix/w_add23_out [16]),
        .O(\r_f1t[4]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[4]_i_4 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [8]),
        .I1(\r_f1t[11]_i_5_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [4]),
        .I3(\r_f1t[11]_i_4__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m1_out [12]),
        .O(\r_f1t[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[4]_i_4__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [8]),
        .I1(\r_f1t[11]_i_5__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [4]),
        .I3(\r_f1t[11]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m3_out [12]),
        .O(\r_f1t[4]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[4]_i_4__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [8]),
        .I1(\r_f1t[11]_i_5__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [4]),
        .I3(\r_f1t[11]_i_4__3_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add23_out [12]),
        .O(\r_f1t[4]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[4]_i_4__2 
       (.I0(\r_f0[8]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_8__2_n_0 ),
        .I2(\r_f0[4]_i_2_n_0 ),
        .I3(\r_f1t[15]_i_9_n_0 ),
        .I4(\r_f0[12]_i_2_n_0 ),
        .O(\r_f1t[4]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[4]_i_5 
       (.I0(\r_f1t[6]_i_6_n_0 ),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[2]_i_5_n_0 ),
        .O(\r_f1t[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[4]_i_5__0 
       (.I0(\r_f1t[6]_i_6__0_n_0 ),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[2]_i_5__0_n_0 ),
        .O(\r_f1t[4]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[4]_i_5__1 
       (.I0(\r_f1t[6]_i_6__1_n_0 ),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[2]_i_5__1_n_0 ),
        .O(\r_f1t[4]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[4]_i_5__2 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [8]),
        .I1(\r_f1t[15]_i_8__2_n_0 ),
        .I2(\u_geo/u_geo_clip/w_add_in_a [4]),
        .I3(\r_f1t[15]_i_9_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [12]),
        .O(\r_f1t[4]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[5]_i_1 
       (.I0(\r_f1t[6]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[5]_i_2_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[5]_i_3__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[5]_i_1__0 
       (.I0(\r_f1t[6]_i_2__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\r_f1t[5]_i_2__0_n_0 ),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[5]_i_3__2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[5]_i_1__1 
       (.I0(\r_f1t[6]_i_2__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[5]_i_2__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[5]_i_3__3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[5]_i_1__2 
       (.I0(\r_f1t[6]_i_3__2_n_0 ),
        .I1(\r_f1t[15]_i_6__2_n_0 ),
        .I2(\r_f1t[5]_i_2__2_n_0 ),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f1t[15]_i_5_n_0 ),
        .I5(\r_f1t[5]_i_3_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[5]_i_1__3 
       (.I0(\r_f1t[13]_i_2__3_n_0 ),
        .I1(\r_f1t[7]_i_2__3_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[6]_i_2__3_n_0 ),
        .I4(\r_f1t[5]_i_2__3_n_0 ),
        .I5(\r_f1t[13]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[5]_i_2 
       (.I0(\r_f1t[7]_i_4_n_0 ),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[5]_i_4_n_0 ),
        .O(\r_f1t[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[5]_i_2__0 
       (.I0(\r_f1t[7]_i_4__0_n_0 ),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[5]_i_4__0_n_0 ),
        .O(\r_f1t[5]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[5]_i_2__1 
       (.I0(\r_f1t[7]_i_4__1_n_0 ),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[5]_i_4__1_n_0 ),
        .O(\r_f1t[5]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[5]_i_2__2 
       (.I0(\r_f1t[7]_i_4__2_n_0 ),
        .I1(\r_f1t[15]_i_2_n_0 ),
        .I2(\r_f1t[5]_i_4__2_n_0 ),
        .O(\r_f1t[5]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[5]_i_2__3 
       (.I0(\r_f1t[7]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_viewport/sel0 [1]),
        .I2(\r_f1t[5]_i_3__0_n_0 ),
        .O(\r_f1t[5]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[5]_i_3 
       (.I0(\r_f1t[7]_i_5__2_n_0 ),
        .I1(\r_f1t[5]_i_5__2_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[8]_i_7__2_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[6]_i_6__2_n_0 ),
        .O(\r_f1t[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE200FFFFE200E200)) 
    \r_f1t[5]_i_3__0 
       (.I0(\u_geo/w_vy_pdiv [9]),
        .I1(\r_f0[15]_i_2_n_0 ),
        .I2(\u_geo/w_vx_pdiv [9]),
        .I3(\r_f1t[11]_i_5__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/sel0 [2]),
        .I5(\r_f1t[1]_i_4__0_n_0 ),
        .O(\r_f1t[5]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFFFB8B80000B8)) 
    \r_f1t[5]_i_3__1 
       (.I0(\r_f1t[5]_i_5_n_0 ),
        .I1(\r_f1t[15]_i_4_n_0 ),
        .I2(\r_f1t[5]_i_6_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [16]),
        .I4(\u_geo/u_geo_matrix/w_m1_out [16]),
        .I5(\r_f1t[6]_i_5_n_0 ),
        .O(\r_f1t[5]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFFFB8B80000B8)) 
    \r_f1t[5]_i_3__2 
       (.I0(\r_f1t[5]_i_5__0_n_0 ),
        .I1(\r_f1t[15]_i_4__0_n_0 ),
        .I2(\r_f1t[5]_i_6__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [16]),
        .I4(\u_geo/u_geo_matrix/w_m3_out [16]),
        .I5(\r_f1t[6]_i_5__0_n_0 ),
        .O(\r_f1t[5]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFFFB8B80000B8)) 
    \r_f1t[5]_i_3__3 
       (.I0(\r_f1t[5]_i_5__1_n_0 ),
        .I1(\r_f1t[15]_i_4__1_n_0 ),
        .I2(\r_f1t[5]_i_6__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [16]),
        .I4(\u_geo/u_geo_matrix/w_add23_out [16]),
        .I5(\r_f1t[6]_i_5__1_n_0 ),
        .O(\r_f1t[5]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[5]_i_4 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [9]),
        .I1(\r_f1t[11]_i_5_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [5]),
        .I3(\r_f1t[11]_i_4__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m1_out [13]),
        .O(\r_f1t[5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[5]_i_4__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [9]),
        .I1(\r_f1t[11]_i_5__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [5]),
        .I3(\r_f1t[11]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m3_out [13]),
        .O(\r_f1t[5]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[5]_i_4__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [9]),
        .I1(\r_f1t[11]_i_5__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [5]),
        .I3(\r_f1t[11]_i_4__3_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add23_out [13]),
        .O(\r_f1t[5]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[5]_i_4__2 
       (.I0(\r_f0[9]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_8__2_n_0 ),
        .I2(\r_f0[5]_i_2_n_0 ),
        .I3(\r_f1t[15]_i_9_n_0 ),
        .I4(\r_f0[13]_i_2_n_0 ),
        .O(\r_f1t[5]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[5]_i_5 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [11]),
        .I1(\r_f1t[11]_i_5_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m0_out [7]),
        .I3(\r_f1t[11]_i_4__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m0_out [15]),
        .O(\r_f1t[5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[5]_i_5__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [11]),
        .I1(\r_f1t[11]_i_5__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m2_out [7]),
        .I3(\r_f1t[11]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m2_out [15]),
        .O(\r_f1t[5]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[5]_i_5__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [11]),
        .I1(\r_f1t[11]_i_5__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add01_out [7]),
        .I3(\r_f1t[11]_i_4__3_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add01_out [15]),
        .O(\r_f1t[5]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[5]_i_5__2 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [9]),
        .I1(\r_f1t[15]_i_8__2_n_0 ),
        .I2(\u_geo/u_geo_clip/w_add_in_a [5]),
        .I3(\r_f1t[15]_i_9_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [13]),
        .O(\r_f1t[5]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[5]_i_6 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [9]),
        .I1(\r_f1t[11]_i_5_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m0_out [5]),
        .I3(\r_f1t[11]_i_4__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m0_out [13]),
        .O(\r_f1t[5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[5]_i_6__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [9]),
        .I1(\r_f1t[11]_i_5__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m2_out [5]),
        .I3(\r_f1t[11]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m2_out [13]),
        .O(\r_f1t[5]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[5]_i_6__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [9]),
        .I1(\r_f1t[11]_i_5__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add01_out [5]),
        .I3(\r_f1t[11]_i_4__3_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add01_out [13]),
        .O(\r_f1t[5]_i_6__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[6]_i_1 
       (.I0(\r_f1t[7]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[6]_i_2_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[6]_i_3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[6]_i_1__0 
       (.I0(\r_f1t[7]_i_2__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\r_f1t[6]_i_2__0_n_0 ),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[6]_i_3__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[6]_i_1__1 
       (.I0(\r_f1t[7]_i_2__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[6]_i_2__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[6]_i_3__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[6]_i_1__2 
       (.I0(\r_f1t[6]_i_2__2_n_0 ),
        .I1(\r_f1t[15]_i_6__2_n_0 ),
        .I2(\r_f1t[6]_i_3__2_n_0 ),
        .I3(\r_f0[15]_i_2__3_n_0 ),
        .I4(\r_f1t[15]_i_5_n_0 ),
        .I5(\r_f1t[6]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[6]_i_1__3 
       (.I0(\r_f1t[14]_i_2__3_n_0 ),
        .I1(\r_f1t[7]_i_2__3_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[7]_i_3__3_n_0 ),
        .I4(\r_f1t[6]_i_2__3_n_0 ),
        .I5(\r_f1t[13]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[6]_i_2 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [8]),
        .I2(\r_f1t[11]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m1_out [12]),
        .I4(\r_f1t[15]_i_4_n_0 ),
        .I5(\r_f1t[6]_i_4_n_0 ),
        .O(\r_f1t[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[6]_i_2__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [8]),
        .I2(\r_f1t[11]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m3_out [12]),
        .I4(\r_f1t[15]_i_4__0_n_0 ),
        .I5(\r_f1t[6]_i_4__0_n_0 ),
        .O(\r_f1t[6]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[6]_i_2__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [8]),
        .I2(\r_f1t[11]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add23_out [12]),
        .I4(\r_f1t[15]_i_4__1_n_0 ),
        .I5(\r_f1t[6]_i_4__1_n_0 ),
        .O(\r_f1t[6]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[6]_i_2__2 
       (.I0(\r_f1t[9]_i_5_n_0 ),
        .I1(\r_f1t[15]_i_2_n_0 ),
        .I2(\r_f1t[7]_i_4__2_n_0 ),
        .O(\r_f1t[6]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF888FFFFF8880000)) 
    \r_f1t[6]_i_2__3 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [12]),
        .I1(\r_f1t[11]_i_5__2_n_0 ),
        .I2(\u_geo/u_geo_viewport/w_fadd_a [8]),
        .I3(\r_f1t[15]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/sel0 [1]),
        .I5(\r_f1t[6]_i_3__3_n_0 ),
        .O(\r_f1t[6]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \r_f1t[6]_i_3 
       (.I0(\r_f1t[6]_i_5_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [16]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [16]),
        .I3(\r_f1t[7]_i_5_n_0 ),
        .O(\r_f1t[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \r_f1t[6]_i_3__0 
       (.I0(\r_f1t[6]_i_5__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [16]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [16]),
        .I3(\r_f1t[7]_i_5__0_n_0 ),
        .O(\r_f1t[6]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \r_f1t[6]_i_3__1 
       (.I0(\r_f1t[6]_i_5__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [16]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [16]),
        .I3(\r_f1t[7]_i_5__1_n_0 ),
        .O(\r_f1t[6]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_f1t[6]_i_3__2 
       (.I0(\r_f1t[8]_i_5__2_n_0 ),
        .I1(\r_f1t[15]_i_2_n_0 ),
        .I2(\r_f1t[6]_i_5__2_n_0 ),
        .O(\r_f1t[6]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE200FFFFE200E200)) 
    \r_f1t[6]_i_3__3 
       (.I0(\u_geo/w_vy_pdiv [10]),
        .I1(\r_f0[15]_i_2_n_0 ),
        .I2(\u_geo/w_vx_pdiv [10]),
        .I3(\r_f1t[11]_i_5__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/sel0 [2]),
        .I5(\r_f1t[6]_i_4__3_n_0 ),
        .O(\r_f1t[6]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[6]_i_4 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [10]),
        .I1(\r_f1t[11]_i_5_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [6]),
        .I3(\r_f1t[11]_i_4__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m1_out [14]),
        .O(\r_f1t[6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[6]_i_4__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [10]),
        .I1(\r_f1t[11]_i_5__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [6]),
        .I3(\r_f1t[11]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m3_out [14]),
        .O(\r_f1t[6]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[6]_i_4__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [10]),
        .I1(\r_f1t[11]_i_5__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [6]),
        .I3(\r_f1t[11]_i_4__3_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add23_out [14]),
        .O(\r_f1t[6]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[6]_i_4__2 
       (.I0(\r_f1t[8]_i_7__2_n_0 ),
        .I1(\r_f1t[6]_i_6__2_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[9]_i_4__2_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[7]_i_5__2_n_0 ),
        .O(\r_f1t[6]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFAFA0C0C0AFA0)) 
    \r_f1t[6]_i_4__3 
       (.I0(\u_geo/w_vy_pdiv [14]),
        .I1(\u_geo/w_vx_pdiv [14]),
        .I2(\u_geo/u_geo_viewport/sel0 [3]),
        .I3(\u_geo/w_vy_pdiv [6]),
        .I4(\r_f0[15]_i_2_n_0 ),
        .I5(\u_geo/w_vx_pdiv [6]),
        .O(\r_f1t[6]_i_4__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[6]_i_5 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [8]),
        .I2(\r_f1t[11]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [12]),
        .I4(\r_f1t[15]_i_4_n_0 ),
        .I5(\r_f1t[6]_i_6_n_0 ),
        .O(\r_f1t[6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[6]_i_5__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [8]),
        .I2(\r_f1t[11]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [12]),
        .I4(\r_f1t[15]_i_4__0_n_0 ),
        .I5(\r_f1t[6]_i_6__0_n_0 ),
        .O(\r_f1t[6]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[6]_i_5__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [8]),
        .I2(\r_f1t[11]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [12]),
        .I4(\r_f1t[15]_i_4__1_n_0 ),
        .I5(\r_f1t[6]_i_6__1_n_0 ),
        .O(\r_f1t[6]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[6]_i_5__2 
       (.I0(\r_f0[10]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_8__2_n_0 ),
        .I2(\r_f0[6]_i_2_n_0 ),
        .I3(\r_f1t[15]_i_9_n_0 ),
        .I4(\r_f0[14]_i_2_n_0 ),
        .O(\r_f1t[6]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[6]_i_6 
       (.I0(\u_geo/u_geo_matrix/w_m0_out [10]),
        .I1(\r_f1t[11]_i_5_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m0_out [6]),
        .I3(\r_f1t[11]_i_4__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m0_out [14]),
        .O(\r_f1t[6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[6]_i_6__0 
       (.I0(\u_geo/u_geo_matrix/w_m2_out [10]),
        .I1(\r_f1t[11]_i_5__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m2_out [6]),
        .I3(\r_f1t[11]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m2_out [14]),
        .O(\r_f1t[6]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[6]_i_6__1 
       (.I0(\u_geo/u_geo_matrix/w_add01_out [10]),
        .I1(\r_f1t[11]_i_5__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add01_out [6]),
        .I3(\r_f1t[11]_i_4__3_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add01_out [14]),
        .O(\r_f1t[6]_i_6__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[6]_i_6__2 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [10]),
        .I1(\r_f1t[15]_i_8__2_n_0 ),
        .I2(\u_geo/u_geo_clip/w_add_in_a [6]),
        .I3(\r_f1t[15]_i_9_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [14]),
        .O(\r_f1t[6]_i_6__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[7]_i_1 
       (.I0(\r_f1t[8]_i_3_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[7]_i_2_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[7]_i_3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[7]_i_1__0 
       (.I0(\r_f1t[8]_i_3__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\r_f1t[7]_i_2__0_n_0 ),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[7]_i_3__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[7]_i_1__1 
       (.I0(\r_f1t[8]_i_3__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[7]_i_2__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[7]_i_3__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4070)) 
    \r_f1t[7]_i_1__2 
       (.I0(\r_f1t[7]_i_2__2_n_0 ),
        .I1(\r_f0[15]_i_2__3_n_0 ),
        .I2(\r_f1t[15]_i_5_n_0 ),
        .I3(\r_f1t[7]_i_3__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[7]_i_1__3 
       (.I0(\r_f1t[11]_i_2__3_n_0 ),
        .I1(\r_f1t[7]_i_2__3_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[8]_i_2__3_n_0 ),
        .I4(\r_f1t[7]_i_3__3_n_0 ),
        .I5(\r_f1t[13]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[7]_i_2 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [9]),
        .I2(\r_f1t[11]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m1_out [13]),
        .I4(\r_f1t[15]_i_4_n_0 ),
        .I5(\r_f1t[7]_i_4_n_0 ),
        .O(\r_f1t[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[7]_i_2__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [9]),
        .I2(\r_f1t[11]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m3_out [13]),
        .I4(\r_f1t[15]_i_4__0_n_0 ),
        .I5(\r_f1t[7]_i_4__0_n_0 ),
        .O(\r_f1t[7]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[7]_i_2__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [9]),
        .I2(\r_f1t[11]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add23_out [13]),
        .I4(\r_f1t[15]_i_4__1_n_0 ),
        .I5(\r_f1t[7]_i_4__1_n_0 ),
        .O(\r_f1t[7]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[7]_i_2__2 
       (.I0(\r_f1t[9]_i_5_n_0 ),
        .I1(\r_f1t[7]_i_4__2_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[8]_i_4__2_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[8]_i_5__2_n_0 ),
        .O(\r_f1t[7]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \r_f1t[7]_i_2__3 
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ),
        .I1(\u_geo/u_geo_viewport/sel0 [3]),
        .I2(\u_geo/u_geo_viewport/sel0 [2]),
        .O(\r_f1t[7]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \r_f1t[7]_i_3 
       (.I0(\r_f1t[7]_i_5_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [16]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [16]),
        .I3(\r_f1t[8]_i_7_n_0 ),
        .O(\r_f1t[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \r_f1t[7]_i_3__0 
       (.I0(\r_f1t[7]_i_5__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [16]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [16]),
        .I3(\r_f1t[8]_i_7__0_n_0 ),
        .O(\r_f1t[7]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \r_f1t[7]_i_3__1 
       (.I0(\r_f1t[7]_i_5__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [16]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [16]),
        .I3(\r_f1t[8]_i_7__1_n_0 ),
        .O(\r_f1t[7]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[7]_i_3__2 
       (.I0(\r_f1t[9]_i_4__2_n_0 ),
        .I1(\r_f1t[7]_i_5__2_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[8]_i_6__2_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[8]_i_7__2_n_0 ),
        .O(\r_f1t[7]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF888FFFFF8880000)) 
    \r_f1t[7]_i_3__3 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [13]),
        .I1(\r_f1t[11]_i_5__2_n_0 ),
        .I2(\u_geo/u_geo_viewport/w_fadd_a [9]),
        .I3(\r_f1t[15]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/sel0 [1]),
        .I5(\r_f1t[7]_i_4__3_n_0 ),
        .O(\r_f1t[7]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[7]_i_4 
       (.I0(\u_geo/u_geo_matrix/w_m1_out [11]),
        .I1(\r_f1t[11]_i_5_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [7]),
        .I3(\r_f1t[11]_i_4__1_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m1_out [15]),
        .O(\r_f1t[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[7]_i_4__0 
       (.I0(\u_geo/u_geo_matrix/w_m3_out [11]),
        .I1(\r_f1t[11]_i_5__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [7]),
        .I3(\r_f1t[11]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_m3_out [15]),
        .O(\r_f1t[7]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[7]_i_4__1 
       (.I0(\u_geo/u_geo_matrix/w_add23_out [11]),
        .I1(\r_f1t[11]_i_5__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [7]),
        .I3(\r_f1t[11]_i_4__3_n_0 ),
        .I4(\u_geo/u_geo_matrix/w_add23_out [15]),
        .O(\r_f1t[7]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[7]_i_4__2 
       (.I0(\r_f0[11]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_8__2_n_0 ),
        .I2(\r_f0[7]_i_2_n_0 ),
        .I3(\r_f1t[15]_i_9_n_0 ),
        .I4(\r_f0[15]_i_3__2_n_0 ),
        .O(\r_f1t[7]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE200FFFFE200E200)) 
    \r_f1t[7]_i_4__3 
       (.I0(\u_geo/w_vy_pdiv [11]),
        .I1(\r_f0[15]_i_2_n_0 ),
        .I2(\u_geo/w_vx_pdiv [11]),
        .I3(\r_f1t[11]_i_5__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/sel0 [2]),
        .I5(\r_f1t[7]_i_5__3_n_0 ),
        .O(\r_f1t[7]_i_4__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[7]_i_5 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [9]),
        .I2(\r_f1t[11]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [13]),
        .I4(\r_f1t[15]_i_4_n_0 ),
        .I5(\r_f1t[5]_i_5_n_0 ),
        .O(\r_f1t[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[7]_i_5__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [9]),
        .I2(\r_f1t[11]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [13]),
        .I4(\r_f1t[15]_i_4__0_n_0 ),
        .I5(\r_f1t[5]_i_5__0_n_0 ),
        .O(\r_f1t[7]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[7]_i_5__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [9]),
        .I2(\r_f1t[11]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [13]),
        .I4(\r_f1t[15]_i_4__1_n_0 ),
        .I5(\r_f1t[5]_i_5__1_n_0 ),
        .O(\r_f1t[7]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCC47FF47)) 
    \r_f1t[7]_i_5__2 
       (.I0(\u_geo/u_geo_clip/w_add_in_a [11]),
        .I1(\r_f1t[15]_i_8__2_n_0 ),
        .I2(\u_geo/u_geo_clip/w_add_in_a [7]),
        .I3(\r_f1t[15]_i_9_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [15]),
        .O(\r_f1t[7]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFCFAFA0C0C0AFA0)) 
    \r_f1t[7]_i_5__3 
       (.I0(\u_geo/w_vy_pdiv [15]),
        .I1(\u_geo/w_vx_pdiv [15]),
        .I2(\u_geo/u_geo_viewport/sel0 [3]),
        .I3(\u_geo/w_vy_pdiv [7]),
        .I4(\r_f0[15]_i_2_n_0 ),
        .I5(\u_geo/w_vx_pdiv [7]),
        .O(\r_f1t[7]_i_5__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[8]_i_1 
       (.I0(\r_f1t[8]_i_2_n_0 ),
        .I1(\r_f1t[15]_i_5__0_n_0 ),
        .I2(\r_f1t[8]_i_3_n_0 ),
        .I3(\r_f0[15]_i_2__0_n_0 ),
        .I4(\r_f1t[15]_i_6_n_0 ),
        .I5(\r_f1t[8]_i_4_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[8]_i_1__0 
       (.I0(\r_f1t[8]_i_2__0_n_0 ),
        .I1(\r_f1t[15]_i_5__1_n_0 ),
        .I2(\r_f1t[8]_i_3__0_n_0 ),
        .I3(\r_f0[15]_i_2__1_n_0 ),
        .I4(\r_f1t[15]_i_6__0_n_0 ),
        .I5(\r_f1t[8]_i_4__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D0000001DFF0000)) 
    \r_f1t[8]_i_1__1 
       (.I0(\r_f1t[8]_i_2__1_n_0 ),
        .I1(\r_f1t[15]_i_5__2_n_0 ),
        .I2(\r_f1t[8]_i_3__1_n_0 ),
        .I3(\r_f0[15]_i_2__2_n_0 ),
        .I4(\r_f1t[15]_i_6__1_n_0 ),
        .I5(\r_f1t[8]_i_4__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4070)) 
    \r_f1t[8]_i_1__2 
       (.I0(\r_f1t[8]_i_2__2_n_0 ),
        .I1(\r_f0[15]_i_2__3_n_0 ),
        .I2(\r_f1t[15]_i_5_n_0 ),
        .I3(\r_f1t[8]_i_3__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[8]_i_1__3 
       (.I0(\r_f1t[12]_i_2__3_n_0 ),
        .I1(\r_f1t[11]_i_3__2_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[9]_i_2__3_n_0 ),
        .I4(\r_f1t[8]_i_2__3_n_0 ),
        .I5(\r_f1t[13]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[8]_i_2 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [11]),
        .I2(\r_f1t[11]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m1_out [15]),
        .I4(\r_f1t[15]_i_4_n_0 ),
        .I5(\r_f1t[8]_i_5_n_0 ),
        .O(\r_f1t[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[8]_i_2__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [11]),
        .I2(\r_f1t[11]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m3_out [15]),
        .I4(\r_f1t[15]_i_4__0_n_0 ),
        .I5(\r_f1t[8]_i_5__0_n_0 ),
        .O(\r_f1t[8]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[8]_i_2__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [11]),
        .I2(\r_f1t[11]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add23_out [15]),
        .I4(\r_f1t[15]_i_4__1_n_0 ),
        .I5(\r_f1t[8]_i_5__1_n_0 ),
        .O(\r_f1t[8]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[8]_i_2__2 
       (.I0(\r_f1t[8]_i_4__2_n_0 ),
        .I1(\r_f1t[8]_i_5__2_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[11]_i_4_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[9]_i_5_n_0 ),
        .O(\r_f1t[8]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF888FFFFF8880000)) 
    \r_f1t[8]_i_2__3 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [14]),
        .I1(\r_f1t[11]_i_5__2_n_0 ),
        .I2(\u_geo/u_geo_viewport/w_fadd_a [10]),
        .I3(\r_f1t[15]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/sel0 [1]),
        .I5(\r_f1t[8]_i_3__3_n_0 ),
        .O(\r_f1t[8]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[8]_i_3 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [10]),
        .I2(\r_f1t[11]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m1_out [14]),
        .I4(\r_f1t[15]_i_4_n_0 ),
        .I5(\r_f1t[8]_i_6_n_0 ),
        .O(\r_f1t[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[8]_i_3__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [10]),
        .I2(\r_f1t[11]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m3_out [14]),
        .I4(\r_f1t[15]_i_4__0_n_0 ),
        .I5(\r_f1t[8]_i_6__0_n_0 ),
        .O(\r_f1t[8]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[8]_i_3__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [10]),
        .I2(\r_f1t[11]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add23_out [14]),
        .I4(\r_f1t[15]_i_4__1_n_0 ),
        .I5(\r_f1t[8]_i_6__1_n_0 ),
        .O(\r_f1t[8]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[8]_i_3__2 
       (.I0(\r_f1t[8]_i_6__2_n_0 ),
        .I1(\r_f1t[8]_i_7__2_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[11]_i_6__2_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[9]_i_4__2_n_0 ),
        .O(\r_f1t[8]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE200E200E200)) 
    \r_f1t[8]_i_3__3 
       (.I0(\u_geo/w_vy_pdiv [12]),
        .I1(\r_f0[15]_i_2_n_0 ),
        .I2(\u_geo/w_vx_pdiv [12]),
        .I3(\r_f1t[11]_i_5__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/w_fadd_a [8]),
        .I5(\r_f1t[15]_i_4__2_n_0 ),
        .O(\r_f1t[8]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \r_f1t[8]_i_4 
       (.I0(\r_f1t[8]_i_7_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [16]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [16]),
        .I3(\r_f1t[9]_i_3_n_0 ),
        .O(\r_f1t[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \r_f1t[8]_i_4__0 
       (.I0(\r_f1t[8]_i_7__0_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [16]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [16]),
        .I3(\r_f1t[9]_i_3__0_n_0 ),
        .O(\r_f1t[8]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \r_f1t[8]_i_4__1 
       (.I0(\r_f1t[8]_i_7__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [16]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [16]),
        .I3(\r_f1t[9]_i_3__1_n_0 ),
        .O(\r_f1t[8]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[8]_i_4__2 
       (.I0(\r_f1t[15]_i_9_n_0 ),
        .I1(\r_f0[10]_i_2_n_0 ),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\r_f0[14]_i_2_n_0 ),
        .O(\r_f1t[8]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[8]_i_5 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [9]),
        .I2(\r_f1t[11]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m1_out [13]),
        .O(\r_f1t[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[8]_i_5__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [9]),
        .I2(\r_f1t[11]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m3_out [13]),
        .O(\r_f1t[8]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[8]_i_5__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [9]),
        .I2(\r_f1t[11]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add23_out [13]),
        .O(\r_f1t[8]_i_5__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[8]_i_5__2 
       (.I0(\r_f1t[15]_i_9_n_0 ),
        .I1(\r_f0[8]_i_2_n_0 ),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\r_f0[12]_i_2_n_0 ),
        .O(\r_f1t[8]_i_5__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[8]_i_6 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m1_out [8]),
        .I2(\r_f1t[11]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m1_out [12]),
        .O(\r_f1t[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[8]_i_6__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m3_out [8]),
        .I2(\r_f1t[11]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m3_out [12]),
        .O(\r_f1t[8]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[8]_i_6__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add23_out [8]),
        .I2(\r_f1t[11]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add23_out [12]),
        .O(\r_f1t[8]_i_6__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBABABABFBFBFB)) 
    \r_f1t[8]_i_6__2 
       (.I0(\r_f1t[15]_i_9_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [10]),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\u_geo/w_vw_mvp [14]),
        .I4(\u_geo/w_state_clip ),
        .I5(\u_geo/w_vw_clip [14]),
        .O(\r_f1t[8]_i_6__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[8]_i_7 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [10]),
        .I2(\r_f1t[11]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [14]),
        .I4(\r_f1t[15]_i_4_n_0 ),
        .I5(\r_f1t[8]_i_8_n_0 ),
        .O(\r_f1t[8]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[8]_i_7__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [10]),
        .I2(\r_f1t[11]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [14]),
        .I4(\r_f1t[15]_i_4__0_n_0 ),
        .I5(\r_f1t[8]_i_8__0_n_0 ),
        .O(\r_f1t[8]_i_7__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[8]_i_7__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [10]),
        .I2(\r_f1t[11]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [14]),
        .I4(\r_f1t[15]_i_4__1_n_0 ),
        .I5(\r_f1t[8]_i_8__1_n_0 ),
        .O(\r_f1t[8]_i_7__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBABABABFBFBFB)) 
    \r_f1t[8]_i_7__2 
       (.I0(\r_f1t[15]_i_9_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [8]),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\u_geo/w_vw_mvp [12]),
        .I4(\u_geo/w_state_clip ),
        .I5(\u_geo/w_vw_clip [12]),
        .O(\r_f1t[8]_i_7__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[8]_i_8 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [8]),
        .I2(\r_f1t[11]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [12]),
        .O(\r_f1t[8]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[8]_i_8__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [8]),
        .I2(\r_f1t[11]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [12]),
        .O(\r_f1t[8]_i_8__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[8]_i_8__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [8]),
        .I2(\r_f1t[11]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [12]),
        .O(\r_f1t[8]_i_8__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_f1t[9]_i_1 
       (.I0(\r_f1t[15]_i_6_n_0 ),
        .I1(\r_f1t[9]_i_2_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_f1t[9]_i_1__0 
       (.I0(\r_f1t[15]_i_6__0_n_0 ),
        .I1(\r_f1t[9]_i_2__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_f1t[9]_i_1__1 
       (.I0(\r_f1t[15]_i_6__1_n_0 ),
        .I1(\r_f1t[9]_i_2__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888FF8FF888)) 
    \r_f1t[9]_i_1__2 
       (.I0(\r_f1t[13]_i_2__3_n_0 ),
        .I1(\r_f1t[11]_i_3__2_n_0 ),
        .I2(\u_geo/u_geo_viewport/sel0 [0]),
        .I3(\r_f1t[10]_i_2__3_n_0 ),
        .I4(\r_f1t[9]_i_2__3_n_0 ),
        .I5(\r_f1t[13]_i_4__2_n_0 ),
        .O(\u_geo/u_geo_viewport/w_f1t [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[9]_i_2 
       (.I0(\r_f1t[8]_i_2_n_0 ),
        .I1(\r_f1t[10]_i_2_n_0 ),
        .I2(\r_f0[15]_i_2__0_n_0 ),
        .I3(\r_f1t[9]_i_3_n_0 ),
        .I4(\r_f1t[15]_i_5__0_n_0 ),
        .I5(\r_f1t[10]_i_4_n_0 ),
        .O(\r_f1t[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[9]_i_2__0 
       (.I0(\r_f1t[8]_i_2__0_n_0 ),
        .I1(\r_f1t[10]_i_2__0_n_0 ),
        .I2(\r_f0[15]_i_2__1_n_0 ),
        .I3(\r_f1t[9]_i_3__0_n_0 ),
        .I4(\r_f1t[15]_i_5__1_n_0 ),
        .I5(\r_f1t[10]_i_4__0_n_0 ),
        .O(\r_f1t[9]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_f1t[9]_i_2__1 
       (.I0(\r_f1t[8]_i_2__1_n_0 ),
        .I1(\r_f1t[10]_i_2__1_n_0 ),
        .I2(\r_f0[15]_i_2__2_n_0 ),
        .I3(\r_f1t[9]_i_3__1_n_0 ),
        .I4(\r_f1t[15]_i_5__2_n_0 ),
        .I5(\r_f1t[10]_i_4__1_n_0 ),
        .O(\r_f1t[9]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h020202A2A2A202A2)) 
    \r_f1t[9]_i_2__2 
       (.I0(\r_f1t[15]_i_5_n_0 ),
        .I1(\r_f1t[10]_i_3__2_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[9]_i_4__2_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[11]_i_6__2_n_0 ),
        .O(\r_f1t[9]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF888FFFFF8880000)) 
    \r_f1t[9]_i_2__3 
       (.I0(\u_geo/u_geo_viewport/w_fadd_a [15]),
        .I1(\r_f1t[11]_i_5__2_n_0 ),
        .I2(\u_geo/u_geo_viewport/w_fadd_a [11]),
        .I3(\r_f1t[15]_i_4__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/sel0 [1]),
        .I5(\r_f1t[9]_i_3__3_n_0 ),
        .O(\r_f1t[9]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[9]_i_3 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [11]),
        .I2(\r_f1t[11]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [15]),
        .I4(\r_f1t[15]_i_4_n_0 ),
        .I5(\r_f1t[9]_i_4_n_0 ),
        .O(\r_f1t[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[9]_i_3__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [11]),
        .I2(\r_f1t[11]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [15]),
        .I4(\r_f1t[15]_i_4__0_n_0 ),
        .I5(\r_f1t[9]_i_4__0_n_0 ),
        .O(\r_f1t[9]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBFFFFABFB0000)) 
    \r_f1t[9]_i_3__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [11]),
        .I2(\r_f1t[11]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [15]),
        .I4(\r_f1t[15]_i_4__1_n_0 ),
        .I5(\r_f1t[9]_i_4__1_n_0 ),
        .O(\r_f1t[9]_i_3__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h020202A2A2A202A2)) 
    \r_f1t[9]_i_3__2 
       (.I0(\r_f1t[15]_i_5_n_0 ),
        .I1(\r_f1t[10]_i_2__2_n_0 ),
        .I2(\r_f1t[15]_i_6__2_n_0 ),
        .I3(\r_f1t[9]_i_5_n_0 ),
        .I4(\r_f1t[15]_i_2_n_0 ),
        .I5(\r_f1t[11]_i_4_n_0 ),
        .O(\r_f1t[9]_i_3__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFE200E200E200)) 
    \r_f1t[9]_i_3__3 
       (.I0(\u_geo/w_vy_pdiv [13]),
        .I1(\r_f0[15]_i_2_n_0 ),
        .I2(\u_geo/w_vx_pdiv [13]),
        .I3(\r_f1t[11]_i_5__2_n_0 ),
        .I4(\u_geo/u_geo_viewport/w_fadd_a [9]),
        .I5(\r_f1t[15]_i_4__2_n_0 ),
        .O(\r_f1t[9]_i_3__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[9]_i_4 
       (.I0(\r_f1t[11]_i_4__1_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m0_out [9]),
        .I2(\r_f1t[11]_i_5_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m0_out [13]),
        .O(\r_f1t[9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[9]_i_4__0 
       (.I0(\r_f1t[11]_i_4__2_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_m2_out [9]),
        .I2(\r_f1t[11]_i_5__0_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_m2_out [13]),
        .O(\r_f1t[9]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[9]_i_4__1 
       (.I0(\r_f1t[11]_i_4__3_n_0 ),
        .I1(\u_geo/u_geo_matrix/w_add01_out [9]),
        .I2(\r_f1t[11]_i_5__1_n_0 ),
        .I3(\u_geo/u_geo_matrix/w_add01_out [13]),
        .O(\r_f1t[9]_i_4__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABFBABABABFBFBFB)) 
    \r_f1t[9]_i_4__2 
       (.I0(\r_f1t[15]_i_9_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [9]),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\u_geo/w_vw_mvp [13]),
        .I4(\u_geo/w_state_clip ),
        .I5(\u_geo/w_vw_clip [13]),
        .O(\r_f1t[9]_i_4__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFB)) 
    \r_f1t[9]_i_5 
       (.I0(\r_f1t[15]_i_9_n_0 ),
        .I1(\r_f0[9]_i_2_n_0 ),
        .I2(\r_f1t[15]_i_8__2_n_0 ),
        .I3(\r_f0[13]_i_2_n_0 ),
        .O(\r_f1t[9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_f1t_reg[14]_i_1 
       (.I0(\r_f1t[14]_i_2_n_0 ),
        .I1(\r_f1t[14]_i_3_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [14]),
        .S(\r_f0[15]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_f1t_reg[14]_i_1__0 
       (.I0(\r_f1t[14]_i_2__0_n_0 ),
        .I1(\r_f1t[14]_i_3__0_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [14]),
        .S(\r_f0[15]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_f1t_reg[14]_i_1__1 
       (.I0(\r_f1t[14]_i_2__1_n_0 ),
        .I1(\r_f1t[14]_i_3__1_n_0 ),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [14]),
        .S(\r_f0[15]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_f1t_reg[9]_i_1 
       (.I0(\r_f1t[9]_i_2__2_n_0 ),
        .I1(\r_f1t[9]_i_3__2_n_0 ),
        .O(\u_geo/u_geo_clip/w_f1t [9]),
        .S(\r_f0[15]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEEEEE0E)) 
    r_int_i_1
       (.I0(\u_sys/p_21_in [0]),
        .I1(\u_sys/w_int_set ),
        .I2(r_int_i_3_n_0),
        .I3(\r_dma_size[15]_i_2_n_0 ),
        .I4(\r_m10[21]_i_2_n_0 ),
        .I5(rst_i),
        .O(r_int_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    r_int_i_2
       (.I0(\u_geo/r_int_i_4_n_0 ),
        .I1(\u_geo/r_int_i_5_n_0 ),
        .I2(w_dma_start),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .I5(w_sy_flag1_carry_i_10_n_0),
        .O(\u_sys/w_int_set ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    r_int_i_3
       (.I0(s_wb_adr_i[6]),
        .I1(s_wb_adr_i[5]),
        .O(r_int_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF02000000)) 
    r_int_mask_i_1
       (.I0(s_wb_dat_i[8]),
        .I1(\r_m10[21]_i_2_n_0 ),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(r_int_i_3_n_0),
        .I4(s_wb_sel_i[1]),
        .I5(\u_sys/p_21_in [8]),
        .O(r_int_mask_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    r_int_out_i_1
       (.I0(\u_sys/p_21_in [0]),
        .I1(\u_sys/p_21_in [8]),
        .O(r_int_out_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \r_ivw[15]_i_1 
       (.I0(\u_geo/u_geo_persdiv/r_state [1]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .O(r_ivw));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \r_ivw[16]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[16] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [16]),
        .O(\u_geo/u_geo_persdiv/w_b_exp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \r_ivw[17]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[17] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [17]),
        .O(\u_geo/u_geo_persdiv/w_b_exp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \r_ivw[18]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[18] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [18]),
        .O(\u_geo/u_geo_persdiv/w_b_exp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \r_ivw[19]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[19] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [19]),
        .O(\u_geo/u_geo_persdiv/w_b_exp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \r_ivw[20]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[20] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [20]),
        .O(\u_geo/u_geo_persdiv/w_b_exp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    \r_ivw[21]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[21] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [21]),
        .O(\r_ivw[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h51)) 
    \r_lat_cnt[8]_i_1 
       (.I0(rst_i),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/w_en_dma ),
        .O(\u_geo/u_geo_matrix/r_lat_cnt ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \r_m00[15]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[2]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[6]),
        .I4(s_wb_adr_i[5]),
        .I5(s_wb_sel_i[1]),
        .O(r_m00));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFCCCDCCC)) 
    \r_m00[15]_i_2 
       (.I0(\r_m00[20]_i_2_n_0 ),
        .I1(s_wb_dat_i[30]),
        .I2(s_wb_dat_i[29]),
        .I3(s_wb_dat_i[28]),
        .I4(s_wb_dat_i[27]),
        .O(\u_sys/w_f22 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF80FF800000)) 
    \r_m00[16]_i_1 
       (.I0(s_wb_dat_i[27]),
        .I1(s_wb_dat_i[28]),
        .I2(s_wb_dat_i[29]),
        .I3(s_wb_dat_i[30]),
        .I4(\u_sys/p_0_in ),
        .I5(s_wb_dat_i[23]),
        .O(\u_sys/w_f22 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2A80)) 
    \r_m00[17]_i_1 
       (.I0(\r_m00[19]_i_2_n_0 ),
        .I1(s_wb_dat_i[23]),
        .I2(\u_sys/p_0_in ),
        .I3(s_wb_dat_i[24]),
        .O(\u_sys/w_f22 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    \r_m00[18]_i_1 
       (.I0(\r_m00[19]_i_2_n_0 ),
        .I1(s_wb_dat_i[24]),
        .I2(\u_sys/p_0_in ),
        .I3(s_wb_dat_i[23]),
        .I4(s_wb_dat_i[25]),
        .O(\u_sys/w_f22 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7FFF000080000000)) 
    \r_m00[19]_i_1 
       (.I0(s_wb_dat_i[24]),
        .I1(\u_sys/p_0_in ),
        .I2(s_wb_dat_i[23]),
        .I3(s_wb_dat_i[25]),
        .I4(\r_m00[19]_i_2_n_0 ),
        .I5(s_wb_dat_i[26]),
        .O(\u_sys/w_f22 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF80)) 
    \r_m00[19]_i_2 
       (.I0(s_wb_dat_i[27]),
        .I1(s_wb_dat_i[28]),
        .I2(s_wb_dat_i[29]),
        .I3(s_wb_dat_i[30]),
        .O(\r_m00[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0F08F000)) 
    \r_m00[20]_i_1 
       (.I0(s_wb_dat_i[28]),
        .I1(s_wb_dat_i[29]),
        .I2(\r_m00[20]_i_2_n_0 ),
        .I3(s_wb_dat_i[30]),
        .I4(s_wb_dat_i[27]),
        .O(\u_sys/w_f22 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \r_m00[20]_i_2 
       (.I0(s_wb_dat_i[25]),
        .I1(s_wb_dat_i[23]),
        .I2(\u_sys/p_0_in ),
        .I3(s_wb_dat_i[24]),
        .I4(s_wb_dat_i[26]),
        .O(\r_m00[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \r_m00[21]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[2]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[6]),
        .I4(s_wb_adr_i[5]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m00[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \r_m00[21]_i_2 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_stb_i),
        .I2(s_wb_we_i),
        .O(\r_m00[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_m00[3]_i_5 
       (.I0(s_wb_dat_i[8]),
        .I1(s_wb_dat_i[7]),
        .O(\r_m00[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \r_m00[7]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[2]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[6]),
        .I4(s_wb_adr_i[5]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m00[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_m00_reg[11]_i_1 
       (.CI(\r_m00_reg[7]_i_2_n_0 ),
        .CO(r_m00_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_m00_reg[11]_i_1_n_4 ,\r_m00_reg[11]_i_1_n_5 ,\r_m00_reg[11]_i_1_n_6 ,\r_m00_reg[11]_i_1_n_7 }),
        .S(s_wb_dat_i[19:16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_m00_reg[14]_i_1 
       (.CI(r_m00_reg[3]),
        .CO({\u_sys/p_0_in ,\r_m00_reg[14]_i_1_n_1 ,\r_m00_reg[14]_i_1_n_2 ,\r_m00_reg[14]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_m00_reg[14]_i_1_n_4 ,\r_m00_reg[14]_i_1_n_5 ,\r_m00_reg[14]_i_1_n_6 ,\r_m00_reg[14]_i_1_n_7 }),
        .S({\<const1>__0__0 ,s_wb_dat_i[22:20]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_m00_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\r_m00_reg[3]_i_1_n_0 ,\r_m00_reg[3]_i_1_n_1 ,\r_m00_reg[3]_i_1_n_2 ,\r_m00_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,s_wb_dat_i[8]}),
        .O({\r_m00_reg[3]_i_1_n_4 ,\r_m00_reg[3]_i_1_n_5 ,\r_m00_reg[3]_i_1_n_6 ,\r_m00_reg[3]_i_1_n_7 }),
        .S({s_wb_dat_i[11:9],\r_m00[3]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_m00_reg[7]_i_2 
       (.CI(\r_m00_reg[3]_i_1_n_0 ),
        .CO({\r_m00_reg[7]_i_2_n_0 ,\r_m00_reg[7]_i_2_n_1 ,\r_m00_reg[7]_i_2_n_2 ,\r_m00_reg[7]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_m00_reg[7]_i_2_n_4 ,\r_m00_reg[7]_i_2_n_5 ,\r_m00_reg[7]_i_2_n_6 ,\r_m00_reg[7]_i_2_n_7 }),
        .S(s_wb_dat_i[15:12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m01[15]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[1]),
        .O(r_m01));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m01[21]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m01[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m01[7]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m01[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m02[15]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[2]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[1]),
        .O(r_m02));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m02[21]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[2]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m02[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m02[7]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[2]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m02[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m03[15]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[1]),
        .O(r_m03));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m03[21]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m03[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m03[7]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m03[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \r_m10[15]_i_1 
       (.I0(\r_m10[21]_i_2_n_0 ),
        .I1(\r_m10[21]_i_3_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[1]),
        .O(r_m10));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \r_m10[21]_i_1 
       (.I0(\r_m10[21]_i_2_n_0 ),
        .I1(\r_m10[21]_i_3_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m10[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_m10[21]_i_2 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .O(\r_m10[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r_m10[21]_i_3 
       (.I0(s_wb_we_i),
        .I1(s_wb_stb_i),
        .O(\r_m10[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \r_m10[7]_i_1 
       (.I0(\r_m10[21]_i_2_n_0 ),
        .I1(\r_m10[21]_i_3_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m10[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m11[15]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[1]),
        .O(r_m11));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m11[21]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m11[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m11[7]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m11[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m12[15]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[1]),
        .O(r_m12));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m12[21]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m12[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m12[7]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m12[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m13[15]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[5]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[1]),
        .O(r_m13));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m13[21]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[5]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m13[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m13[7]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[5]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m13[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m20[15]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[2]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[1]),
        .O(r_m20));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m20[21]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[2]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m20[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m20[7]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[2]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m20[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m21[15]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[5]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[1]),
        .O(r_m21));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m21[21]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[5]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m21[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m21[7]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[5]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m21[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m22[15]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[5]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[1]),
        .O(r_m22));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m22[21]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[5]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m22[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m22[7]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[5]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m22[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \r_m23[15]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[6]),
        .I4(s_wb_adr_i[5]),
        .I5(s_wb_sel_i[1]),
        .O(r_m23));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \r_m23[21]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[6]),
        .I4(s_wb_adr_i[5]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m23[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \r_m23[7]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[6]),
        .I4(s_wb_adr_i[5]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m23[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \r_m30[15]_i_1 
       (.I0(\r_m10[21]_i_2_n_0 ),
        .I1(\r_m10[21]_i_3_n_0 ),
        .I2(s_wb_adr_i[6]),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[2]),
        .I5(s_wb_sel_i[1]),
        .O(r_m30));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \r_m30[21]_i_1 
       (.I0(\r_m10[21]_i_2_n_0 ),
        .I1(\r_m10[21]_i_3_n_0 ),
        .I2(s_wb_adr_i[6]),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[2]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m30[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \r_m30[7]_i_1 
       (.I0(\r_m10[21]_i_2_n_0 ),
        .I1(\r_m10[21]_i_3_n_0 ),
        .I2(s_wb_adr_i[6]),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[2]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m30[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m31[15]_i_1 
       (.I0(s_wb_adr_i[6]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[1]),
        .O(r_m31));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m31[21]_i_1 
       (.I0(s_wb_adr_i[6]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m31[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m31[7]_i_1 
       (.I0(s_wb_adr_i[6]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m31[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m32[15]_i_1 
       (.I0(s_wb_adr_i[6]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[2]),
        .I5(s_wb_sel_i[1]),
        .O(r_m32));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m32[21]_i_1 
       (.I0(s_wb_adr_i[6]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[2]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m32[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_m32[7]_i_1 
       (.I0(s_wb_adr_i[6]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_top_address[29]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[2]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m32[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m33[15]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[6]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[4]),
        .I5(s_wb_sel_i[1]),
        .O(r_m33));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m33[21]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[6]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[4]),
        .I5(s_wb_sel_i[2]),
        .O(\r_m33[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_m33[7]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[6]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[4]),
        .I5(s_wb_sel_i[0]),
        .O(\r_m33[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[11]_i_1 
       (.CI(\r_mats_reg[7]_i_1_n_0 ),
        .CO({\r_mats_reg[11]_i_1_n_0 ,\r_mats_reg[11]_i_1_n_1 ,\r_mats_reg[11]_i_1_n_2 ,\r_mats_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [11:8]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [11:8]),
        .S({\u_fadd_m01/r_mats ,\u_fadd_m01/r_mats[11]_i_3_n_0 ,\u_fadd_m01/r_mats[11]_i_4_n_0 ,\u_fadd_m01/r_mats[11]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[11]_i_1__0 
       (.CI(\r_mats_reg[7]_i_1__0_n_0 ),
        .CO(r_mats_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [11:8]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [11:8]),
        .S({\u_fadd_m23/r_mats ,\u_fadd_m23/r_mats[11]_i_3_n_0 ,\u_fadd_m23/r_mats[11]_i_4_n_0 ,\u_fadd_m23/r_mats[11]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[11]_i_1__1 
       (.CI(\r_mats_reg[7]_i_1__1_n_0 ),
        .CO({\r_mats_reg[11]_i_1__1_n_0 ,\r_mats_reg[11]_i_1__1_n_1 ,\r_mats_reg[11]_i_1__1_n_2 ,\r_mats_reg[11]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [11:8]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [11:8]),
        .S({\u_fadd_m0123/r_mats ,\u_fadd_m0123/r_mats[11]_i_3_n_0 ,\u_fadd_m0123/r_mats[11]_i_4_n_0 ,\u_fadd_m0123/r_mats[11]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[11]_i_1__2 
       (.CI(\r_mats_reg[7]_i_1__2_n_0 ),
        .CO({\r_mats_reg[11]_i_1__2_n_0 ,\r_mats_reg[11]_i_1__2_n_1 ,\r_mats_reg[11]_i_1__2_n_2 ,\r_mats_reg[11]_i_1__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_clip/r_f0 [11:8]),
        .O(\u_geo/u_geo_clip/w_mats [11:8]),
        .S({\u_fadd/r_mats[11]_i_2_n_0 ,\u_fadd/r_mats[11]_i_3_n_0 ,\u_fadd/r_mats[11]_i_4_n_0 ,\u_fadd/r_mats[11]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[11]_i_1__3 
       (.CI(\r_mats_reg[7]_i_1__3_n_0 ),
        .CO({\r_mats_reg[11]_i_1__3_n_0 ,\r_mats_reg[11]_i_1__3_n_1 ,\r_mats_reg[11]_i_1__3_n_2 ,\r_mats_reg[11]_i_1__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_viewport/r_f0 [11:8]),
        .O(\u_geo/u_geo_viewport/w_mats [11:8]),
        .S({\u_fadd/r_mats ,\u_fadd/r_mats[11]_i_3__0_n_0 ,\u_fadd/r_mats[11]_i_4__0_n_0 ,\u_fadd/r_mats[11]_i_5__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[15]_i_1 
       (.CI(\r_mats_reg[11]_i_1_n_0 ),
        .CO({\r_mats_reg[15]_i_1_n_0 ,\r_mats_reg[15]_i_1_n_1 ,\r_mats_reg[15]_i_1_n_2 ,\r_mats_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [15:12]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [15:12]),
        .S({\u_fadd_m01/r_mats[15]_i_2_n_0 ,\u_fadd_m01/r_mats[15]_i_3_n_0 ,\u_fadd_m01/r_mats[15]_i_4_n_0 ,\u_fadd_m01/r_mats[15]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[15]_i_1__0 
       (.CI(r_mats_reg[3]),
        .CO({\r_mats_reg[15]_i_1__0_n_0 ,\r_mats_reg[15]_i_1__0_n_1 ,\r_mats_reg[15]_i_1__0_n_2 ,\r_mats_reg[15]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [15:12]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [15:12]),
        .S({\u_fadd_m23/r_mats[15]_i_2_n_0 ,\u_fadd_m23/r_mats[15]_i_3_n_0 ,\u_fadd_m23/r_mats[15]_i_4_n_0 ,\u_fadd_m23/r_mats[15]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[15]_i_1__1 
       (.CI(\r_mats_reg[11]_i_1__1_n_0 ),
        .CO({\r_mats_reg[15]_i_1__1_n_0 ,\r_mats_reg[15]_i_1__1_n_1 ,\r_mats_reg[15]_i_1__1_n_2 ,\r_mats_reg[15]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [15:12]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [15:12]),
        .S({\u_fadd_m0123/r_mats[15]_i_2_n_0 ,\u_fadd_m0123/r_mats[15]_i_3_n_0 ,\u_fadd_m0123/r_mats[15]_i_4_n_0 ,\u_fadd_m0123/r_mats[15]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[15]_i_1__2 
       (.CI(\r_mats_reg[11]_i_1__2_n_0 ),
        .CO({\r_mats_reg[15]_i_1__2_n_0 ,\r_mats_reg[15]_i_1__2_n_1 ,\r_mats_reg[15]_i_1__2_n_2 ,\r_mats_reg[15]_i_1__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_clip/r_f0 [15:12]),
        .O(\u_geo/u_geo_clip/w_mats [15:12]),
        .S({\u_fadd/r_mats[15]_i_2_n_0 ,\u_fadd/r_mats[15]_i_3_n_0 ,\u_fadd/r_mats[15]_i_4_n_0 ,\u_fadd/r_mats[15]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[15]_i_1__3 
       (.CI(\r_mats_reg[11]_i_1__3_n_0 ),
        .CO({\r_mats_reg[15]_i_1__3_n_0 ,\r_mats_reg[15]_i_1__3_n_1 ,\r_mats_reg[15]_i_1__3_n_2 ,\r_mats_reg[15]_i_1__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_viewport/r_f0 [15:12]),
        .O(\u_geo/u_geo_viewport/w_mats [15:12]),
        .S({\u_fadd/r_mats[15]_i_2__0_n_0 ,\u_fadd/r_mats[15]_i_3__0_n_0 ,\u_fadd/r_mats[15]_i_4__0_n_0 ,\u_fadd/r_mats[15]_i_5__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[16]_i_1 
       (.CI(\r_mats_reg[15]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_mats_reg[16]_i_1_n_4 ,\r_mats_reg[16]_i_1_n_5 ,\r_mats_reg[16]_i_1_n_6 ,\u_geo/u_geo_matrix/u_fadd_m01/w_mats [16]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fadd_m01/r_sub }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[16]_i_1__0 
       (.CI(\r_mats_reg[15]_i_1__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_mats_reg[16]_i_1__0_n_4 ,\r_mats_reg[16]_i_1__0_n_5 ,\r_mats_reg[16]_i_1__0_n_6 ,\u_geo/u_geo_matrix/u_fadd_m23/w_mats [16]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fadd_m23/r_sub }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[16]_i_1__1 
       (.CI(\r_mats_reg[15]_i_1__1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_mats_reg[16]_i_1__1_n_4 ,\r_mats_reg[16]_i_1__1_n_5 ,\r_mats_reg[16]_i_1__1_n_6 ,\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [16]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fadd_m0123/r_sub }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[16]_i_1__2 
       (.CI(\r_mats_reg[15]_i_1__2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_mats_reg[16]_i_1__2_n_4 ,\r_mats_reg[16]_i_1__2_n_5 ,\r_mats_reg[16]_i_1__2_n_6 ,\u_geo/u_geo_clip/w_mats [16]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_clip/r_sub }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[16]_i_1__3 
       (.CI(\r_mats_reg[15]_i_1__3_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_mats_reg[16]_i_1__3_n_4 ,\r_mats_reg[16]_i_1__3_n_5 ,\r_mats_reg[16]_i_1__3_n_6 ,\u_geo/u_geo_viewport/w_mats [16]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_viewport/r_sub }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\r_mats_reg[3]_i_1_n_0 ,\r_mats_reg[3]_i_1_n_1 ,\r_mats_reg[3]_i_1_n_2 ,\r_mats_reg[3]_i_1_n_3 }),
        .CYINIT(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [0]),
        .DI({\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [3:1],\u_geo/u_geo_matrix/u_fadd_m01/r_sub }),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [3:0]),
        .S({\u_fadd_m01/r_mats[3]_i_2_n_0 ,\u_fadd_m01/r_mats[3]_i_3_n_0 ,\u_fadd_m01/r_mats[3]_i_4_n_0 ,\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [0]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[3]_i_1__0 
       (.CI(\<const0>__0__0 ),
        .CO({\r_mats_reg[3]_i_1__0_n_0 ,\r_mats_reg[3]_i_1__0_n_1 ,\r_mats_reg[3]_i_1__0_n_2 ,\r_mats_reg[3]_i_1__0_n_3 }),
        .CYINIT(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [0]),
        .DI({\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [3:1],\u_geo/u_geo_matrix/u_fadd_m23/r_sub }),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [3:0]),
        .S({\u_fadd_m23/r_mats[3]_i_2_n_0 ,\u_fadd_m23/r_mats[3]_i_3_n_0 ,\u_fadd_m23/r_mats[3]_i_4_n_0 ,\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [0]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[3]_i_1__1 
       (.CI(\<const0>__0__0 ),
        .CO({\r_mats_reg[3]_i_1__1_n_0 ,\r_mats_reg[3]_i_1__1_n_1 ,\r_mats_reg[3]_i_1__1_n_2 ,\r_mats_reg[3]_i_1__1_n_3 }),
        .CYINIT(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [0]),
        .DI({\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [3:1],\u_geo/u_geo_matrix/u_fadd_m0123/r_sub }),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [3:0]),
        .S({\u_fadd_m0123/r_mats[3]_i_2_n_0 ,\u_fadd_m0123/r_mats[3]_i_3_n_0 ,\u_fadd_m0123/r_mats[3]_i_4_n_0 ,\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [0]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[3]_i_1__2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_mats_reg[3]_i_1__2_n_0 ,\r_mats_reg[3]_i_1__2_n_1 ,\r_mats_reg[3]_i_1__2_n_2 ,\r_mats_reg[3]_i_1__2_n_3 }),
        .CYINIT(\u_geo/u_geo_clip/r_f0 [0]),
        .DI({\u_geo/u_geo_clip/r_f0 [3:1],\u_geo/u_geo_clip/r_sub }),
        .O(\u_geo/u_geo_clip/w_mats [3:0]),
        .S({\u_fadd/r_mats[3]_i_2_n_0 ,\u_fadd/r_mats[3]_i_3_n_0 ,\u_fadd/r_mats[3]_i_4_n_0 ,\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_ }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[3]_i_1__3 
       (.CI(\<const0>__0__0 ),
        .CO({\r_mats_reg[3]_i_1__3_n_0 ,\r_mats_reg[3]_i_1__3_n_1 ,\r_mats_reg[3]_i_1__3_n_2 ,\r_mats_reg[3]_i_1__3_n_3 }),
        .CYINIT(\u_geo/u_geo_viewport/r_f0 [0]),
        .DI({\u_geo/u_geo_viewport/r_f0 [3:1],\u_geo/u_geo_viewport/r_sub }),
        .O(\u_geo/u_geo_viewport/w_mats [3:0]),
        .S({\u_fadd/r_mats[3]_i_2__0_n_0 ,\u_fadd/r_mats[3]_i_3__0_n_0 ,\u_fadd/r_mats[3]_i_4__0_n_0 ,\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_ }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[7]_i_1 
       (.CI(\r_mats_reg[3]_i_1_n_0 ),
        .CO({\r_mats_reg[7]_i_1_n_0 ,\r_mats_reg[7]_i_1_n_1 ,\r_mats_reg[7]_i_1_n_2 ,\r_mats_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [7:4]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [7:4]),
        .S({\u_fadd_m01/r_mats[7]_i_2_n_0 ,\u_fadd_m01/r_mats[7]_i_3_n_0 ,\u_fadd_m01/r_mats[7]_i_4_n_0 ,\u_fadd_m01/r_mats[7]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[7]_i_1__0 
       (.CI(\r_mats_reg[3]_i_1__0_n_0 ),
        .CO({\r_mats_reg[7]_i_1__0_n_0 ,\r_mats_reg[7]_i_1__0_n_1 ,\r_mats_reg[7]_i_1__0_n_2 ,\r_mats_reg[7]_i_1__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [7:4]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [7:4]),
        .S({\u_fadd_m23/r_mats[7]_i_2_n_0 ,\u_fadd_m23/r_mats[7]_i_3_n_0 ,\u_fadd_m23/r_mats[7]_i_4_n_0 ,\u_fadd_m23/r_mats[7]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[7]_i_1__1 
       (.CI(\r_mats_reg[3]_i_1__1_n_0 ),
        .CO({\r_mats_reg[7]_i_1__1_n_0 ,\r_mats_reg[7]_i_1__1_n_1 ,\r_mats_reg[7]_i_1__1_n_2 ,\r_mats_reg[7]_i_1__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [7:4]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [7:4]),
        .S({\u_fadd_m0123/r_mats[7]_i_2_n_0 ,\u_fadd_m0123/r_mats[7]_i_3_n_0 ,\u_fadd_m0123/r_mats[7]_i_4_n_0 ,\u_fadd_m0123/r_mats[7]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[7]_i_1__2 
       (.CI(\r_mats_reg[3]_i_1__2_n_0 ),
        .CO({\r_mats_reg[7]_i_1__2_n_0 ,\r_mats_reg[7]_i_1__2_n_1 ,\r_mats_reg[7]_i_1__2_n_2 ,\r_mats_reg[7]_i_1__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_clip/r_f0 [7:4]),
        .O(\u_geo/u_geo_clip/w_mats [7:4]),
        .S({\u_fadd/r_mats[7]_i_2_n_0 ,\u_fadd/r_mats[7]_i_3_n_0 ,\u_fadd/r_mats[7]_i_4_n_0 ,\u_fadd/r_mats[7]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_mats_reg[7]_i_1__3 
       (.CI(\r_mats_reg[3]_i_1__3_n_0 ),
        .CO({\r_mats_reg[7]_i_1__3_n_0 ,\r_mats_reg[7]_i_1__3_n_1 ,\r_mats_reg[7]_i_1__3_n_2 ,\r_mats_reg[7]_i_1__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_viewport/r_f0 [7:4]),
        .O(\u_geo/u_geo_viewport/w_mats [7:4]),
        .S({\u_fadd/r_mats[7]_i_2__0_n_0 ,\u_fadd/r_mats[7]_i_3__0_n_0 ,\u_fadd/r_mats[7]_i_4__0_n_0 ,\u_fadd/r_mats[7]_i_5__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \r_outcode[5]_i_1 
       (.I0(\u_geo/u_geo_persdiv/r_state [1]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\u_geo/w_state_pd ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \r_outcode[5]_i_1__0 
       (.I0(\u_geo/u_geo_viewport/r_state [2]),
        .I1(\u_geo/u_geo_viewport/r_state [1]),
        .I2(\u_geo/u_geo_viewport/r_state [0]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .O(\u_geo/w_state_view ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_pixel_color[7]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[5]),
        .I2(r_pixel_color),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[2]),
        .I5(s_wb_sel_i[0]),
        .O(\u_sys/r_pixel_color ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \r_pixel_color[7]_i_2 
       (.I0(s_wb_adr_i[6]),
        .I1(s_wb_stb_i),
        .I2(s_wb_we_i),
        .O(r_pixel_color));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_pixel_top_address[13]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[6]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[1]),
        .O(r_pixel_top_address));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_pixel_top_address[21]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[6]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[2]),
        .O(\r_pixel_top_address[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_pixel_top_address[29]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[6]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[3]),
        .O(\r_pixel_top_address[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_pixel_top_address[5]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[6]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[0]),
        .O(\r_pixel_top_address[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0A0ACCCCCACAC0CC)) 
    \r_rd[0]_i_1 
       (.I0(r_rd_reg),
        .I1(\r_rd[0]_i_3_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[6]),
        .I5(\r_rd[0]_i_4_n_0 ),
        .O(\r_rd[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB833B800)) 
    \r_rd[0]_i_10 
       (.I0(w_dma_size[0]),
        .I1(s_wb_adr_i[3]),
        .I2(\u_sys/p_21_in [0]),
        .I3(s_wb_adr_i[2]),
        .I4(w_dma_start),
        .O(r_rd));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[0]_i_11 
       (.I0(w_m03[0]),
        .I1(w_m02[0]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[0]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[0]),
        .O(\r_rd[0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[0]_i_12 
       (.I0(w_m13[0]),
        .I1(w_m12[0]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[0]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[0]),
        .O(\r_rd[0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[0]_i_13 
       (.I0(w_m23[0]),
        .I1(w_m22[0]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[0]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[0]),
        .O(\r_rd[0]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888B888B8BBB888)) 
    \r_rd[0]_i_3 
       (.I0(\r_rd_reg[0]_i_7_n_0 ),
        .I1(\r_rd[31]_i_6_n_0 ),
        .I2(\^m_wb_dat_o [24]),
        .I3(\r_rd[31]_i_4_n_0 ),
        .I4(w_scr_w[0]),
        .I5(\r_rd[31]_i_5_n_0 ),
        .O(\r_rd[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_rd[0]_i_4 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[2]),
        .O(\r_rd[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[0]_i_5 
       (.I0(w_m33[0]),
        .I1(w_m32[0]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[0]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[0]),
        .O(\r_rd[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[0]_i_6 
       (.I0(w_scr_h_m1[0]),
        .I1(w_scr_w_m1[0]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[0]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[0]),
        .O(\r_rd[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[10]_i_1 
       (.I0(\r_rd[10]_i_2_n_0 ),
        .I1(\r_rd[10]_i_3_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[10]_i_4_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[10]_i_5_n_0 ),
        .O(\r_rd[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[10]_i_2 
       (.I0(\r_rd[10]_i_6_n_0 ),
        .I1(\r_rd[10]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[10]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[10]_i_9_n_0 ),
        .O(\r_rd[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000000E2)) 
    \r_rd[10]_i_3 
       (.I0(w_scr_w[10]),
        .I1(s_wb_adr_i[2]),
        .I2(w_pixel_top_address[8]),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[3]),
        .O(\r_rd[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[10]_i_4 
       (.I0(w_scr_h_m1[10]),
        .I1(w_scr_w_m1[10]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[10]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[10]),
        .O(\r_rd[10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[10]_i_5 
       (.I0(w_m33[10]),
        .I1(w_m32[10]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[10]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[10]),
        .O(\r_rd[10]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[10]_i_6 
       (.I0(w_m23[10]),
        .I1(w_m22[10]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[10]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[10]),
        .O(\r_rd[10]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[10]_i_7 
       (.I0(w_m13[10]),
        .I1(w_m12[10]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[10]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[10]),
        .O(\r_rd[10]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[10]_i_8 
       (.I0(w_m03[10]),
        .I1(w_m02[10]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[10]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[10]),
        .O(\r_rd[10]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[10]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[8]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[10]),
        .O(\r_rd[10]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[11]_i_1 
       (.I0(\r_rd[11]_i_2_n_0 ),
        .I1(\r_rd[11]_i_3_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[11]_i_4_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[11]_i_5_n_0 ),
        .O(\r_rd[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[11]_i_2 
       (.I0(\r_rd[11]_i_6_n_0 ),
        .I1(\r_rd[11]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[11]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[11]_i_9_n_0 ),
        .O(\r_rd[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000000E2)) 
    \r_rd[11]_i_3 
       (.I0(w_scr_w[11]),
        .I1(s_wb_adr_i[2]),
        .I2(w_pixel_top_address[9]),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[3]),
        .O(\r_rd[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[11]_i_4 
       (.I0(w_scr_h_m1[11]),
        .I1(w_scr_w_m1[11]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[11]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[11]),
        .O(\r_rd[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[11]_i_5 
       (.I0(w_m33[11]),
        .I1(w_m32[11]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[11]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[11]),
        .O(\r_rd[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[11]_i_6 
       (.I0(w_m23[11]),
        .I1(w_m22[11]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[11]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[11]),
        .O(\r_rd[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[11]_i_7 
       (.I0(w_m13[11]),
        .I1(w_m12[11]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[11]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[11]),
        .O(\r_rd[11]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[11]_i_8 
       (.I0(w_m03[11]),
        .I1(w_m02[11]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[11]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[11]),
        .O(\r_rd[11]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[11]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[9]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[11]),
        .O(\r_rd[11]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[12]_i_1 
       (.I0(\r_rd[12]_i_2_n_0 ),
        .I1(\r_rd[12]_i_3_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[12]_i_4_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[12]_i_5_n_0 ),
        .O(\r_rd[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[12]_i_2 
       (.I0(\r_rd[12]_i_6_n_0 ),
        .I1(\r_rd[12]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[12]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[12]_i_9_n_0 ),
        .O(\r_rd[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000000E2)) 
    \r_rd[12]_i_3 
       (.I0(w_scr_w[12]),
        .I1(s_wb_adr_i[2]),
        .I2(w_pixel_top_address[10]),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[3]),
        .O(\r_rd[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[12]_i_4 
       (.I0(w_scr_h_m1[12]),
        .I1(w_scr_w_m1[12]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[12]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[12]),
        .O(\r_rd[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[12]_i_5 
       (.I0(w_m33[12]),
        .I1(w_m32[12]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[12]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[12]),
        .O(\r_rd[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[12]_i_6 
       (.I0(w_m23[12]),
        .I1(w_m22[12]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[12]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[12]),
        .O(\r_rd[12]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[12]_i_7 
       (.I0(w_m13[12]),
        .I1(w_m12[12]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[12]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[12]),
        .O(\r_rd[12]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[12]_i_8 
       (.I0(w_m03[12]),
        .I1(w_m02[12]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[12]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[12]),
        .O(\r_rd[12]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[12]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[10]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[12]),
        .O(\r_rd[12]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[13]_i_1 
       (.I0(\r_rd[13]_i_2_n_0 ),
        .I1(\r_rd[13]_i_3_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[13]_i_4_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[13]_i_5_n_0 ),
        .O(\r_rd[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[13]_i_2 
       (.I0(\r_rd[13]_i_6_n_0 ),
        .I1(\r_rd[13]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[13]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[13]_i_9_n_0 ),
        .O(\r_rd[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000000E2)) 
    \r_rd[13]_i_3 
       (.I0(w_scr_w[13]),
        .I1(s_wb_adr_i[2]),
        .I2(w_pixel_top_address[11]),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[3]),
        .O(\r_rd[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[13]_i_4 
       (.I0(w_scr_h_m1[13]),
        .I1(w_scr_w_m1[13]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[13]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[13]),
        .O(\r_rd[13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[13]_i_5 
       (.I0(w_m33[13]),
        .I1(w_m32[13]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[13]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[13]),
        .O(\r_rd[13]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[13]_i_6 
       (.I0(w_m23[13]),
        .I1(w_m22[13]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[13]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[13]),
        .O(\r_rd[13]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[13]_i_7 
       (.I0(w_m13[13]),
        .I1(w_m12[13]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[13]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[13]),
        .O(\r_rd[13]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[13]_i_8 
       (.I0(w_m03[13]),
        .I1(w_m02[13]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[13]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[13]),
        .O(\r_rd[13]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[13]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[11]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[13]),
        .O(\r_rd[13]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[14]_i_1 
       (.I0(\r_rd[14]_i_2_n_0 ),
        .I1(\r_rd[14]_i_3_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[14]_i_4_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[14]_i_5_n_0 ),
        .O(\r_rd[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[14]_i_2 
       (.I0(\r_rd[14]_i_6_n_0 ),
        .I1(\r_rd[14]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[14]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[14]_i_9_n_0 ),
        .O(\r_rd[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000000E2)) 
    \r_rd[14]_i_3 
       (.I0(w_scr_w[14]),
        .I1(s_wb_adr_i[2]),
        .I2(w_pixel_top_address[12]),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[3]),
        .O(\r_rd[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[14]_i_4 
       (.I0(w_scr_h_m1[14]),
        .I1(w_scr_w_m1[14]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[14]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[14]),
        .O(\r_rd[14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[14]_i_5 
       (.I0(w_m33[14]),
        .I1(w_m32[14]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[14]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[14]),
        .O(\r_rd[14]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[14]_i_6 
       (.I0(w_m23[14]),
        .I1(w_m22[14]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[14]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[14]),
        .O(\r_rd[14]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[14]_i_7 
       (.I0(w_m13[14]),
        .I1(w_m12[14]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[14]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[14]),
        .O(\r_rd[14]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[14]_i_8 
       (.I0(w_m03[14]),
        .I1(w_m02[14]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[14]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[14]),
        .O(\r_rd[14]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[14]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[12]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[14]),
        .O(\r_rd[14]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE001)) 
    \r_rd[15]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[6]),
        .I3(s_wb_adr_i[5]),
        .O(\u_sys/w_rd [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[15]_i_10 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[13]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[15]),
        .O(\r_rd[15]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[15]_i_2 
       (.I0(\r_rd[15]_i_3_n_0 ),
        .I1(\r_rd[15]_i_4_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[15]_i_5_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[15]_i_6_n_0 ),
        .O(\r_rd[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[15]_i_3 
       (.I0(\r_rd[15]_i_7_n_0 ),
        .I1(\r_rd[15]_i_8_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[15]_i_9_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[15]_i_10_n_0 ),
        .O(\r_rd[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000000E2)) 
    \r_rd[15]_i_4 
       (.I0(w_scr_w[15]),
        .I1(s_wb_adr_i[2]),
        .I2(w_pixel_top_address[13]),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[3]),
        .O(\r_rd[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[15]_i_5 
       (.I0(w_scr_h_m1[15]),
        .I1(w_scr_w_m1[15]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[15]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[15]),
        .O(\r_rd[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[15]_i_6 
       (.I0(w_m33[15]),
        .I1(w_m32[15]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[15]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[15]),
        .O(\r_rd[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[15]_i_7 
       (.I0(w_m23[15]),
        .I1(w_m22[15]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[15]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[15]),
        .O(\r_rd[15]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[15]_i_8 
       (.I0(w_m13[15]),
        .I1(w_m12[15]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[15]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[15]),
        .O(\r_rd[15]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[15]_i_9 
       (.I0(w_m03[15]),
        .I1(w_m02[15]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[15]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[15]),
        .O(\r_rd[15]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0022AA8A20AAAA8A)) 
    \r_rd[16]_i_1 
       (.I0(\r_rd_reg[16]_i_2_n_0 ),
        .I1(s_wb_adr_i[4]),
        .I2(s_wb_adr_i[2]),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_adr_i[3]),
        .O(\r_rd[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \r_rd[16]_i_10 
       (.I0(w_dma_top_address[14]),
        .I1(s_wb_adr_i[3]),
        .I2(w_ccw),
        .I3(s_wb_adr_i[2]),
        .O(\r_rd[16]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \r_rd[16]_i_3 
       (.I0(w_vw[16]),
        .I1(s_wb_adr_i[2]),
        .I2(w_vh[16]),
        .I3(s_wb_adr_i[3]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[16]_i_5_n_0 ),
        .O(\r_rd[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h888888888888B888)) 
    \r_rd[16]_i_4 
       (.I0(\r_rd[16]_i_6_n_0 ),
        .I1(\r_rd[31]_i_6_n_0 ),
        .I2(w_pixel_top_address[14]),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[4]),
        .I5(s_wb_adr_i[3]),
        .O(\r_rd[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[16]_i_5 
       (.I0(w_m33[16]),
        .I1(w_m32[16]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[16]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[16]),
        .O(\r_rd[16]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[16]_i_6 
       (.I0(\r_rd[16]_i_7_n_0 ),
        .I1(\r_rd[16]_i_8_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[16]_i_9_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[16]_i_10_n_0 ),
        .O(\r_rd[16]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[16]_i_7 
       (.I0(w_m23[16]),
        .I1(w_m22[16]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[16]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[16]),
        .O(\r_rd[16]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[16]_i_8 
       (.I0(w_m13[16]),
        .I1(w_m12[16]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[16]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[16]),
        .O(\r_rd[16]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[16]_i_9 
       (.I0(w_m03[16]),
        .I1(w_m02[16]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[16]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[16]),
        .O(\r_rd[16]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \r_rd[17]_i_2 
       (.I0(w_vw[17]),
        .I1(s_wb_adr_i[2]),
        .I2(w_vh[17]),
        .I3(s_wb_adr_i[3]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[17]_i_4_n_0 ),
        .O(\r_rd[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h888888888888B888)) 
    \r_rd[17]_i_3 
       (.I0(\r_rd[17]_i_5_n_0 ),
        .I1(\r_rd[31]_i_6_n_0 ),
        .I2(w_pixel_top_address[15]),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[4]),
        .I5(s_wb_adr_i[3]),
        .O(\r_rd[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[17]_i_4 
       (.I0(w_m33[17]),
        .I1(w_m32[17]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[17]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[17]),
        .O(\r_rd[17]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[17]_i_5 
       (.I0(\r_rd[17]_i_6_n_0 ),
        .I1(\r_rd[17]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[17]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[17]_i_9_n_0 ),
        .O(\r_rd[17]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[17]_i_6 
       (.I0(w_m23[17]),
        .I1(w_m22[17]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[17]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[17]),
        .O(\r_rd[17]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[17]_i_7 
       (.I0(w_m13[17]),
        .I1(w_m12[17]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[17]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[17]),
        .O(\r_rd[17]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[17]_i_8 
       (.I0(w_m03[17]),
        .I1(w_m02[17]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[17]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[17]),
        .O(\r_rd[17]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \r_rd[17]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[2]),
        .I2(w_dma_top_address[15]),
        .O(\r_rd[17]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \r_rd[18]_i_2 
       (.I0(w_vw[18]),
        .I1(s_wb_adr_i[2]),
        .I2(w_vh[18]),
        .I3(s_wb_adr_i[3]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[18]_i_4_n_0 ),
        .O(\r_rd[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h888888888888B888)) 
    \r_rd[18]_i_3 
       (.I0(\r_rd[18]_i_5_n_0 ),
        .I1(\r_rd[31]_i_6_n_0 ),
        .I2(w_pixel_top_address[16]),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[4]),
        .I5(s_wb_adr_i[3]),
        .O(\r_rd[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[18]_i_4 
       (.I0(w_m33[18]),
        .I1(w_m32[18]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[18]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[18]),
        .O(\r_rd[18]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[18]_i_5 
       (.I0(\r_rd[18]_i_6_n_0 ),
        .I1(\r_rd[18]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[18]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[18]_i_9_n_0 ),
        .O(\r_rd[18]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[18]_i_6 
       (.I0(w_m23[18]),
        .I1(w_m22[18]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[18]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[18]),
        .O(\r_rd[18]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[18]_i_7 
       (.I0(w_m13[18]),
        .I1(w_m12[18]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[18]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[18]),
        .O(\r_rd[18]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[18]_i_8 
       (.I0(w_m03[18]),
        .I1(w_m02[18]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[18]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[18]),
        .O(\r_rd[18]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \r_rd[18]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[2]),
        .I2(w_dma_top_address[16]),
        .O(\r_rd[18]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \r_rd[19]_i_2 
       (.I0(w_vw[19]),
        .I1(s_wb_adr_i[2]),
        .I2(w_vh[19]),
        .I3(s_wb_adr_i[3]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[19]_i_4_n_0 ),
        .O(\r_rd[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h888888888888B888)) 
    \r_rd[19]_i_3 
       (.I0(\r_rd[19]_i_5_n_0 ),
        .I1(\r_rd[31]_i_6_n_0 ),
        .I2(w_pixel_top_address[17]),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[4]),
        .I5(s_wb_adr_i[3]),
        .O(\r_rd[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[19]_i_4 
       (.I0(w_m33[19]),
        .I1(w_m32[19]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[19]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[19]),
        .O(\r_rd[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[19]_i_5 
       (.I0(\r_rd[19]_i_6_n_0 ),
        .I1(\r_rd[19]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[19]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[19]_i_9_n_0 ),
        .O(\r_rd[19]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[19]_i_6 
       (.I0(w_m23[19]),
        .I1(w_m22[19]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[19]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[19]),
        .O(\r_rd[19]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[19]_i_7 
       (.I0(w_m13[19]),
        .I1(w_m12[19]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[19]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[19]),
        .O(\r_rd[19]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[19]_i_8 
       (.I0(w_m03[19]),
        .I1(w_m02[19]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[19]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[19]),
        .O(\r_rd[19]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \r_rd[19]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[2]),
        .I2(w_dma_top_address[17]),
        .O(\r_rd[19]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0A0A2A2AAAAAA8A0)) 
    \r_rd[1]_i_1 
       (.I0(\r_rd[1]_i_2_n_0 ),
        .I1(s_wb_adr_i[2]),
        .I2(s_wb_adr_i[5]),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[4]),
        .I5(s_wb_adr_i[6]),
        .O(\r_rd[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \r_rd[1]_i_10 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_size[1]),
        .I2(s_wb_adr_i[2]),
        .O(\r_rd[1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[1]_i_2 
       (.I0(\r_rd[1]_i_3_n_0 ),
        .I1(\r_rd[1]_i_4_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[1]_i_5_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[1]_i_6_n_0 ),
        .O(\r_rd[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[1]_i_3 
       (.I0(\r_rd[1]_i_7_n_0 ),
        .I1(\r_rd[1]_i_8_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[1]_i_9_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[1]_i_10_n_0 ),
        .O(\r_rd[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8A8ABA8)) 
    \r_rd[1]_i_4 
       (.I0(\^m_wb_dat_o [25]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[4]),
        .I3(w_scr_w[1]),
        .I4(s_wb_adr_i[2]),
        .O(\r_rd[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[1]_i_5 
       (.I0(w_scr_h_m1[1]),
        .I1(w_scr_w_m1[1]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[1]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[1]),
        .O(\r_rd[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[1]_i_6 
       (.I0(w_m33[1]),
        .I1(w_m32[1]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[1]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[1]),
        .O(\r_rd[1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[1]_i_7 
       (.I0(w_m23[1]),
        .I1(w_m22[1]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[1]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[1]),
        .O(\r_rd[1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[1]_i_8 
       (.I0(w_m13[1]),
        .I1(w_m12[1]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[1]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[1]),
        .O(\r_rd[1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[1]_i_9 
       (.I0(w_m03[1]),
        .I1(w_m02[1]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[1]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[1]),
        .O(\r_rd[1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \r_rd[20]_i_2 
       (.I0(w_vw[20]),
        .I1(s_wb_adr_i[2]),
        .I2(w_vh[20]),
        .I3(s_wb_adr_i[3]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[20]_i_4_n_0 ),
        .O(\r_rd[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h888888888888B888)) 
    \r_rd[20]_i_3 
       (.I0(\r_rd[20]_i_5_n_0 ),
        .I1(\r_rd[31]_i_6_n_0 ),
        .I2(w_pixel_top_address[18]),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[4]),
        .I5(s_wb_adr_i[3]),
        .O(\r_rd[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[20]_i_4 
       (.I0(w_m33[20]),
        .I1(w_m32[20]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[20]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[20]),
        .O(\r_rd[20]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[20]_i_5 
       (.I0(\r_rd[20]_i_6_n_0 ),
        .I1(\r_rd[20]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[20]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[20]_i_9_n_0 ),
        .O(\r_rd[20]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[20]_i_6 
       (.I0(w_m23[20]),
        .I1(w_m22[20]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[20]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[20]),
        .O(\r_rd[20]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[20]_i_7 
       (.I0(w_m13[20]),
        .I1(w_m12[20]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[20]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[20]),
        .O(\r_rd[20]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[20]_i_8 
       (.I0(w_m03[20]),
        .I1(w_m02[20]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[20]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[20]),
        .O(\r_rd[20]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \r_rd[20]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[2]),
        .I2(w_dma_top_address[18]),
        .O(\r_rd[20]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hE805EA01)) 
    \r_rd[21]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[4]),
        .I3(s_wb_adr_i[6]),
        .I4(s_wb_adr_i[2]),
        .O(\u_sys/w_rd [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \r_rd[21]_i_10 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[2]),
        .I2(w_dma_top_address[19]),
        .O(\r_rd[21]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \r_rd[21]_i_3 
       (.I0(w_vw[21]),
        .I1(s_wb_adr_i[2]),
        .I2(w_vh[21]),
        .I3(s_wb_adr_i[3]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[21]_i_5_n_0 ),
        .O(\r_rd[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h888888888888B888)) 
    \r_rd[21]_i_4 
       (.I0(\r_rd[21]_i_6_n_0 ),
        .I1(\r_rd[31]_i_6_n_0 ),
        .I2(w_pixel_top_address[19]),
        .I3(s_wb_adr_i[2]),
        .I4(s_wb_adr_i[4]),
        .I5(s_wb_adr_i[3]),
        .O(\r_rd[21]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[21]_i_5 
       (.I0(w_m33[21]),
        .I1(w_m32[21]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[21]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[21]),
        .O(\r_rd[21]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[21]_i_6 
       (.I0(\r_rd[21]_i_7_n_0 ),
        .I1(\r_rd[21]_i_8_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[21]_i_9_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[21]_i_10_n_0 ),
        .O(\r_rd[21]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[21]_i_7 
       (.I0(w_m23[21]),
        .I1(w_m22[21]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[21]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[21]),
        .O(\r_rd[21]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[21]_i_8 
       (.I0(w_m13[21]),
        .I1(w_m12[21]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[21]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[21]),
        .O(\r_rd[21]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[21]_i_9 
       (.I0(w_m03[21]),
        .I1(w_m02[21]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[21]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[21]),
        .O(\r_rd[21]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA200000002000)) 
    \r_rd[22]_i_1 
       (.I0(\r_rd[31]_i_3_n_0 ),
        .I1(\r_rd[31]_i_4_n_0 ),
        .I2(\r_rd[31]_i_5_n_0 ),
        .I3(w_pixel_top_address[20]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[22]_i_2_n_0 ),
        .O(\r_rd[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \r_rd[22]_i_2 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_top_address[20]),
        .I4(s_wb_adr_i[5]),
        .O(\r_rd[22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA200000002000)) 
    \r_rd[23]_i_1 
       (.I0(\r_rd[31]_i_3_n_0 ),
        .I1(\r_rd[31]_i_4_n_0 ),
        .I2(\r_rd[31]_i_5_n_0 ),
        .I3(w_pixel_top_address[21]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[23]_i_2_n_0 ),
        .O(\r_rd[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \r_rd[23]_i_2 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_top_address[21]),
        .I4(s_wb_adr_i[5]),
        .O(\r_rd[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA200000002000)) 
    \r_rd[24]_i_1 
       (.I0(\r_rd[31]_i_3_n_0 ),
        .I1(\r_rd[31]_i_4_n_0 ),
        .I2(\r_rd[31]_i_5_n_0 ),
        .I3(w_pixel_top_address[22]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[24]_i_2_n_0 ),
        .O(\r_rd[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \r_rd[24]_i_2 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_top_address[22]),
        .I4(s_wb_adr_i[5]),
        .O(\r_rd[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA200000002000)) 
    \r_rd[25]_i_1 
       (.I0(\r_rd[31]_i_3_n_0 ),
        .I1(\r_rd[31]_i_4_n_0 ),
        .I2(\r_rd[31]_i_5_n_0 ),
        .I3(w_pixel_top_address[23]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[25]_i_2_n_0 ),
        .O(\r_rd[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \r_rd[25]_i_2 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_top_address[23]),
        .I4(s_wb_adr_i[5]),
        .O(\r_rd[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA200000002000)) 
    \r_rd[26]_i_1 
       (.I0(\r_rd[31]_i_3_n_0 ),
        .I1(\r_rd[31]_i_4_n_0 ),
        .I2(\r_rd[31]_i_5_n_0 ),
        .I3(w_pixel_top_address[24]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[26]_i_2_n_0 ),
        .O(\r_rd[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \r_rd[26]_i_2 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_top_address[24]),
        .I4(s_wb_adr_i[5]),
        .O(\r_rd[26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA200000002000)) 
    \r_rd[27]_i_1 
       (.I0(\r_rd[31]_i_3_n_0 ),
        .I1(\r_rd[31]_i_4_n_0 ),
        .I2(\r_rd[31]_i_5_n_0 ),
        .I3(w_pixel_top_address[25]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[27]_i_2_n_0 ),
        .O(\r_rd[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \r_rd[27]_i_2 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_top_address[25]),
        .I4(s_wb_adr_i[5]),
        .O(\r_rd[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA200000002000)) 
    \r_rd[28]_i_1 
       (.I0(\r_rd[31]_i_3_n_0 ),
        .I1(\r_rd[31]_i_4_n_0 ),
        .I2(\r_rd[31]_i_5_n_0 ),
        .I3(w_pixel_top_address[26]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[28]_i_2_n_0 ),
        .O(\r_rd[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \r_rd[28]_i_2 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_top_address[26]),
        .I4(s_wb_adr_i[5]),
        .O(\r_rd[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA200000002000)) 
    \r_rd[29]_i_1 
       (.I0(\r_rd[31]_i_3_n_0 ),
        .I1(\r_rd[31]_i_4_n_0 ),
        .I2(\r_rd[31]_i_5_n_0 ),
        .I3(w_pixel_top_address[27]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[29]_i_2_n_0 ),
        .O(\r_rd[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \r_rd[29]_i_2 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_top_address[27]),
        .I4(s_wb_adr_i[5]),
        .O(\r_rd[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[2]_i_1 
       (.I0(\r_rd[2]_i_2_n_0 ),
        .I1(\r_rd[2]_i_3_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[2]_i_4_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[2]_i_5_n_0 ),
        .O(\r_rd[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[2]_i_2 
       (.I0(\r_rd[2]_i_6_n_0 ),
        .I1(\r_rd[2]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[2]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[2]_i_9_n_0 ),
        .O(\r_rd[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABA8ABABABA8A8A8)) 
    \r_rd[2]_i_3 
       (.I0(\^m_wb_dat_o [26]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[4]),
        .I3(w_pixel_top_address[0]),
        .I4(s_wb_adr_i[2]),
        .I5(w_scr_w[2]),
        .O(\r_rd[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[2]_i_4 
       (.I0(w_scr_h_m1[2]),
        .I1(w_scr_w_m1[2]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[2]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[2]),
        .O(\r_rd[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[2]_i_5 
       (.I0(w_m33[2]),
        .I1(w_m32[2]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[2]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[2]),
        .O(\r_rd[2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[2]_i_6 
       (.I0(w_m23[2]),
        .I1(w_m22[2]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[2]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[2]),
        .O(\r_rd[2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[2]_i_7 
       (.I0(w_m13[2]),
        .I1(w_m12[2]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[2]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[2]),
        .O(\r_rd[2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[2]_i_8 
       (.I0(w_m03[2]),
        .I1(w_m02[2]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[2]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[2]),
        .O(\r_rd[2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[2]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[0]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[2]),
        .O(\r_rd[2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA200000002000)) 
    \r_rd[30]_i_1 
       (.I0(\r_rd[31]_i_3_n_0 ),
        .I1(\r_rd[31]_i_4_n_0 ),
        .I2(\r_rd[31]_i_5_n_0 ),
        .I3(w_pixel_top_address[28]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[30]_i_2_n_0 ),
        .O(\r_rd[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \r_rd[30]_i_2 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_top_address[28]),
        .I4(s_wb_adr_i[5]),
        .O(\r_rd[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFBFFD)) 
    \r_rd[31]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[2]),
        .I2(s_wb_adr_i[5]),
        .I3(s_wb_adr_i[6]),
        .I4(s_wb_adr_i[4]),
        .O(\u_sys/w_rd [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA200000002000)) 
    \r_rd[31]_i_2 
       (.I0(\r_rd[31]_i_3_n_0 ),
        .I1(\r_rd[31]_i_4_n_0 ),
        .I2(\r_rd[31]_i_5_n_0 ),
        .I3(w_pixel_top_address[29]),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[31]_i_7_n_0 ),
        .O(\r_rd[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \r_rd[31]_i_3 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[6]),
        .O(\r_rd[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_rd[31]_i_4 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[4]),
        .O(\r_rd[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBA)) 
    \r_rd[31]_i_5 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[2]),
        .O(\r_rd[31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h5D)) 
    \r_rd[31]_i_6 
       (.I0(s_wb_adr_i[6]),
        .I1(s_wb_adr_i[4]),
        .I2(s_wb_adr_i[5]),
        .O(\r_rd[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \r_rd[31]_i_7 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_top_address[29]),
        .I4(s_wb_adr_i[5]),
        .O(\r_rd[31]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[3]_i_1 
       (.I0(\r_rd[3]_i_2_n_0 ),
        .I1(\r_rd[3]_i_3_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[3]_i_4_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[3]_i_5_n_0 ),
        .O(\r_rd[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[3]_i_2 
       (.I0(\r_rd[3]_i_6_n_0 ),
        .I1(\r_rd[3]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[3]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[3]_i_9_n_0 ),
        .O(\r_rd[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABA8ABABABA8A8A8)) 
    \r_rd[3]_i_3 
       (.I0(\^m_wb_dat_o [27]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[4]),
        .I3(w_pixel_top_address[1]),
        .I4(s_wb_adr_i[2]),
        .I5(w_scr_w[3]),
        .O(\r_rd[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[3]_i_4 
       (.I0(w_scr_h_m1[3]),
        .I1(w_scr_w_m1[3]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[3]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[3]),
        .O(\r_rd[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[3]_i_5 
       (.I0(w_m33[3]),
        .I1(w_m32[3]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[3]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[3]),
        .O(\r_rd[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[3]_i_6 
       (.I0(w_m23[3]),
        .I1(w_m22[3]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[3]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[3]),
        .O(\r_rd[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[3]_i_7 
       (.I0(w_m13[3]),
        .I1(w_m12[3]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[3]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[3]),
        .O(\r_rd[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[3]_i_8 
       (.I0(w_m03[3]),
        .I1(w_m02[3]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[3]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[3]),
        .O(\r_rd[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[3]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[1]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[3]),
        .O(\r_rd[3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[4]_i_1 
       (.I0(\r_rd[4]_i_2_n_0 ),
        .I1(\r_rd[4]_i_3_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[4]_i_4_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[4]_i_5_n_0 ),
        .O(\r_rd[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[4]_i_2 
       (.I0(\r_rd[4]_i_6_n_0 ),
        .I1(\r_rd[4]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[4]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[4]_i_9_n_0 ),
        .O(\r_rd[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABA8ABABABA8A8A8)) 
    \r_rd[4]_i_3 
       (.I0(\^m_wb_dat_o [28]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[4]),
        .I3(w_pixel_top_address[2]),
        .I4(s_wb_adr_i[2]),
        .I5(w_scr_w[4]),
        .O(\r_rd[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[4]_i_4 
       (.I0(w_scr_h_m1[4]),
        .I1(w_scr_w_m1[4]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[4]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[4]),
        .O(\r_rd[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[4]_i_5 
       (.I0(w_m33[4]),
        .I1(w_m32[4]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[4]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[4]),
        .O(\r_rd[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[4]_i_6 
       (.I0(w_m23[4]),
        .I1(w_m22[4]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[4]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[4]),
        .O(\r_rd[4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[4]_i_7 
       (.I0(w_m13[4]),
        .I1(w_m12[4]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[4]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[4]),
        .O(\r_rd[4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[4]_i_8 
       (.I0(w_m03[4]),
        .I1(w_m02[4]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[4]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[4]),
        .O(\r_rd[4]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[4]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[2]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[4]),
        .O(\r_rd[4]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[5]_i_1 
       (.I0(\r_rd[5]_i_2_n_0 ),
        .I1(\r_rd[5]_i_3_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[5]_i_4_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[5]_i_5_n_0 ),
        .O(\r_rd[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[5]_i_2 
       (.I0(\r_rd[5]_i_6_n_0 ),
        .I1(\r_rd[5]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[5]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[5]_i_9_n_0 ),
        .O(\r_rd[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABA8ABABABA8A8A8)) 
    \r_rd[5]_i_3 
       (.I0(\^m_wb_dat_o [29]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[4]),
        .I3(w_pixel_top_address[3]),
        .I4(s_wb_adr_i[2]),
        .I5(w_scr_w[5]),
        .O(\r_rd[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[5]_i_4 
       (.I0(w_scr_h_m1[5]),
        .I1(w_scr_w_m1[5]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[5]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[5]),
        .O(\r_rd[5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[5]_i_5 
       (.I0(w_m33[5]),
        .I1(w_m32[5]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[5]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[5]),
        .O(\r_rd[5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[5]_i_6 
       (.I0(w_m23[5]),
        .I1(w_m22[5]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[5]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[5]),
        .O(\r_rd[5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[5]_i_7 
       (.I0(w_m13[5]),
        .I1(w_m12[5]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[5]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[5]),
        .O(\r_rd[5]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[5]_i_8 
       (.I0(w_m03[5]),
        .I1(w_m02[5]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[5]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[5]),
        .O(\r_rd[5]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[5]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[3]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[5]),
        .O(\r_rd[5]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[6]_i_1 
       (.I0(\r_rd[6]_i_2_n_0 ),
        .I1(\r_rd[6]_i_3_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[6]_i_4_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[6]_i_5_n_0 ),
        .O(\r_rd[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[6]_i_2 
       (.I0(\r_rd[6]_i_6_n_0 ),
        .I1(\r_rd[6]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[6]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[6]_i_9_n_0 ),
        .O(\r_rd[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABA8ABABABA8A8A8)) 
    \r_rd[6]_i_3 
       (.I0(\^m_wb_dat_o [30]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[4]),
        .I3(w_pixel_top_address[4]),
        .I4(s_wb_adr_i[2]),
        .I5(w_scr_w[6]),
        .O(\r_rd[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[6]_i_4 
       (.I0(w_scr_h_m1[6]),
        .I1(w_scr_w_m1[6]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[6]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[6]),
        .O(\r_rd[6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[6]_i_5 
       (.I0(w_m33[6]),
        .I1(w_m32[6]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[6]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[6]),
        .O(\r_rd[6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[6]_i_6 
       (.I0(w_m23[6]),
        .I1(w_m22[6]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[6]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[6]),
        .O(\r_rd[6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[6]_i_7 
       (.I0(w_m13[6]),
        .I1(w_m12[6]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[6]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[6]),
        .O(\r_rd[6]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[6]_i_8 
       (.I0(w_m03[6]),
        .I1(w_m02[6]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[6]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[6]),
        .O(\r_rd[6]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[6]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[4]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[6]),
        .O(\r_rd[6]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC0C08003)) 
    \r_rd[7]_i_1 
       (.I0(s_wb_adr_i[2]),
        .I1(s_wb_adr_i[6]),
        .I2(s_wb_adr_i[5]),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[4]),
        .O(\u_sys/w_rd [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[7]_i_10 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[5]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[7]),
        .O(\r_rd[7]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[7]_i_2 
       (.I0(\r_rd[7]_i_3_n_0 ),
        .I1(\r_rd[7]_i_4_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[7]_i_5_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[7]_i_6_n_0 ),
        .O(\r_rd[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[7]_i_3 
       (.I0(\r_rd[7]_i_7_n_0 ),
        .I1(\r_rd[7]_i_8_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[7]_i_9_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[7]_i_10_n_0 ),
        .O(\r_rd[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABA8ABABABA8A8A8)) 
    \r_rd[7]_i_4 
       (.I0(\^m_wb_dat_o [31]),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[4]),
        .I3(w_pixel_top_address[5]),
        .I4(s_wb_adr_i[2]),
        .I5(w_scr_w[7]),
        .O(\r_rd[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[7]_i_5 
       (.I0(w_scr_h_m1[7]),
        .I1(w_scr_w_m1[7]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[7]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[7]),
        .O(\r_rd[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[7]_i_6 
       (.I0(w_m33[7]),
        .I1(w_m32[7]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[7]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[7]),
        .O(\r_rd[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[7]_i_7 
       (.I0(w_m23[7]),
        .I1(w_m22[7]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[7]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[7]),
        .O(\r_rd[7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[7]_i_8 
       (.I0(w_m13[7]),
        .I1(w_m12[7]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[7]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[7]),
        .O(\r_rd[7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[7]_i_9 
       (.I0(w_m03[7]),
        .I1(w_m02[7]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[7]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[7]),
        .O(\r_rd[7]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2A2A2AAA2AAA2AAA)) 
    \r_rd[8]_i_1 
       (.I0(\r_rd[8]_i_2_n_0 ),
        .I1(s_wb_adr_i[6]),
        .I2(s_wb_adr_i[5]),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[2]),
        .I5(s_wb_adr_i[3]),
        .O(\r_rd[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[8]_i_10 
       (.I0(w_m03[8]),
        .I1(w_m02[8]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[8]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[8]),
        .O(\r_rd[8]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[8]_i_11 
       (.I0(w_m13[8]),
        .I1(w_m12[8]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[8]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[8]),
        .O(\r_rd[8]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[8]_i_12 
       (.I0(w_m23[8]),
        .I1(w_m22[8]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[8]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[8]),
        .O(\r_rd[8]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[8]_i_2 
       (.I0(\r_rd_reg[8]_i_3_n_0 ),
        .I1(\r_rd[8]_i_4_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[8]_i_5_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[8]_i_6_n_0 ),
        .O(\r_rd[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hABA8ABABABA8A8A8)) 
    \r_rd[8]_i_4 
       (.I0(w_y_flip),
        .I1(s_wb_adr_i[3]),
        .I2(s_wb_adr_i[4]),
        .I3(w_pixel_top_address[6]),
        .I4(s_wb_adr_i[2]),
        .I5(w_scr_w[8]),
        .O(\r_rd[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[8]_i_5 
       (.I0(w_scr_h_m1[8]),
        .I1(w_scr_w_m1[8]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[8]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[8]),
        .O(\r_rd[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[8]_i_6 
       (.I0(w_m33[8]),
        .I1(w_m32[8]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[8]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[8]),
        .O(\r_rd[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[8]_i_9 
       (.I0(w_dma_size[8]),
        .I1(w_dma_top_address[6]),
        .I2(s_wb_adr_i[3]),
        .I3(\u_sys/p_21_in [8]),
        .I4(s_wb_adr_i[2]),
        .I5(w_en_cull),
        .O(\r_rd[8]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[9]_i_1 
       (.I0(\r_rd[9]_i_2_n_0 ),
        .I1(\r_rd[9]_i_3_n_0 ),
        .I2(\r_rd[31]_i_3_n_0 ),
        .I3(\r_rd[9]_i_4_n_0 ),
        .I4(\r_rd[31]_i_6_n_0 ),
        .I5(\r_rd[9]_i_5_n_0 ),
        .O(\r_rd[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[9]_i_2 
       (.I0(\r_rd[9]_i_6_n_0 ),
        .I1(\r_rd[9]_i_7_n_0 ),
        .I2(s_wb_adr_i[5]),
        .I3(\r_rd[9]_i_8_n_0 ),
        .I4(s_wb_adr_i[4]),
        .I5(\r_rd[9]_i_9_n_0 ),
        .O(\r_rd[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000000E2)) 
    \r_rd[9]_i_3 
       (.I0(w_scr_w[9]),
        .I1(s_wb_adr_i[2]),
        .I2(w_pixel_top_address[7]),
        .I3(s_wb_adr_i[4]),
        .I4(s_wb_adr_i[3]),
        .O(\r_rd[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[9]_i_4 
       (.I0(w_scr_h_m1[9]),
        .I1(w_scr_w_m1[9]),
        .I2(s_wb_adr_i[3]),
        .I3(w_vh[9]),
        .I4(s_wb_adr_i[2]),
        .I5(w_vw[9]),
        .O(\r_rd[9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[9]_i_5 
       (.I0(w_m33[9]),
        .I1(w_m32[9]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m31[9]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m30[9]),
        .O(\r_rd[9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[9]_i_6 
       (.I0(w_m23[9]),
        .I1(w_m22[9]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m21[9]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m20[9]),
        .O(\r_rd[9]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[9]_i_7 
       (.I0(w_m13[9]),
        .I1(w_m12[9]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m11[9]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m10[9]),
        .O(\r_rd[9]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_rd[9]_i_8 
       (.I0(w_m03[9]),
        .I1(w_m02[9]),
        .I2(s_wb_adr_i[3]),
        .I3(w_m01[9]),
        .I4(s_wb_adr_i[2]),
        .I5(w_m00[9]),
        .O(\r_rd[9]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \r_rd[9]_i_9 
       (.I0(s_wb_adr_i[3]),
        .I1(w_dma_top_address[7]),
        .I2(s_wb_adr_i[2]),
        .I3(w_dma_size[9]),
        .O(\r_rd[9]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_rd_reg[0]_i_2 
       (.I0(\r_rd[0]_i_5_n_0 ),
        .I1(\r_rd[0]_i_6_n_0 ),
        .O(r_rd_reg),
        .S(\r_rd[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \r_rd_reg[0]_i_7 
       (.I0(\r_rd_reg[0]_i_8_n_0 ),
        .I1(\r_rd_reg[0]_i_9_n_0 ),
        .O(\r_rd_reg[0]_i_7_n_0 ),
        .S(s_wb_adr_i[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_rd_reg[0]_i_8 
       (.I0(r_rd),
        .I1(\r_rd[0]_i_11_n_0 ),
        .O(\r_rd_reg[0]_i_8_n_0 ),
        .S(s_wb_adr_i[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_rd_reg[0]_i_9 
       (.I0(\r_rd[0]_i_12_n_0 ),
        .I1(\r_rd[0]_i_13_n_0 ),
        .O(\r_rd_reg[0]_i_9_n_0 ),
        .S(s_wb_adr_i[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_rd_reg[16]_i_2 
       (.I0(\r_rd[16]_i_3_n_0 ),
        .I1(\r_rd[16]_i_4_n_0 ),
        .O(\r_rd_reg[16]_i_2_n_0 ),
        .S(\r_rd[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_rd_reg[17]_i_1 
       (.I0(\r_rd[17]_i_2_n_0 ),
        .I1(\r_rd[17]_i_3_n_0 ),
        .O(\r_rd_reg[17]_i_1_n_0 ),
        .S(\r_rd[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_rd_reg[18]_i_1 
       (.I0(\r_rd[18]_i_2_n_0 ),
        .I1(\r_rd[18]_i_3_n_0 ),
        .O(\r_rd_reg[18]_i_1_n_0 ),
        .S(\r_rd[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_rd_reg[19]_i_1 
       (.I0(\r_rd[19]_i_2_n_0 ),
        .I1(\r_rd[19]_i_3_n_0 ),
        .O(\r_rd_reg[19]_i_1_n_0 ),
        .S(\r_rd[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_rd_reg[20]_i_1 
       (.I0(\r_rd[20]_i_2_n_0 ),
        .I1(\r_rd[20]_i_3_n_0 ),
        .O(\r_rd_reg[20]_i_1_n_0 ),
        .S(\r_rd[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_rd_reg[21]_i_2 
       (.I0(\r_rd[21]_i_3_n_0 ),
        .I1(\r_rd[21]_i_4_n_0 ),
        .O(\r_rd_reg[21]_i_2_n_0 ),
        .S(\r_rd[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \r_rd_reg[8]_i_3 
       (.I0(\r_rd_reg[8]_i_7_n_0 ),
        .I1(\r_rd_reg[8]_i_8_n_0 ),
        .O(\r_rd_reg[8]_i_3_n_0 ),
        .S(s_wb_adr_i[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_rd_reg[8]_i_7 
       (.I0(\r_rd[8]_i_9_n_0 ),
        .I1(\r_rd[8]_i_10_n_0 ),
        .O(\r_rd_reg[8]_i_7_n_0 ),
        .S(s_wb_adr_i[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_rd_reg[8]_i_8 
       (.I0(\r_rd[8]_i_11_n_0 ),
        .I1(\r_rd[8]_i_12_n_0 ),
        .O(\r_rd_reg[8]_i_8_n_0 ),
        .S(s_wb_adr_i[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0044)) 
    r_req_geo_i_1
       (.I0(m_wb_ack_i),
        .I1(w_req_geo),
        .I2(\u_ras/u_ras_mem/r_state ),
        .I3(\u_mem_arb/r_state ),
        .I4(\u_mem_arb/r_req_geo ),
        .O(r_req_geo_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    r_rstr_i_1
       (.I0(s_wb_stb_i),
        .I1(s_wb_we_i),
        .O(r_rstr_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \r_scr_h_m1[15]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[1]),
        .O(r_scr_h_m1));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \r_scr_h_m1[7]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[4]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[6]),
        .I5(s_wb_sel_i[0]),
        .O(\r_scr_h_m1[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_scr_w[15]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[4]),
        .I2(r_pixel_color),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[2]),
        .I5(s_wb_sel_i[1]),
        .O(r_scr_w));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_scr_w[7]_i_1 
       (.I0(s_wb_adr_i[5]),
        .I1(s_wb_adr_i[4]),
        .I2(r_pixel_color),
        .I3(s_wb_adr_i[3]),
        .I4(s_wb_adr_i[2]),
        .I5(s_wb_sel_i[0]),
        .O(\r_scr_w[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_scr_w_m1[15]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[6]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[2]),
        .I5(s_wb_sel_i[1]),
        .O(r_scr_w_m1));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_scr_w_m1[7]_i_1 
       (.I0(s_wb_adr_i[3]),
        .I1(s_wb_adr_i[6]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[2]),
        .I5(s_wb_sel_i[0]),
        .O(\r_scr_w_m1[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    r_sign_1z_i_1
       (.I0(\u_geo/u_geo_matrix/r_vx_in [21]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/w_vx_dma [21]),
        .I3(r_sign_1z_i_2_n_0),
        .I4(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I5(w_m10[21]),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/w_sign ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    r_sign_1z_i_1__0
       (.I0(\u_geo/u_geo_matrix/r_vy_in [21]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/w_vy_dma [21]),
        .I3(r_sign_1z_i_2__0_n_0),
        .I4(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I5(w_m11[21]),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/w_sign ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D1D1DE2E2E21DE2)) 
    r_sign_1z_i_1__1
       (.I0(\u_geo/u_geo_matrix/r_vz_in [21]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/w_vz_dma [21]),
        .I3(r_sign_1z_i_2__1_n_0),
        .I4(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I5(w_m12[21]),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/w_sign ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_sign_1z_i_1__2
       (.I0(\u_geo/u_geo_matrix/w_m0_out [21]),
        .I1(\r_f0[15]_i_2__0_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m1_out [21]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_sign ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_sign_1z_i_1__3
       (.I0(\u_geo/u_geo_matrix/w_m2_out [21]),
        .I1(\r_f0[15]_i_2__1_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_m3_out [21]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_sign ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_sign_1z_i_1__4
       (.I0(\u_geo/u_geo_matrix/w_add01_out [21]),
        .I1(\r_f0[15]_i_2__2_n_0 ),
        .I2(\u_geo/u_geo_matrix/w_add23_out [21]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_sign ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_sign_1z_i_1__5
       (.I0(w_m13[21]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(r_sign_1z_i_2__2_n_0),
        .O(r_sign_1z_i_1__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B800FF)) 
    r_sign_1z_i_1__6
       (.I0(\u_geo/w_vw_mvp [21]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [21]),
        .I3(r_sub_i_2_n_0),
        .I4(\r_f0[15]_i_2__3_n_0 ),
        .O(\u_geo/u_geo_clip/u_fadd/w_sign ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h474747B8B8B847B8)) 
    r_sign_1z_i_1__7
       (.I0(\u_geo/w_vx_pdiv [21]),
        .I1(\r_ce_tmp_1z[4]_i_3__2_n_0 ),
        .I2(\u_geo/w_vy_pdiv [21]),
        .I3(\u_geo/u_geo_persdiv/r_ivw [21]),
        .I4(r_ivw),
        .I5(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[21] ),
        .O(\u_geo/u_geo_persdiv/u_fmul/w_sign ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    r_sign_1z_i_1__8
       (.I0(\u_geo/u_geo_viewport/w_fadd_out ),
        .I1(\r_ce_tmp_1z[4]_i_3__3_n_0 ),
        .I2(w_vh[21]),
        .I3(w_vw[21]),
        .O(\u_geo/u_geo_viewport/u_fmul/w_sign ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    r_sign_1z_i_2
       (.I0(w_m20[21]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[21]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[21]),
        .O(r_sign_1z_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    r_sign_1z_i_2__0
       (.I0(w_m21[21]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[21]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[21]),
        .O(r_sign_1z_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    r_sign_1z_i_2__1
       (.I0(w_m22[21]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[21]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[21]),
        .O(r_sign_1z_i_2__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    r_sign_1z_i_2__2
       (.I0(w_m23[21]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[21]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[21]),
        .O(r_sign_1z_i_2__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00FE)) 
    \r_size[0]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\u_geo/u_geo_mem/r_size__0 [0]),
        .O(r_size));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[10]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[12]_i_2_n_6 ),
        .O(\u_geo/u_geo_mem/r_size [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[11]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[12]_i_2_n_5 ),
        .O(\u_geo/u_geo_mem/r_size [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[12]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[12]_i_2_n_4 ),
        .O(\u_geo/u_geo_mem/r_size [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[13]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[15]_i_3_n_7 ),
        .O(\u_geo/u_geo_mem/r_size [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[14]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[15]_i_3_n_6 ),
        .O(\u_geo/u_geo_mem/r_size [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF8888888)) 
    \r_size[15]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .I1(w_dma_start),
        .I2(m_wb_ack_i),
        .I3(\u_mem_arb/w_pri__0 ),
        .I4(\FSM_onehot_r_state[5]_i_4_n_0 ),
        .O(\r_size[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[15]_i_2 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[15]_i_3_n_5 ),
        .O(\u_geo/u_geo_mem/r_size [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[1]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[4]_i_2_n_7 ),
        .O(\u_geo/u_geo_mem/r_size [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[2]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[4]_i_2_n_6 ),
        .O(\u_geo/u_geo_mem/r_size [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[3]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[4]_i_2_n_5 ),
        .O(\u_geo/u_geo_mem/r_size [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[4]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[4]_i_2_n_4 ),
        .O(\u_geo/u_geo_mem/r_size [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[5]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[8]_i_2_n_7 ),
        .O(\u_geo/u_geo_mem/r_size [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[6]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[8]_i_2_n_6 ),
        .O(\u_geo/u_geo_mem/r_size [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[7]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[8]_i_2_n_5 ),
        .O(\u_geo/u_geo_mem/r_size [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[8]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[8]_i_2_n_4 ),
        .O(\u_geo/u_geo_mem/r_size [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_size[9]_i_1 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(\r_size_reg[12]_i_2_n_7 ),
        .O(\u_geo/u_geo_mem/r_size [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_size_reg[12]_i_2 
       (.CI(\r_size_reg[8]_i_2_n_0 ),
        .CO(r_size_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_size_reg[12]_i_2_n_4 ,\r_size_reg[12]_i_2_n_5 ,\r_size_reg[12]_i_2_n_6 ,\r_size_reg[12]_i_2_n_7 }),
        .S(\u_geo/u_geo_mem/r_size__0 [12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_size_reg[15]_i_3 
       (.CI(r_size_reg[3]),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_size_reg[15]_i_3_n_4 ,\r_size_reg[15]_i_3_n_5 ,\r_size_reg[15]_i_3_n_6 ,\r_size_reg[15]_i_3_n_7 }),
        .S({\<const0>__0__0 ,\u_geo/u_geo_mem/r_size__0 [15:13]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_size_reg[4]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_size_reg[4]_i_2_n_0 ,\r_size_reg[4]_i_2_n_1 ,\r_size_reg[4]_i_2_n_2 ,\r_size_reg[4]_i_2_n_3 }),
        .CYINIT(\u_geo/u_geo_mem/r_size__0 [0]),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_size_reg[4]_i_2_n_4 ,\r_size_reg[4]_i_2_n_5 ,\r_size_reg[4]_i_2_n_6 ,\r_size_reg[4]_i_2_n_7 }),
        .S(\u_geo/u_geo_mem/r_size__0 [4:1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_size_reg[8]_i_2 
       (.CI(\r_size_reg[4]_i_2_n_0 ),
        .CO({\r_size_reg[8]_i_2_n_0 ,\r_size_reg[8]_i_2_n_1 ,\r_size_reg[8]_i_2_n_2 ,\r_size_reg[8]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_size_reg[8]_i_2_n_4 ,\r_size_reg[8]_i_2_n_5 ,\r_size_reg[8]_i_2_n_6 ,\r_size_reg[8]_i_2_n_7 }),
        .S(\u_geo/u_geo_mem/r_size__0 [8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h44FC)) 
    \r_state[0]_i_1 
       (.I0(\r_state[1]_i_2_n_0 ),
        .I1(\u_geo/u_geo_cull/r_state [1]),
        .I2(\u_geo/w_en_tri ),
        .I3(\u_geo/u_geo_cull/r_state [0]),
        .O(r_state));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h33DCFFDC)) 
    \r_state[1]_i_1 
       (.I0(w_en_cull),
        .I1(\u_geo/u_geo_cull/r_state [0]),
        .I2(\u_geo/w_en_tri ),
        .I3(\u_geo/u_geo_cull/r_state [1]),
        .I4(\r_state[1]_i_2_n_0 ),
        .O(\r_state[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF11111F1)) 
    \r_state[1]_i_2 
       (.I0(\u_ras/u_ras_state/r_state [1]),
        .I1(\u_ras/u_ras_state/r_state [0]),
        .I2(w_en_cull),
        .I3(w_ccw),
        .I4(\u_geo/u_geo_cull/p_0_in ),
        .O(\r_state[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAABBAFAAFFBBAFAA)) 
    \r_state[1]_i_3 
       (.I0(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .I1(\u_ras/u_ras_state/f_reject0_return ),
        .I2(\u_ras/u_ras_state/f_reject_return ),
        .I3(\u_ras/u_ras_state/r_state [0]),
        .I4(\u_ras/u_ras_state/r_state [1]),
        .I5(\u_ras/u_ras_state/f_reject1_return ),
        .O(\r_state[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFFFFE)) 
    \r_state[1]_i_4 
       (.I0(\u_ras/w_y ),
        .I1(\u_ras/u_ras_line/w_reject1__7 ),
        .I2(\u_ras/w_x ),
        .I3(\u_ras/u_ras_line/w_reject0__7 ),
        .I4(\u_ras/w_ack_pix ),
        .I5(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_state[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \r_state[1]_i_5 
       (.I0(\u_ras/u_ras_mem/r_state ),
        .I1(\u_mem_arb/w_pri__0 ),
        .I2(m_wb_ack_i),
        .O(\u_ras/w_ack_pix ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFD0)) 
    r_state_i_1
       (.I0(m_wb_ack_i),
        .I1(\u_mem_arb/w_pri__0 ),
        .I2(\u_ras/u_ras_mem/r_state ),
        .I3(\u_ras/w_en_pix ),
        .O(r_state_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFFFFE)) 
    r_state_i_1__0
       (.I0(\u_mem_arb/r_state ),
        .I1(\u_ras/u_ras_mem/r_state ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I3(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I4(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I5(m_wb_ack_i),
        .O(r_state_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \r_state_reg[1]_i_2 
       (.I0(\r_state[1]_i_3_n_0 ),
        .I1(\r_state[1]_i_4_n_0 ),
        .O(r_state_reg),
        .S(\u_ras/u_ras_line/r_state_reg_n_0_ ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    r_sub_i_1
       (.I0(\u_geo/u_geo_matrix/w_m0_out [21]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [21]),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/w_sub11_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    r_sub_i_1__0
       (.I0(\u_geo/u_geo_matrix/w_m2_out [21]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [21]),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/w_sub11_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    r_sub_i_1__1
       (.I0(\u_geo/u_geo_matrix/w_add01_out [21]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [21]),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/w_sub11_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAA8)) 
    r_sub_i_1__2
       (.I0(\u_geo/w_vy_pdiv [21]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .I5(\u_geo/w_vx_pdiv [21]),
        .O(\u_geo/u_geo_viewport/w_fadd_a [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE21D)) 
    r_sub_i_1__3
       (.I0(\u_geo/w_vw_clip [21]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_mvp [21]),
        .I3(r_sub_i_2_n_0),
        .O(r_sub_i_1__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hAAA9)) 
    r_sub_i_2
       (.I0(r_sub_i_3_n_0),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(\u_geo/w_state_clip ),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .O(r_sub_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCAACCAACCAACCF0)) 
    r_sub_i_3
       (.I0(\u_geo/w_vy_clip [21]),
        .I1(\u_geo/w_vx_clip [21]),
        .I2(r_sub_i_4_n_0),
        .I3(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .I4(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .I5(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(r_sub_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    r_sub_i_4
       (.I0(\u_geo/u_geo_clip/r_vz [21]),
        .I1(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .I3(\u_geo/w_vx_mvp [21]),
        .O(r_sub_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[0]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [0]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_105 ),
        .O(\u_geo/u_geo_cull/p_1_in [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[10]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [10]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_95 ),
        .O(\u_geo/u_geo_cull/p_1_in [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[11]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [11]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_94 ),
        .O(\u_geo/u_geo_cull/p_1_in [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[11]_i_3 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[11] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_94 ),
        .O(r_sum));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[11]_i_4 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[10] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_95 ),
        .O(\r_sum[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[11]_i_5 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[9] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_96 ),
        .O(\r_sum[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[11]_i_6 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[8] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_97 ),
        .O(\r_sum[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[12]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [12]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_93 ),
        .O(\u_geo/u_geo_cull/p_1_in [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[13]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [13]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_92 ),
        .O(\u_geo/u_geo_cull/p_1_in [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[14]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [14]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_91 ),
        .O(\u_geo/u_geo_cull/p_1_in [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[15]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [15]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_90 ),
        .O(\u_geo/u_geo_cull/p_1_in [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[15]_i_3 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[15] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_90 ),
        .O(\r_sum[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[15]_i_4 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[14] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_91 ),
        .O(\r_sum[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[15]_i_5 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[13] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_92 ),
        .O(\r_sum[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[15]_i_6 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[12] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_93 ),
        .O(\r_sum[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[16]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [16]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_89 ),
        .O(\u_geo/u_geo_cull/p_1_in [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[17]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [17]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_88 ),
        .O(\u_geo/u_geo_cull/p_1_in [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[18]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [18]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_87 ),
        .O(\u_geo/u_geo_cull/p_1_in [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[19]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [19]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_86 ),
        .O(\u_geo/u_geo_cull/p_1_in [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[19]_i_3 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[19] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_86 ),
        .O(\r_sum[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[19]_i_4 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[18] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_87 ),
        .O(\r_sum[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[19]_i_5 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[17] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_88 ),
        .O(\r_sum[19]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[19]_i_6 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[16] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_89 ),
        .O(\r_sum[19]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[1]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [1]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_104 ),
        .O(\u_geo/u_geo_cull/p_1_in [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[20]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [20]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_85 ),
        .O(\u_geo/u_geo_cull/p_1_in [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[21]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [21]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_84 ),
        .O(\u_geo/u_geo_cull/p_1_in [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[22]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [22]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_83 ),
        .O(\u_geo/u_geo_cull/p_1_in [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEA55EA)) 
    \r_sum[23]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(w_en_cull),
        .I2(\u_geo/w_en_tri ),
        .I3(\u_geo/u_geo_cull/r_state [1]),
        .I4(\r_state[1]_i_2_n_0 ),
        .O(\r_sum[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[23]_i_2 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [23]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_82 ),
        .O(\u_geo/u_geo_cull/p_1_in [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[23]_i_4 
       (.I0(\u_geo/u_geo_cull/p_0_in ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_82 ),
        .O(\r_sum[23]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[23]_i_5 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[22] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_83 ),
        .O(\r_sum[23]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[23]_i_6 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[21] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_84 ),
        .O(\r_sum[23]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[23]_i_7 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[20] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_85 ),
        .O(\r_sum[23]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[2]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [2]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_103 ),
        .O(\u_geo/u_geo_cull/p_1_in [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[3]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [3]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_102 ),
        .O(\u_geo/u_geo_cull/p_1_in [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[3]_i_3 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_102 ),
        .O(\r_sum[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[3]_i_4 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[2] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_103 ),
        .O(\r_sum[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[3]_i_5 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[1] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_104 ),
        .O(\r_sum[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[3]_i_6 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_ ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_105 ),
        .O(\r_sum[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[4]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [4]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_101 ),
        .O(\u_geo/u_geo_cull/p_1_in [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[5]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [5]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_100 ),
        .O(\u_geo/u_geo_cull/p_1_in [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[6]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [6]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_99 ),
        .O(\u_geo/u_geo_cull/p_1_in [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[7]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [7]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_98 ),
        .O(\u_geo/u_geo_cull/p_1_in [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[7]_i_3 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[7] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_98 ),
        .O(\r_sum[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[7]_i_4 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[6] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_99 ),
        .O(\r_sum[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[7]_i_5 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[5] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_100 ),
        .O(\r_sum[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_sum[7]_i_6 
       (.I0(\u_geo/u_geo_cull/r_sum_reg_n_0_[4] ),
        .I1(\u_geo/u_geo_cull/f_multi_return_n_101 ),
        .O(\r_sum[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[8]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [8]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_97 ),
        .O(\u_geo/u_geo_cull/p_1_in [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4D48)) 
    \r_sum[9]_i_1 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_sum0 [9]),
        .I2(\u_geo/u_geo_cull/r_state [1]),
        .I3(\u_geo/u_geo_cull/f_multi_return_n_96 ),
        .O(\u_geo/u_geo_cull/p_1_in [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_sum_reg[11]_i_2 
       (.CI(\r_sum_reg[7]_i_2_n_0 ),
        .CO(r_sum_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\u_geo/u_geo_cull/r_sum_reg_n_0_[11] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[10] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[9] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[8] }),
        .O(\u_geo/u_geo_cull/r_sum0 [11:8]),
        .S({r_sum,\r_sum[11]_i_4_n_0 ,\r_sum[11]_i_5_n_0 ,\r_sum[11]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_sum_reg[15]_i_2 
       (.CI(r_sum_reg[3]),
        .CO({\r_sum_reg[15]_i_2_n_0 ,\r_sum_reg[15]_i_2_n_1 ,\r_sum_reg[15]_i_2_n_2 ,\r_sum_reg[15]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\u_geo/u_geo_cull/r_sum_reg_n_0_[15] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[14] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[13] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[12] }),
        .O(\u_geo/u_geo_cull/r_sum0 [15:12]),
        .S({\r_sum[15]_i_3_n_0 ,\r_sum[15]_i_4_n_0 ,\r_sum[15]_i_5_n_0 ,\r_sum[15]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_sum_reg[19]_i_2 
       (.CI(\r_sum_reg[15]_i_2_n_0 ),
        .CO({\r_sum_reg[19]_i_2_n_0 ,\r_sum_reg[19]_i_2_n_1 ,\r_sum_reg[19]_i_2_n_2 ,\r_sum_reg[19]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\u_geo/u_geo_cull/r_sum_reg_n_0_[19] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[18] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[17] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[16] }),
        .O(\u_geo/u_geo_cull/r_sum0 [19:16]),
        .S({\r_sum[19]_i_3_n_0 ,\r_sum[19]_i_4_n_0 ,\r_sum[19]_i_5_n_0 ,\r_sum[19]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_sum_reg[23]_i_3 
       (.CI(\r_sum_reg[19]_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\u_geo/u_geo_cull/r_sum_reg_n_0_[22] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[21] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[20] }),
        .O(\u_geo/u_geo_cull/r_sum0 [23:20]),
        .S({\r_sum[23]_i_4_n_0 ,\r_sum[23]_i_5_n_0 ,\r_sum[23]_i_6_n_0 ,\r_sum[23]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_sum_reg[3]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_sum_reg[3]_i_2_n_0 ,\r_sum_reg[3]_i_2_n_1 ,\r_sum_reg[3]_i_2_n_2 ,\r_sum_reg[3]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\u_geo/u_geo_cull/r_sum_reg_n_0_[3] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[2] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[1] ,\u_geo/u_geo_cull/r_sum_reg_n_0_ }),
        .O(\u_geo/u_geo_cull/r_sum0 [3:0]),
        .S({\r_sum[3]_i_3_n_0 ,\r_sum[3]_i_4_n_0 ,\r_sum[3]_i_5_n_0 ,\r_sum[3]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_sum_reg[7]_i_2 
       (.CI(\r_sum_reg[3]_i_2_n_0 ),
        .CO({\r_sum_reg[7]_i_2_n_0 ,\r_sum_reg[7]_i_2_n_1 ,\r_sum_reg[7]_i_2_n_2 ,\r_sum_reg[7]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\u_geo/u_geo_cull/r_sum_reg_n_0_[7] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[6] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[5] ,\u_geo/u_geo_cull/r_sum_reg_n_0_[4] }),
        .O(\u_geo/u_geo_cull/r_sum0 [7:4]),
        .S({\r_sum[7]_i_3_n_0 ,\r_sum[7]_i_4_n_0 ,\r_sum[7]_i_5_n_0 ,\r_sum[7]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000008)) 
    \r_v0_outcode[5]_i_1 
       (.I0(\u_geo/w_state_if ),
        .I1(\u_geo/u_geo_viewport/r_state [3]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_tri/w_set_v0_x ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8A80BABF)) 
    \r_v0_x[0]_i_1 
       (.I0(\u_geo/u_geo_tri/w_ui_2c [1]),
        .I1(\u_geo/w_vx_view [21]),
        .I2(\u_geo/u_geo_tri/w_set_y ),
        .I3(\u_geo/u_geo_tri/r_vy [21]),
        .I4(\r_v0_x[3]_i_8_n_0 ),
        .O(\u_geo/u_geo_tri/p_0_in__0 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF084C3B7F)) 
    \r_v0_x[0]_i_2 
       (.I0(\r_v0_x[11]_i_9_n_0 ),
        .I1(\r_v0_x[10]_i_4_n_0 ),
        .I2(r_v0_x),
        .I3(\r_v0_x[4]_i_3_n_0 ),
        .I4(\r_v0_x[8]_i_2_n_0 ),
        .I5(\r_v0_x[10]_i_5_n_0 ),
        .O(\r_v0_x[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFACA0ACA)) 
    \r_v0_x[0]_i_3 
       (.I0(\r_v0_x[2]_i_4_n_0 ),
        .I1(\r_v0_x[0]_i_4_n_0 ),
        .I2(\r_v0_x[9]_i_5_n_0 ),
        .I3(\u_geo/u_geo_tri/exp ),
        .I4(\r_v0_x[0]_i_5_n_0 ),
        .O(r_v0_x));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[0]_i_4 
       (.I0(\u_geo/w_vx_view [1]),
        .I1(\u_geo/u_geo_tri/w_set_y ),
        .I2(\u_geo/u_geo_tri/r_vy [1]),
        .O(\r_v0_x[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[0]_i_5 
       (.I0(\u_geo/w_vx_view [2]),
        .I1(\u_geo/u_geo_tri/w_set_y ),
        .I2(\u_geo/u_geo_tri/r_vy [2]),
        .O(\r_v0_x[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF088F0F0F0888888)) 
    \r_v0_x[10]_i_1 
       (.I0(\r_v0_x[10]_i_2_n_0 ),
        .I1(\r_v0_x[10]_i_3_n_0 ),
        .I2(\u_geo/u_geo_tri/w_ui_2c [11]),
        .I3(\u_geo/w_vx_view [21]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [21]),
        .O(\u_geo/u_geo_tri/p_0_in__0 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[10]_i_10 
       (.I0(\u_geo/w_vx_view [12]),
        .I1(\u_geo/u_geo_tri/r_vy [12]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [11]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [11]),
        .O(\r_v0_x[10]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[10]_i_11 
       (.I0(\u_geo/w_vx_view [14]),
        .I1(\u_geo/u_geo_tri/r_vy [14]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [13]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [13]),
        .O(\r_v0_x[10]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_v0_x[10]_i_2 
       (.I0(\r_v0_x[10]_i_4_n_0 ),
        .I1(\r_v0_x[10]_i_5_n_0 ),
        .O(\r_v0_x[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[10]_i_3 
       (.I0(\r_v0_x[10]_i_6_n_0 ),
        .I1(\r_v0_x[11]_i_9_n_0 ),
        .I2(\r_v0_x[10]_i_7_n_0 ),
        .O(\r_v0_x[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h77775FA088885FA0)) 
    \r_v0_x[10]_i_4 
       (.I0(\r_v0_x[10]_i_8_n_0 ),
        .I1(\u_geo/w_vx_view [18]),
        .I2(\u_geo/u_geo_tri/r_vy [18]),
        .I3(\u_geo/u_geo_tri/r_vy [19]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/w_vx_view [19]),
        .O(\r_v0_x[10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB88B744747474747)) 
    \r_v0_x[10]_i_5 
       (.I0(\u_geo/w_vx_view [20]),
        .I1(\u_geo/u_geo_tri/w_set_y ),
        .I2(\u_geo/u_geo_tri/r_vy [20]),
        .I3(\u_geo/u_geo_tri/r_vy [19]),
        .I4(\u_geo/w_vx_view [19]),
        .I5(\r_v0_x[10]_i_9_n_0 ),
        .O(\r_v0_x[10]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[10]_i_6 
       (.I0(\r_v0_x[10]_i_10_n_0 ),
        .I1(\r_v0_x[9]_i_5_n_0 ),
        .I2(\r_v0_x[10]_i_11_n_0 ),
        .O(\r_v0_x[10]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4703440000000000)) 
    \r_v0_x[10]_i_7 
       (.I0(\u_geo/w_vx_view [16]),
        .I1(\u_geo/u_geo_tri/w_set_y ),
        .I2(\u_geo/u_geo_tri/r_vy [16]),
        .I3(\u_geo/w_vx_view [15]),
        .I4(\u_geo/u_geo_tri/r_vy [15]),
        .I5(\r_v0_x[9]_i_5_n_0 ),
        .O(\r_v0_x[10]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCA000A0)) 
    \r_v0_x[10]_i_8 
       (.I0(\u_geo/u_geo_tri/r_vy [17]),
        .I1(\u_geo/w_vx_view [17]),
        .I2(\u_geo/u_geo_tri/r_vy [16]),
        .I3(\u_geo/u_geo_tri/w_set_y ),
        .I4(\u_geo/w_vx_view [16]),
        .O(\r_v0_x[10]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC000A0A0C0000000)) 
    \r_v0_x[10]_i_9 
       (.I0(\u_geo/u_geo_tri/r_vy [18]),
        .I1(\u_geo/w_vx_view [18]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [17]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [17]),
        .O(\r_v0_x[10]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBABF8A80)) 
    \r_v0_x[11]_i_1 
       (.I0(\u_geo/u_geo_tri/w_ui_2c [12]),
        .I1(\u_geo/w_vx_view [21]),
        .I2(\u_geo/u_geo_tri/w_set_y ),
        .I3(\u_geo/u_geo_tri/r_vy [21]),
        .I4(\u_geo/u_geo_tri/u_ftoi/f_ftoi__60 ),
        .O(\u_geo/u_geo_tri/p_0_in__0 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[11]_i_10 
       (.I0(\u_geo/w_vx_view [13]),
        .I1(\u_geo/u_geo_tri/r_vy [13]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [12]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [12]),
        .O(\r_v0_x[11]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[11]_i_11 
       (.I0(\u_geo/w_vx_view [16]),
        .I1(\u_geo/u_geo_tri/w_set_y ),
        .I2(\u_geo/u_geo_tri/r_vy [16]),
        .O(\u_geo/u_geo_tri/exp ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \r_v0_x[11]_i_3 
       (.I0(\r_v0_x[11]_i_8_n_0 ),
        .I1(\r_v0_x[11]_i_9_n_0 ),
        .I2(\r_v0_x[10]_i_2_n_0 ),
        .O(\u_geo/u_geo_tri/u_ftoi/f_ftoi__60 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \r_v0_x[11]_i_4 
       (.I0(\r_v0_x[10]_i_2_n_0 ),
        .I1(\r_v0_x[11]_i_9_n_0 ),
        .I2(\r_v0_x[11]_i_8_n_0 ),
        .O(\r_v0_x[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \r_v0_x[11]_i_5 
       (.I0(\r_v0_x[10]_i_2_n_0 ),
        .I1(\r_v0_x[10]_i_3_n_0 ),
        .O(\r_v0_x[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \r_v0_x[11]_i_6 
       (.I0(\r_v0_x[10]_i_2_n_0 ),
        .I1(\r_v0_x[9]_i_2_n_0 ),
        .O(\r_v0_x[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \r_v0_x[11]_i_7 
       (.I0(\r_v0_x[10]_i_2_n_0 ),
        .I1(\r_v0_x[8]_i_2_n_0 ),
        .O(\r_v0_x[11]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[11]_i_8 
       (.I0(\r_v0_x[11]_i_10_n_0 ),
        .I1(\r_v0_x[9]_i_5_n_0 ),
        .I2(\r_v0_x[9]_i_4_n_0 ),
        .O(\r_v0_x[11]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h77775FA088885FA0)) 
    \r_v0_x[11]_i_9 
       (.I0(\u_geo/u_geo_tri/exp ),
        .I1(\u_geo/w_vx_view [17]),
        .I2(\u_geo/u_geo_tri/r_vy [17]),
        .I3(\u_geo/u_geo_tri/r_vy [18]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/w_vx_view [18]),
        .O(\r_v0_x[11]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8A80BABF)) 
    \r_v0_x[1]_i_1 
       (.I0(\u_geo/u_geo_tri/w_ui_2c [2]),
        .I1(\u_geo/w_vx_view [21]),
        .I2(\u_geo/u_geo_tri/w_set_y ),
        .I3(\u_geo/u_geo_tri/r_vy [21]),
        .I4(\r_v0_x[3]_i_7_n_0 ),
        .O(\u_geo/u_geo_tri/p_0_in__0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT4 #(
    .INIT(16'hDDCF)) 
    \r_v0_x[1]_i_2 
       (.I0(\r_v0_x[1]_i_3_n_0 ),
        .I1(\r_v0_x[10]_i_5_n_0 ),
        .I2(\r_v0_x[9]_i_2_n_0 ),
        .I3(\r_v0_x[10]_i_4_n_0 ),
        .O(\r_v0_x[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFACA0ACA)) 
    \r_v0_x[1]_i_3 
       (.I0(\r_v0_x[5]_i_3_n_0 ),
        .I1(\r_v0_x[3]_i_11_n_0 ),
        .I2(\r_v0_x[11]_i_9_n_0 ),
        .I3(\r_v0_x[9]_i_5_n_0 ),
        .I4(\r_v0_x[1]_i_4_n_0 ),
        .O(\r_v0_x[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[1]_i_4 
       (.I0(\u_geo/w_vx_view [3]),
        .I1(\u_geo/u_geo_tri/r_vy [3]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [2]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [2]),
        .O(\r_v0_x[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8A80BABF)) 
    \r_v0_x[2]_i_1 
       (.I0(\u_geo/u_geo_tri/w_ui_2c [3]),
        .I1(\u_geo/w_vx_view [21]),
        .I2(\u_geo/u_geo_tri/w_set_y ),
        .I3(\u_geo/u_geo_tri/r_vy [21]),
        .I4(\r_v0_x[3]_i_6_n_0 ),
        .O(\u_geo/u_geo_tri/p_0_in__0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hDDCF)) 
    \r_v0_x[2]_i_2 
       (.I0(\r_v0_x[2]_i_3_n_0 ),
        .I1(\r_v0_x[10]_i_5_n_0 ),
        .I2(\r_v0_x[10]_i_3_n_0 ),
        .I3(\r_v0_x[10]_i_4_n_0 ),
        .O(\r_v0_x[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFACA0ACA)) 
    \r_v0_x[2]_i_3 
       (.I0(\r_v0_x[6]_i_3_n_0 ),
        .I1(\r_v0_x[4]_i_4_n_0 ),
        .I2(\r_v0_x[11]_i_9_n_0 ),
        .I3(\r_v0_x[9]_i_5_n_0 ),
        .I4(\r_v0_x[2]_i_4_n_0 ),
        .O(\r_v0_x[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[2]_i_4 
       (.I0(\u_geo/w_vx_view [4]),
        .I1(\u_geo/u_geo_tri/r_vy [4]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [3]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [3]),
        .O(\r_v0_x[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8A80BABF)) 
    \r_v0_x[3]_i_1 
       (.I0(\u_geo/u_geo_tri/w_ui_2c [4]),
        .I1(\u_geo/w_vx_view [21]),
        .I2(\u_geo/u_geo_tri/w_set_y ),
        .I3(\u_geo/u_geo_tri/r_vy [21]),
        .I4(\r_v0_x[3]_i_5_n_0 ),
        .O(\u_geo/u_geo_tri/p_0_in__0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0AACCAA)) 
    \r_v0_x[3]_i_10 
       (.I0(\r_v0_x[3]_i_9_n_0 ),
        .I1(\r_v0_x[1]_i_4_n_0 ),
        .I2(\r_v0_x[3]_i_12_n_0 ),
        .I3(\r_v0_x[11]_i_9_n_0 ),
        .I4(\r_v0_x[9]_i_5_n_0 ),
        .O(\r_v0_x[3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[3]_i_11 
       (.I0(\u_geo/w_vx_view [5]),
        .I1(\u_geo/u_geo_tri/r_vy [5]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [4]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [4]),
        .O(\r_v0_x[3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFC0CFAFAFC0C0A0A)) 
    \r_v0_x[3]_i_12 
       (.I0(\u_geo/u_geo_tri/r_vy [0]),
        .I1(\u_geo/w_vx_view [0]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [1]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [1]),
        .O(\r_v0_x[3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF193B5D7F)) 
    \r_v0_x[3]_i_3 
       (.I0(\r_v0_x[11]_i_9_n_0 ),
        .I1(\r_v0_x[10]_i_4_n_0 ),
        .I2(\r_v0_x[3]_i_9_n_0 ),
        .I3(\r_v0_x[11]_i_8_n_0 ),
        .I4(\r_v0_x[7]_i_4_n_0 ),
        .I5(\r_v0_x[10]_i_5_n_0 ),
        .O(\r_v0_x[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hAFBB)) 
    \r_v0_x[3]_i_4 
       (.I0(\r_v0_x[10]_i_5_n_0 ),
        .I1(\r_v0_x[7]_i_2_n_0 ),
        .I2(\r_v0_x[3]_i_10_n_0 ),
        .I3(\r_v0_x[10]_i_4_n_0 ),
        .O(\r_v0_x[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[3]_i_9 
       (.I0(\r_v0_x[3]_i_11_n_0 ),
        .I1(\r_v0_x[9]_i_5_n_0 ),
        .I2(\r_v0_x[5]_i_5_n_0 ),
        .O(\r_v0_x[3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8A80BABF)) 
    \r_v0_x[4]_i_1 
       (.I0(\u_geo/u_geo_tri/w_ui_2c [5]),
        .I1(\u_geo/w_vx_view [21]),
        .I2(\u_geo/u_geo_tri/w_set_y ),
        .I3(\u_geo/u_geo_tri/r_vy [21]),
        .I4(\r_v0_x[7]_i_8_n_0 ),
        .O(\u_geo/u_geo_tri/p_0_in__0 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF193B5D7F)) 
    \r_v0_x[4]_i_2 
       (.I0(\r_v0_x[11]_i_9_n_0 ),
        .I1(\r_v0_x[10]_i_4_n_0 ),
        .I2(\r_v0_x[4]_i_3_n_0 ),
        .I3(\r_v0_x[8]_i_4_n_0 ),
        .I4(\r_v0_x[8]_i_3_n_0 ),
        .I5(\r_v0_x[10]_i_5_n_0 ),
        .O(\r_v0_x[7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[4]_i_3 
       (.I0(\r_v0_x[4]_i_4_n_0 ),
        .I1(\r_v0_x[9]_i_5_n_0 ),
        .I2(\r_v0_x[6]_i_4_n_0 ),
        .O(\r_v0_x[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[4]_i_4 
       (.I0(\u_geo/w_vx_view [6]),
        .I1(\u_geo/u_geo_tri/r_vy [6]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [5]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [5]),
        .O(\r_v0_x[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8A80BABF)) 
    \r_v0_x[5]_i_1 
       (.I0(\u_geo/u_geo_tri/w_ui_2c [6]),
        .I1(\u_geo/w_vx_view [21]),
        .I2(\u_geo/u_geo_tri/w_set_y ),
        .I3(\u_geo/u_geo_tri/r_vy [21]),
        .I4(\r_v0_x[7]_i_7_n_0 ),
        .O(\u_geo/u_geo_tri/p_0_in__0 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF193B5D7F)) 
    \r_v0_x[5]_i_2 
       (.I0(\r_v0_x[11]_i_9_n_0 ),
        .I1(\r_v0_x[10]_i_4_n_0 ),
        .I2(\r_v0_x[5]_i_3_n_0 ),
        .I3(\r_v0_x[5]_i_4_n_0 ),
        .I4(\r_v0_x[9]_i_3_n_0 ),
        .I5(\r_v0_x[10]_i_5_n_0 ),
        .O(\r_v0_x[7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[5]_i_3 
       (.I0(\r_v0_x[5]_i_5_n_0 ),
        .I1(\r_v0_x[9]_i_5_n_0 ),
        .I2(\r_v0_x[7]_i_9_n_0 ),
        .O(\r_v0_x[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h202A808A2A208A80)) 
    \r_v0_x[5]_i_4 
       (.I0(\r_v0_x[9]_i_4_n_0 ),
        .I1(\u_geo/w_vx_view [17]),
        .I2(\u_geo/u_geo_tri/w_set_y ),
        .I3(\u_geo/u_geo_tri/r_vy [17]),
        .I4(\u_geo/w_vx_view [16]),
        .I5(\u_geo/u_geo_tri/r_vy [16]),
        .O(\r_v0_x[5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[5]_i_5 
       (.I0(\u_geo/w_vx_view [7]),
        .I1(\u_geo/u_geo_tri/r_vy [7]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [6]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [6]),
        .O(\r_v0_x[5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8A80BABF)) 
    \r_v0_x[6]_i_1 
       (.I0(\u_geo/u_geo_tri/w_ui_2c [7]),
        .I1(\u_geo/w_vx_view [21]),
        .I2(\u_geo/u_geo_tri/w_set_y ),
        .I3(\u_geo/u_geo_tri/r_vy [21]),
        .I4(\r_v0_x[7]_i_6_n_0 ),
        .O(\u_geo/u_geo_tri/p_0_in__0 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF193B5D7F)) 
    \r_v0_x[6]_i_2 
       (.I0(\r_v0_x[11]_i_9_n_0 ),
        .I1(\r_v0_x[10]_i_4_n_0 ),
        .I2(\r_v0_x[6]_i_3_n_0 ),
        .I3(\r_v0_x[10]_i_7_n_0 ),
        .I4(\r_v0_x[10]_i_6_n_0 ),
        .I5(\r_v0_x[10]_i_5_n_0 ),
        .O(\r_v0_x[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[6]_i_3 
       (.I0(\r_v0_x[6]_i_4_n_0 ),
        .I1(\r_v0_x[9]_i_5_n_0 ),
        .I2(\r_v0_x[8]_i_5_n_0 ),
        .O(\r_v0_x[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[6]_i_4 
       (.I0(\u_geo/w_vx_view [8]),
        .I1(\u_geo/u_geo_tri/r_vy [8]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [7]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [7]),
        .O(\r_v0_x[6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF088F0F0F0888888)) 
    \r_v0_x[7]_i_1 
       (.I0(\r_v0_x[10]_i_2_n_0 ),
        .I1(\r_v0_x[7]_i_2_n_0 ),
        .I2(\u_geo/u_geo_tri/w_ui_2c [8]),
        .I3(\u_geo/w_vx_view [21]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [21]),
        .O(\u_geo/u_geo_tri/p_0_in__0 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[7]_i_2 
       (.I0(\r_v0_x[7]_i_4_n_0 ),
        .I1(\r_v0_x[11]_i_9_n_0 ),
        .I2(\r_v0_x[11]_i_8_n_0 ),
        .O(\r_v0_x[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[7]_i_4 
       (.I0(\r_v0_x[7]_i_9_n_0 ),
        .I1(\r_v0_x[9]_i_5_n_0 ),
        .I2(\r_v0_x[9]_i_6_n_0 ),
        .O(\r_v0_x[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \r_v0_x[7]_i_5 
       (.I0(\r_v0_x[10]_i_2_n_0 ),
        .I1(\r_v0_x[7]_i_2_n_0 ),
        .O(\r_v0_x[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[7]_i_9 
       (.I0(\u_geo/w_vx_view [9]),
        .I1(\u_geo/u_geo_tri/r_vy [9]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [8]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [8]),
        .O(\r_v0_x[7]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF088F0F0F0888888)) 
    \r_v0_x[8]_i_1 
       (.I0(\r_v0_x[10]_i_2_n_0 ),
        .I1(\r_v0_x[8]_i_2_n_0 ),
        .I2(\u_geo/u_geo_tri/w_ui_2c [9]),
        .I3(\u_geo/w_vx_view [21]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [21]),
        .O(\u_geo/u_geo_tri/p_0_in__0 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[8]_i_2 
       (.I0(\r_v0_x[8]_i_3_n_0 ),
        .I1(\r_v0_x[11]_i_9_n_0 ),
        .I2(\r_v0_x[8]_i_4_n_0 ),
        .O(\r_v0_x[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[8]_i_3 
       (.I0(\r_v0_x[8]_i_5_n_0 ),
        .I1(\r_v0_x[9]_i_5_n_0 ),
        .I2(\r_v0_x[10]_i_10_n_0 ),
        .O(\r_v0_x[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888BBB888B8)) 
    \r_v0_x[8]_i_4 
       (.I0(\r_v0_x[10]_i_11_n_0 ),
        .I1(\r_v0_x[9]_i_5_n_0 ),
        .I2(\u_geo/u_geo_tri/r_vy [15]),
        .I3(\u_geo/u_geo_tri/w_set_y ),
        .I4(\u_geo/w_vx_view [15]),
        .I5(\u_geo/u_geo_tri/exp ),
        .O(\r_v0_x[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[8]_i_5 
       (.I0(\u_geo/w_vx_view [10]),
        .I1(\u_geo/u_geo_tri/r_vy [10]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [9]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [9]),
        .O(\r_v0_x[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF088F0F0F0888888)) 
    \r_v0_x[9]_i_1 
       (.I0(\r_v0_x[10]_i_2_n_0 ),
        .I1(\r_v0_x[9]_i_2_n_0 ),
        .I2(\u_geo/u_geo_tri/w_ui_2c [10]),
        .I3(\u_geo/w_vx_view [21]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [21]),
        .O(\u_geo/u_geo_tri/p_0_in__0 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB888)) 
    \r_v0_x[9]_i_2 
       (.I0(\r_v0_x[9]_i_3_n_0 ),
        .I1(\r_v0_x[11]_i_9_n_0 ),
        .I2(\r_v0_x[9]_i_4_n_0 ),
        .I3(\r_v0_x[9]_i_5_n_0 ),
        .O(\r_v0_x[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_v0_x[9]_i_3 
       (.I0(\r_v0_x[9]_i_6_n_0 ),
        .I1(\r_v0_x[9]_i_5_n_0 ),
        .I2(\r_v0_x[11]_i_10_n_0 ),
        .O(\r_v0_x[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[9]_i_4 
       (.I0(\u_geo/w_vx_view [15]),
        .I1(\u_geo/u_geo_tri/r_vy [15]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [14]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [14]),
        .O(\r_v0_x[9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h335ACC5A)) 
    \r_v0_x[9]_i_5 
       (.I0(\u_geo/u_geo_tri/r_vy [16]),
        .I1(\u_geo/w_vx_view [16]),
        .I2(\u_geo/u_geo_tri/r_vy [17]),
        .I3(\u_geo/u_geo_tri/w_set_y ),
        .I4(\u_geo/w_vx_view [17]),
        .O(\r_v0_x[9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \r_v0_x[9]_i_6 
       (.I0(\u_geo/w_vx_view [11]),
        .I1(\u_geo/u_geo_tri/r_vy [11]),
        .I2(\u_geo/u_geo_tri/exp ),
        .I3(\u_geo/w_vx_view [10]),
        .I4(\u_geo/u_geo_tri/w_set_y ),
        .I5(\u_geo/u_geo_tri/r_vy [10]),
        .O(\r_v0_x[9]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_v0_x_reg[11]_i_2 
       (.CI(\r_v0_x_reg[7]_i_3_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_tri/w_ui_2c [12:9]),
        .S({\r_v0_x[11]_i_4_n_0 ,\r_v0_x[11]_i_5_n_0 ,\r_v0_x[11]_i_6_n_0 ,\r_v0_x[11]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_v0_x_reg[3]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO(r_v0_x_reg),
        .CYINIT(\r_v0_x[3]_i_4_n_0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_tri/w_ui_2c [4:1]),
        .S({\r_v0_x[3]_i_5_n_0 ,\r_v0_x[3]_i_6_n_0 ,\r_v0_x[3]_i_7_n_0 ,\r_v0_x[3]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_v0_x_reg[7]_i_3 
       (.CI(r_v0_x_reg[3]),
        .CO({\r_v0_x_reg[7]_i_3_n_0 ,\r_v0_x_reg[7]_i_3_n_1 ,\r_v0_x_reg[7]_i_3_n_2 ,\r_v0_x_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_tri/w_ui_2c [8:5]),
        .S({\r_v0_x[7]_i_5_n_0 ,\r_v0_x[7]_i_6_n_0 ,\r_v0_x[7]_i_7_n_0 ,\r_v0_x[7]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h28AA000000000000)) 
    \r_v0_y[11]_i_1 
       (.I0(w_ack),
        .I1(\u_geo/u_geo_cull/p_0_in ),
        .I2(w_ccw),
        .I3(w_en_cull),
        .I4(\u_geo/u_geo_cull/r_state [0]),
        .I5(\u_geo/u_geo_cull/r_state [1]),
        .O(\u_ras/u_ras_state/w_set_vtx ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000008)) 
    \r_v1_outcode[5]_i_1 
       (.I0(\u_geo/u_geo_tri/p_0_in0_in ),
        .I1(\u_geo/u_geo_viewport/r_state [3]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_tri/w_set_v1_x ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000008)) 
    \r_v2_outcode[5]_i_1 
       (.I0(\u_geo/u_geo_tri/p_0_in ),
        .I1(\u_geo/u_geo_viewport/r_state [3]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [1]),
        .I4(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_tri/w_set_v2_x ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_vh[15]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[6]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[1]),
        .O(r_vh));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_vh[21]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[6]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[2]),
        .O(\r_vh[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r_vh[7]_i_1 
       (.I0(s_wb_adr_i[4]),
        .I1(s_wb_adr_i[6]),
        .I2(\r_dma_size[15]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[0]),
        .O(\r_vh[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_vw[15]_i_1 
       (.I0(s_wb_adr_i[6]),
        .I1(s_wb_adr_i[2]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[1]),
        .O(r_vw));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r_vw[21]_i_1 
       (.I0(\u_geo/w_en_mvp ),
        .I1(\u_geo/w_state_clip ),
        .O(\r_vw[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_vw[21]_i_1__0 
       (.I0(s_wb_adr_i[6]),
        .I1(s_wb_adr_i[2]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[2]),
        .O(\r_vw[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \r_vw[7]_i_1 
       (.I0(s_wb_adr_i[6]),
        .I1(s_wb_adr_i[2]),
        .I2(\r_m00[21]_i_2_n_0 ),
        .I3(s_wb_adr_i[5]),
        .I4(s_wb_adr_i[3]),
        .I5(s_wb_sel_i[0]),
        .O(\r_vw[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[0]_i_1 
       (.I0(\u_geo/w_vx_clip [0]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_ ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(r_vx));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[10]_i_1 
       (.I0(\u_geo/w_vx_clip [10]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[10] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[11]_i_1 
       (.I0(\u_geo/w_vx_clip [11]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[11] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[12]_i_1 
       (.I0(\u_geo/w_vx_clip [12]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[12] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[13]_i_1 
       (.I0(\u_geo/w_vx_clip [13]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[13] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[14]_i_1 
       (.I0(\u_geo/w_vx_clip [14]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[14] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFCCCDCCC)) 
    \r_vx[15]_i_1 
       (.I0(\r_vx[20]_i_2_n_0 ),
        .I1(m_wb_dat_i[30]),
        .I2(m_wb_dat_i[29]),
        .I3(m_wb_dat_i[28]),
        .I4(m_wb_dat_i[27]),
        .O(\u_geo/u_geo_mem/w_f22 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[15]_i_1__0 
       (.I0(\u_geo/w_vx_clip [15]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[15] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[15]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF80FF800000)) 
    \r_vx[16]_i_1 
       (.I0(m_wb_dat_i[27]),
        .I1(m_wb_dat_i[28]),
        .I2(m_wb_dat_i[29]),
        .I3(m_wb_dat_i[30]),
        .I4(\u_geo/u_geo_mem/p_0_in ),
        .I5(m_wb_dat_i[23]),
        .O(\u_geo/u_geo_mem/w_f22 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[16]_i_1__0 
       (.I0(\u_geo/w_vx_clip [16]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[16] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[16]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2A80)) 
    \r_vx[17]_i_1 
       (.I0(\r_vx[19]_i_2_n_0 ),
        .I1(m_wb_dat_i[23]),
        .I2(\u_geo/u_geo_mem/p_0_in ),
        .I3(m_wb_dat_i[24]),
        .O(\u_geo/u_geo_mem/w_f22 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[17]_i_1__0 
       (.I0(\u_geo/w_vx_clip [17]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[17] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[17]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h2AAA8000)) 
    \r_vx[18]_i_1 
       (.I0(\r_vx[19]_i_2_n_0 ),
        .I1(m_wb_dat_i[24]),
        .I2(\u_geo/u_geo_mem/p_0_in ),
        .I3(m_wb_dat_i[23]),
        .I4(m_wb_dat_i[25]),
        .O(\u_geo/u_geo_mem/w_f22 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[18]_i_1__0 
       (.I0(\u_geo/w_vx_clip [18]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[18] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[18]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7FFF000080000000)) 
    \r_vx[19]_i_1 
       (.I0(m_wb_dat_i[24]),
        .I1(\u_geo/u_geo_mem/p_0_in ),
        .I2(m_wb_dat_i[23]),
        .I3(m_wb_dat_i[25]),
        .I4(\r_vx[19]_i_2_n_0 ),
        .I5(m_wb_dat_i[26]),
        .O(\u_geo/u_geo_mem/w_f22 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[19]_i_1__0 
       (.I0(\u_geo/w_vx_clip [19]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[19] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[19]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF80)) 
    \r_vx[19]_i_2 
       (.I0(m_wb_dat_i[27]),
        .I1(m_wb_dat_i[28]),
        .I2(m_wb_dat_i[29]),
        .I3(m_wb_dat_i[30]),
        .O(\r_vx[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[1]_i_1 
       (.I0(\u_geo/w_vx_clip [1]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0F08F000)) 
    \r_vx[20]_i_1 
       (.I0(m_wb_dat_i[28]),
        .I1(m_wb_dat_i[29]),
        .I2(\r_vx[20]_i_2_n_0 ),
        .I3(m_wb_dat_i[30]),
        .I4(m_wb_dat_i[27]),
        .O(\u_geo/u_geo_mem/w_f22 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[20]_i_1__0 
       (.I0(\u_geo/w_vx_clip [20]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[20] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[20]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \r_vx[20]_i_2 
       (.I0(m_wb_dat_i[25]),
        .I1(m_wb_dat_i[23]),
        .I2(\u_geo/u_geo_mem/p_0_in ),
        .I3(m_wb_dat_i[24]),
        .I4(m_wb_dat_i[26]),
        .O(\r_vx[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB000)) 
    \r_vx[21]_i_1 
       (.I0(\u_mem_arb/r_req_geo ),
        .I1(\u_mem_arb/r_state ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I3(m_wb_ack_i),
        .O(\u_geo/u_geo_mem/r_vx ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h09)) 
    \r_vx[21]_i_1__0 
       (.I0(\u_geo/u_geo_persdiv/r_state [2]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .O(\r_vx[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0008)) 
    \r_vx[21]_i_1__1 
       (.I0(\u_geo/u_geo_viewport/r_state [1]),
        .I1(\u_geo/u_geo_viewport/r_state [2]),
        .I2(\u_geo/u_geo_viewport/r_state [3]),
        .I3(\u_geo/u_geo_viewport/r_state [0]),
        .O(\r_vx[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[21]_i_2 
       (.I0(\u_geo/w_vx_clip [21]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[21] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[2]_i_1 
       (.I0(\u_geo/w_vx_clip [2]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[2] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[3]_i_1 
       (.I0(\u_geo/w_vx_clip [3]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[3] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \r_vx[3]_i_5 
       (.I0(m_wb_dat_i[8]),
        .I1(m_wb_dat_i[7]),
        .O(\r_vx[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[4]_i_1 
       (.I0(\u_geo/w_vx_clip [4]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[4] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[5]_i_1 
       (.I0(\u_geo/w_vx_clip [5]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[5] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[6]_i_1 
       (.I0(\u_geo/w_vx_clip [6]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[6] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[7]_i_1 
       (.I0(\u_geo/w_vx_clip [7]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[7] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[8]_i_1 
       (.I0(\u_geo/w_vx_clip [8]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[8] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCCCCA)) 
    \r_vx[9]_i_1 
       (.I0(\u_geo/w_vx_clip [9]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[9] ),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [0]),
        .I4(\u_geo/u_geo_persdiv/r_state [2]),
        .O(\r_vx[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_vx_reg[11]_i_1 
       (.CI(\r_vx_reg[7]_i_1_n_0 ),
        .CO(r_vx_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_vx_reg[11]_i_1_n_4 ,\r_vx_reg[11]_i_1_n_5 ,\r_vx_reg[11]_i_1_n_6 ,\r_vx_reg[11]_i_1_n_7 }),
        .S(m_wb_dat_i[19:16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_vx_reg[14]_i_1 
       (.CI(r_vx_reg[3]),
        .CO({\u_geo/u_geo_mem/p_0_in ,\r_vx_reg[14]_i_1_n_1 ,\r_vx_reg[14]_i_1_n_2 ,\r_vx_reg[14]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_vx_reg[14]_i_1_n_4 ,\r_vx_reg[14]_i_1_n_5 ,\r_vx_reg[14]_i_1_n_6 ,\r_vx_reg[14]_i_1_n_7 }),
        .S({\<const1>__0__0 ,m_wb_dat_i[22:20]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_vx_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\r_vx_reg[3]_i_1_n_0 ,\r_vx_reg[3]_i_1_n_1 ,\r_vx_reg[3]_i_1_n_2 ,\r_vx_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,m_wb_dat_i[8]}),
        .O({\r_vx_reg[3]_i_1_n_4 ,\r_vx_reg[3]_i_1_n_5 ,\r_vx_reg[3]_i_1_n_6 ,\r_vx_reg[3]_i_1_n_7 }),
        .S({m_wb_dat_i[11:9],\r_vx[3]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_vx_reg[7]_i_1 
       (.CI(\r_vx_reg[3]_i_1_n_0 ),
        .CO({\r_vx_reg[7]_i_1_n_0 ,\r_vx_reg[7]_i_1_n_1 ,\r_vx_reg[7]_i_1_n_2 ,\r_vx_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_vx_reg[7]_i_1_n_4 ,\r_vx_reg[7]_i_1_n_5 ,\r_vx_reg[7]_i_1_n_6 ,\r_vx_reg[7]_i_1_n_7 }),
        .S(m_wb_dat_i[15:12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[0]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_ ),
        .I1(\u_geo/w_vy_clip [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(r_vy));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[10]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[10] ),
        .I1(\u_geo/w_vy_clip [10]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[11]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[11] ),
        .I1(\u_geo/w_vy_clip [11]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[12]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[12] ),
        .I1(\u_geo/w_vy_clip [12]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[13]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[13] ),
        .I1(\u_geo/w_vy_clip [13]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[14]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[14] ),
        .I1(\u_geo/w_vy_clip [14]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[15]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[15] ),
        .I1(\u_geo/w_vy_clip [15]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[16]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[16] ),
        .I1(\u_geo/w_vy_clip [16]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[17]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[17] ),
        .I1(\u_geo/w_vy_clip [17]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[18]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[18] ),
        .I1(\u_geo/w_vy_clip [18]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[19]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[19] ),
        .I1(\u_geo/w_vy_clip [19]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[1]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[1] ),
        .I1(\u_geo/w_vy_clip [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[20]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[20] ),
        .I1(\u_geo/w_vy_clip [20]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB000)) 
    \r_vy[21]_i_1 
       (.I0(\u_mem_arb/r_req_geo ),
        .I1(\u_mem_arb/r_state ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .I3(m_wb_ack_i),
        .O(\u_geo/u_geo_mem/r_vy ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h21)) 
    \r_vy[21]_i_1__0 
       (.I0(\u_geo/u_geo_persdiv/r_state [2]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .O(\r_vy[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0080)) 
    \r_vy[21]_i_1__1 
       (.I0(\u_geo/u_geo_viewport/r_state [0]),
        .I1(\u_geo/u_geo_viewport/r_state [1]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .O(\u_geo/u_geo_viewport/w_set_vy ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE00)) 
    \r_vy[21]_i_1__2 
       (.I0(\u_geo/w_state_if ),
        .I1(\u_geo/u_geo_tri/p_0_in ),
        .I2(\u_geo/u_geo_tri/p_0_in0_in ),
        .I3(\u_geo/w_en_view ),
        .O(\u_geo/u_geo_tri/w_set_y ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[21]_i_2 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[21] ),
        .I1(\u_geo/w_vy_clip [21]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[2]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[2] ),
        .I1(\u_geo/w_vy_clip [2]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[3]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[3] ),
        .I1(\u_geo/w_vy_clip [3]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[4]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[4] ),
        .I1(\u_geo/w_vy_clip [4]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[5]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[5] ),
        .I1(\u_geo/w_vy_clip [5]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[6]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[6] ),
        .I1(\u_geo/w_vy_clip [6]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[7]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[7] ),
        .I1(\u_geo/w_vy_clip [7]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[8]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[8] ),
        .I1(\u_geo/w_vy_clip [8]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCCCACCC)) 
    \r_vy[9]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[9] ),
        .I1(\u_geo/w_vy_clip [9]),
        .I2(\u_geo/u_geo_persdiv/r_state [2]),
        .I3(\u_geo/u_geo_persdiv/r_state [1]),
        .I4(\u_geo/u_geo_persdiv/r_state [0]),
        .O(\r_vy[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB000)) 
    \r_vz[21]_i_1 
       (.I0(\u_mem_arb/r_req_geo ),
        .I1(\u_mem_arb/r_state ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I3(m_wb_ack_i),
        .O(\u_geo/u_geo_mem/r_vz ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r_vz_in[21]_i_1 
       (.I0(\u_geo/w_state_mat ),
        .I1(\u_geo/w_en_dma ),
        .O(r_vz_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_x0_carry__0_i_1
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[7] ),
        .I1(\u_ras/u_ras_line/r_x_reg_n_0_[8] ),
        .O(r_x0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_x0_carry__0_i_2
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[6] ),
        .I1(\u_ras/u_ras_line/r_x_reg_n_0_[7] ),
        .O(r_x0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_x0_carry__0_i_3
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[5] ),
        .I1(\u_ras/u_ras_line/r_x_reg_n_0_[6] ),
        .O(r_x0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_x0_carry__0_i_4
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[4] ),
        .I1(\u_ras/u_ras_line/r_x_reg_n_0_[5] ),
        .O(r_x0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_x0_carry__1_i_1
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[10] ),
        .I1(\u_ras/w_x ),
        .O(r_x0_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_x0_carry__1_i_2
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[9] ),
        .I1(\u_ras/u_ras_line/r_x_reg_n_0_[10] ),
        .O(r_x0_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_x0_carry__1_i_3
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[8] ),
        .I1(\u_ras/u_ras_line/r_x_reg_n_0_[9] ),
        .O(r_x0_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    r_x0_carry_i_1
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[1] ),
        .O(r_x0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_x0_carry_i_2
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[3] ),
        .I1(\u_ras/u_ras_line/r_x_reg_n_0_[4] ),
        .O(r_x0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_x0_carry_i_3
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[2] ),
        .I1(\u_ras/u_ras_line/r_x_reg_n_0_[3] ),
        .O(r_x0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_x0_carry_i_4
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[1] ),
        .I1(\u_ras/u_ras_line/r_x_reg_n_0_[2] ),
        .O(r_x0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA9A9A9A95959A959)) 
    r_x0_carry_i_5
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[1] ),
        .I1(r_x0_carry_i_6_n_0),
        .I2(r_y0_carry_i_7_n_0),
        .I3(\u_ras/u_ras_line/w_sx_flag1__5 ),
        .I4(\u_ras/u_ras_line/r_x1 [11]),
        .I5(\u_ras/u_ras_line/r_x0 [11]),
        .O(r_x0_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFD79AF7BFD58AD08)) 
    r_x0_carry_i_6
       (.I0(\u_ras/u_ras_state/r_state [0]),
        .I1(\u_ras/u_ras_state/p_0_in ),
        .I2(\u_ras/u_ras_state/r_state [1]),
        .I3(\u_ras/u_ras_state/p_1_in ),
        .I4(\u_ras/u_ras_state/p_1_in8_in ),
        .I5(\u_ras/u_ras_line/w_sx_flag1__5 ),
        .O(r_x0_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    \r_x[0]_i_1 
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_ ),
        .I1(\u_ras/w_v0_x [0]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(r_x));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_x[10]_i_1 
       (.I0(\u_ras_line/r_x0_carry__1_n_6 ),
        .I1(\u_ras/w_v0_x [10]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_x[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5055004455555555)) 
    \r_x[11]_i_1 
       (.I0(\u_ras/u_ras_line/r_state_reg_n_0_ ),
        .I1(r_x_reg[1]),
        .I2(\u_ras/u_ras_line/result0_carry__0_n_2 ),
        .I3(\u_ras/u_ras_line/r_e2 ),
        .I4(\u_ras/u_ras_line/w_dym__22 ),
        .I5(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\u_ras/u_ras_line/r_x ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \r_x[11]_i_10 
       (.I0(\u_ras/r_e2 [4]),
        .I1(\u_ras/u_ras_line/w_dym_carry__0_n_7 ),
        .I2(\u_ras/u_ras_line/w_dym_carry__0_n_6 ),
        .I3(\u_ras/r_e2 [5]),
        .O(\r_x[11]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \r_x[11]_i_11 
       (.I0(\u_ras/r_e2 [2]),
        .I1(\u_ras/u_ras_line/w_dym_carry_n_5 ),
        .I2(\u_ras/u_ras_line/w_dym_carry_n_4 ),
        .I3(\u_ras/r_e2 [3]),
        .O(\r_x[11]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_x[11]_i_12 
       (.I0(\u_ras/r_e2 [1]),
        .I1(\u_ras/u_ras_line/w_dym_carry_n_6 ),
        .O(\r_x[11]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r_x[11]_i_13 
       (.I0(\u_ras/r_e2 [6]),
        .I1(\u_ras/u_ras_line/w_dym_carry__0_n_5 ),
        .I2(\u_ras/r_e2 [7]),
        .I3(\u_ras/u_ras_line/w_dym_carry__0_n_4 ),
        .O(\r_x[11]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r_x[11]_i_14 
       (.I0(\u_ras/r_e2 [4]),
        .I1(\u_ras/u_ras_line/w_dym_carry__0_n_7 ),
        .I2(\u_ras/r_e2 [5]),
        .I3(\u_ras/u_ras_line/w_dym_carry__0_n_6 ),
        .O(\r_x[11]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r_x[11]_i_15 
       (.I0(\u_ras/r_e2 [2]),
        .I1(\u_ras/u_ras_line/w_dym_carry_n_5 ),
        .I2(\u_ras/r_e2 [3]),
        .I3(\u_ras/u_ras_line/w_dym_carry_n_4 ),
        .O(\r_x[11]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h09)) 
    \r_x[11]_i_16 
       (.I0(\u_ras/r_e2 [1]),
        .I1(\u_ras/u_ras_line/w_dym_carry_n_6 ),
        .I2(\u_ras/u_ras_line/w_dym_carry_n_7 ),
        .O(\r_x[11]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_x[11]_i_2 
       (.I0(\u_ras_line/r_x0_carry__1_n_5 ),
        .I1(\u_ras/w_v0_x [11]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_x[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_x[11]_i_5 
       (.I0(\u_ras/r_e2 [10]),
        .I1(\u_ras/u_ras_line/w_dym_carry__1_n_5 ),
        .O(\r_x[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \r_x[11]_i_6 
       (.I0(\u_ras/r_e2 [8]),
        .I1(\u_ras/u_ras_line/w_dym_carry__1_n_7 ),
        .I2(\u_ras/u_ras_line/w_dym_carry__1_n_6 ),
        .I3(\u_ras/r_e2 [9]),
        .O(\r_x[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r_x[11]_i_7 
       (.I0(\u_ras/u_ras_line/w_dym_carry__1_n_5 ),
        .I1(\u_ras/r_e2 [10]),
        .O(\r_x[11]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \r_x[11]_i_8 
       (.I0(\u_ras/r_e2 [8]),
        .I1(\u_ras/u_ras_line/w_dym_carry__1_n_7 ),
        .I2(\u_ras/r_e2 [9]),
        .I3(\u_ras/u_ras_line/w_dym_carry__1_n_6 ),
        .O(\r_x[11]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \r_x[11]_i_9 
       (.I0(\u_ras/r_e2 [6]),
        .I1(\u_ras/u_ras_line/w_dym_carry__0_n_5 ),
        .I2(\u_ras/u_ras_line/w_dym_carry__0_n_4 ),
        .I3(\u_ras/r_e2 [7]),
        .O(\r_x[11]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_x[1]_i_1 
       (.I0(\u_ras_line/r_x0_carry_n_7 ),
        .I1(\u_ras/w_v0_x [1]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_x[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_x[2]_i_1 
       (.I0(\u_ras_line/r_x0_carry_n_6 ),
        .I1(\u_ras/w_v0_x [2]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_x[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_x[3]_i_1 
       (.I0(\u_ras_line/r_x0_carry_n_5 ),
        .I1(\u_ras/w_v0_x [3]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_x[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_x[4]_i_1 
       (.I0(\u_ras_line/r_x0_carry_n_4 ),
        .I1(\u_ras/w_v0_x [4]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_x[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_x[5]_i_1 
       (.I0(\u_ras_line/r_x0_carry__0_n_7 ),
        .I1(\u_ras/w_v0_x [5]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_x[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_x[6]_i_1 
       (.I0(\u_ras_line/r_x0_carry__0_n_6 ),
        .I1(\u_ras/w_v0_x [6]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_x[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_x[7]_i_1 
       (.I0(\u_ras_line/r_x0_carry__0_n_5 ),
        .I1(\u_ras/w_v0_x [7]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_x[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_x[8]_i_1 
       (.I0(\u_ras_line/r_x0_carry__0_n_4 ),
        .I1(\u_ras/w_v0_x [8]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_x[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_x[9]_i_1 
       (.I0(\u_ras_line/r_x0_carry__1_n_7 ),
        .I1(\u_ras/w_v0_x [9]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_x[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_x_reg[11]_i_3 
       (.CI(\r_x_reg[11]_i_4_n_0 ),
        .CO(r_x_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r_x[11]_i_5_n_0 ,\r_x[11]_i_6_n_0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\r_x[11]_i_7_n_0 ,\r_x[11]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \r_x_reg[11]_i_4 
       (.CI(\<const0>__0__0 ),
        .CO({\r_x_reg[11]_i_4_n_0 ,\r_x_reg[11]_i_4_n_1 ,\r_x_reg[11]_i_4_n_2 ,\r_x_reg[11]_i_4_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\r_x[11]_i_9_n_0 ,\r_x[11]_i_10_n_0 ,\r_x[11]_i_11_n_0 ,\r_x[11]_i_12_n_0 }),
        .S({\r_x[11]_i_13_n_0 ,\r_x[11]_i_14_n_0 ,\r_x[11]_i_15_n_0 ,\r_x[11]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_y0_carry__0_i_1
       (.I0(\u_ras/r_y [7]),
        .I1(\u_ras/r_y [8]),
        .O(r_y0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_y0_carry__0_i_2
       (.I0(\u_ras/r_y [6]),
        .I1(\u_ras/r_y [7]),
        .O(r_y0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_y0_carry__0_i_3
       (.I0(\u_ras/r_y [5]),
        .I1(\u_ras/r_y [6]),
        .O(r_y0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_y0_carry__0_i_4
       (.I0(\u_ras/r_y [4]),
        .I1(\u_ras/r_y [5]),
        .O(r_y0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_y0_carry__1_i_1
       (.I0(\u_ras/r_y [10]),
        .I1(\u_ras/w_y ),
        .O(r_y0_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_y0_carry__1_i_2
       (.I0(\u_ras/r_y [9]),
        .I1(\u_ras/r_y [10]),
        .O(r_y0_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_y0_carry__1_i_3
       (.I0(\u_ras/r_y [8]),
        .I1(\u_ras/r_y [9]),
        .O(r_y0_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    r_y0_carry_i_1
       (.I0(\u_ras/r_y [1]),
        .O(r_y0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_y0_carry_i_2
       (.I0(\u_ras/r_y [3]),
        .I1(\u_ras/r_y [4]),
        .O(r_y0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_y0_carry_i_3
       (.I0(\u_ras/r_y [2]),
        .I1(\u_ras/r_y [3]),
        .O(r_y0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    r_y0_carry_i_4
       (.I0(\u_ras/r_y [1]),
        .I1(\u_ras/r_y [2]),
        .O(r_y0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA9A9A9A95959A959)) 
    r_y0_carry_i_5
       (.I0(\u_ras/r_y [1]),
        .I1(r_y0_carry_i_6_n_0),
        .I2(r_y0_carry_i_7_n_0),
        .I3(\u_ras/u_ras_line/w_sy_flag1__5 ),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[11] ),
        .I5(\u_ras/u_ras_line/r_y0 [11]),
        .O(r_y0_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFD79AF7BFD58AD08)) 
    r_y0_carry_i_6
       (.I0(\u_ras/u_ras_state/r_state [0]),
        .I1(\u_ras/u_ras_state/p_0_in0_in ),
        .I2(\u_ras/u_ras_state/r_state [1]),
        .I3(\u_ras/u_ras_state/p_1_in1_in ),
        .I4(\u_ras/u_ras_state/p_1_in10_in ),
        .I5(\u_ras/u_ras_line/w_sy_flag1__5 ),
        .O(r_y0_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    r_y0_carry_i_7
       (.I0(\u_ras/u_ras_line/r_state_reg_n_0_ ),
        .I1(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(r_y0_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r_y1[11]_i_1 
       (.I0(\u_ras/u_ras_line/r_state_reg_n_0_ ),
        .I1(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\u_ras/u_ras_line/r_y1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    \r_y[0]_i_1 
       (.I0(\u_ras/r_y [0]),
        .I1(\u_ras/w_v0_y [0]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(r_y));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_y[10]_i_1 
       (.I0(\u_ras_line/r_y0_carry__1_n_6 ),
        .I1(\u_ras/w_v0_y [10]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_y[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45045555)) 
    \r_y[11]_i_1 
       (.I0(\u_ras/u_ras_line/r_state_reg_n_0_ ),
        .I1(\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ),
        .I2(\u_ras/u_ras_line/w_dx ),
        .I3(\u_ras/u_ras_line/r_e2 ),
        .I4(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\u_ras/u_ras_line/r_y ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_y[11]_i_2 
       (.I0(\u_ras_line/r_y0_carry__1_n_5 ),
        .I1(\u_ras/w_v0_y [11]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_y[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_y[1]_i_1 
       (.I0(\u_ras_line/r_y0_carry_n_7 ),
        .I1(\u_ras/w_v0_y [1]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_y[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_y[2]_i_1 
       (.I0(\u_ras_line/r_y0_carry_n_6 ),
        .I1(\u_ras/w_v0_y [2]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_y[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_y[3]_i_1 
       (.I0(\u_ras_line/r_y0_carry_n_5 ),
        .I1(\u_ras/w_v0_y [3]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_y[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_y[4]_i_1 
       (.I0(\u_ras_line/r_y0_carry_n_4 ),
        .I1(\u_ras/w_v0_y [4]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_y[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_y[5]_i_1 
       (.I0(\u_ras_line/r_y0_carry__0_n_7 ),
        .I1(\u_ras/w_v0_y [5]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_y[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_y[6]_i_1 
       (.I0(\u_ras_line/r_y0_carry__0_n_6 ),
        .I1(\u_ras/w_v0_y [6]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_y[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_y[7]_i_1 
       (.I0(\u_ras_line/r_y0_carry__0_n_5 ),
        .I1(\u_ras/w_v0_y [7]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_y[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_y[8]_i_1 
       (.I0(\u_ras_line/r_y0_carry__0_n_4 ),
        .I1(\u_ras/w_v0_y [8]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_y[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_y[9]_i_1 
       (.I0(\u_ras_line/r_y0_carry__1_n_7 ),
        .I1(\u_ras/w_v0_y [9]),
        .I2(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\r_y[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBF80)) 
    r_y_flip_i_1
       (.I0(s_wb_dat_i[8]),
        .I1(s_wb_sel_i[1]),
        .I2(\u_sys/w_hit1A_w__2 ),
        .I3(w_y_flip),
        .O(r_y_flip_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    r_y_flip_i_2
       (.I0(s_wb_adr_i[2]),
        .I1(s_wb_adr_i[4]),
        .I2(s_wb_adr_i[6]),
        .I3(\r_m10[21]_i_3_n_0 ),
        .I4(s_wb_adr_i[5]),
        .I5(s_wb_adr_i[3]),
        .O(\u_sys/w_hit1A_w__2 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result0_carry__0_i_1
       (.I0(\u_ras/r_e2 [10]),
        .I1(\u_ras/u_ras_line/w_dym_carry__1_n_5 ),
        .I2(\u_ras/u_ras_line/w_dym__22 ),
        .I3(\u_ras/u_ras_line/r_e2 ),
        .O(result0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result0_carry__0_i_2
       (.I0(\u_ras/r_e2 [8]),
        .I1(\u_ras/u_ras_line/w_dym_carry__1_n_7 ),
        .I2(\u_ras/u_ras_line/w_dym_carry__1_n_6 ),
        .I3(\u_ras/r_e2 [9]),
        .O(result0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result0_carry__0_i_3
       (.I0(\u_ras/r_e2 [10]),
        .I1(\u_ras/u_ras_line/w_dym_carry__1_n_5 ),
        .I2(\u_ras/u_ras_line/r_e2 ),
        .I3(\u_ras/u_ras_line/w_dym__22 ),
        .O(result0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result0_carry__0_i_4
       (.I0(\u_ras/r_e2 [8]),
        .I1(\u_ras/u_ras_line/w_dym_carry__1_n_7 ),
        .I2(\u_ras/r_e2 [9]),
        .I3(\u_ras/u_ras_line/w_dym_carry__1_n_6 ),
        .O(result0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result0_carry_i_1
       (.I0(\u_ras/r_e2 [6]),
        .I1(\u_ras/u_ras_line/w_dym_carry__0_n_5 ),
        .I2(\u_ras/u_ras_line/w_dym_carry__0_n_4 ),
        .I3(\u_ras/r_e2 [7]),
        .O(result0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result0_carry_i_2
       (.I0(\u_ras/r_e2 [4]),
        .I1(\u_ras/u_ras_line/w_dym_carry__0_n_7 ),
        .I2(\u_ras/u_ras_line/w_dym_carry__0_n_6 ),
        .I3(\u_ras/r_e2 [5]),
        .O(result0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result0_carry_i_3
       (.I0(\u_ras/r_e2 [2]),
        .I1(\u_ras/u_ras_line/w_dym_carry_n_5 ),
        .I2(\u_ras/u_ras_line/w_dym_carry_n_4 ),
        .I3(\u_ras/r_e2 [3]),
        .O(result0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    result0_carry_i_4
       (.I0(\u_ras/r_e2 [1]),
        .I1(\u_ras/u_ras_line/w_dym_carry_n_6 ),
        .O(result0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result0_carry_i_5
       (.I0(\u_ras/r_e2 [6]),
        .I1(\u_ras/u_ras_line/w_dym_carry__0_n_5 ),
        .I2(\u_ras/r_e2 [7]),
        .I3(\u_ras/u_ras_line/w_dym_carry__0_n_4 ),
        .O(result0_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result0_carry_i_6
       (.I0(\u_ras/r_e2 [4]),
        .I1(\u_ras/u_ras_line/w_dym_carry__0_n_7 ),
        .I2(\u_ras/r_e2 [5]),
        .I3(\u_ras/u_ras_line/w_dym_carry__0_n_6 ),
        .O(result0_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result0_carry_i_7
       (.I0(\u_ras/r_e2 [2]),
        .I1(\u_ras/u_ras_line/w_dym_carry_n_5 ),
        .I2(\u_ras/r_e2 [3]),
        .I3(\u_ras/u_ras_line/w_dym_carry_n_4 ),
        .O(result0_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h09)) 
    result0_carry_i_8
       (.I0(\u_ras/r_e2 [1]),
        .I1(\u_ras/u_ras_line/w_dym_carry_n_6 ),
        .I2(\u_ras/u_ras_line/w_dym_carry_n_7 ),
        .O(result0_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result0_inferred__1_carry__0_i_1
       (.I0(\u_ras/u_ras_line/_inferred__5_carry__1_n_5 ),
        .I1(\u_ras/r_e2 [10]),
        .I2(\u_ras/u_ras_line/r_e2 ),
        .I3(\u_ras/u_ras_line/w_dx ),
        .O(result0_inferred__1_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result0_inferred__1_carry__0_i_2
       (.I0(\u_ras/u_ras_line/_inferred__5_carry__1_n_7 ),
        .I1(\u_ras/r_e2 [8]),
        .I2(\u_ras/r_e2 [9]),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__1_n_6 ),
        .O(result0_inferred__1_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result0_inferred__1_carry__0_i_3
       (.I0(\u_ras/u_ras_line/_inferred__5_carry__1_n_5 ),
        .I1(\u_ras/r_e2 [10]),
        .I2(\u_ras/u_ras_line/w_dx ),
        .I3(\u_ras/u_ras_line/r_e2 ),
        .O(result0_inferred__1_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result0_inferred__1_carry__0_i_4
       (.I0(\u_ras/u_ras_line/_inferred__5_carry__1_n_7 ),
        .I1(\u_ras/r_e2 [8]),
        .I2(\u_ras/u_ras_line/_inferred__5_carry__1_n_6 ),
        .I3(\u_ras/r_e2 [9]),
        .O(result0_inferred__1_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result0_inferred__1_carry_i_1
       (.I0(\u_ras/u_ras_line/_inferred__5_carry__0_n_5 ),
        .I1(\u_ras/r_e2 [6]),
        .I2(\u_ras/r_e2 [7]),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__0_n_4 ),
        .O(result0_inferred__1_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result0_inferred__1_carry_i_2
       (.I0(\u_ras/u_ras_line/_inferred__5_carry__0_n_7 ),
        .I1(\u_ras/r_e2 [4]),
        .I2(\u_ras/r_e2 [5]),
        .I3(\u_ras/u_ras_line/_inferred__5_carry__0_n_6 ),
        .O(result0_inferred__1_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result0_inferred__1_carry_i_3
       (.I0(\u_ras/u_ras_line/_inferred__5_carry_n_5 ),
        .I1(\u_ras/r_e2 [2]),
        .I2(\u_ras/r_e2 [3]),
        .I3(\u_ras/u_ras_line/_inferred__5_carry_n_4 ),
        .O(result0_inferred__1_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB2)) 
    result0_inferred__1_carry_i_4
       (.I0(\u_ras/u_ras_line/_inferred__5_carry_n_7 ),
        .I1(\u_ras/r_e2 [1]),
        .I2(\u_ras/u_ras_line/_inferred__5_carry_n_6 ),
        .O(result0_inferred__1_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result0_inferred__1_carry_i_5
       (.I0(\u_ras/u_ras_line/_inferred__5_carry__0_n_5 ),
        .I1(\u_ras/r_e2 [6]),
        .I2(\u_ras/u_ras_line/_inferred__5_carry__0_n_4 ),
        .I3(\u_ras/r_e2 [7]),
        .O(result0_inferred__1_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result0_inferred__1_carry_i_6
       (.I0(\u_ras/u_ras_line/_inferred__5_carry__0_n_7 ),
        .I1(\u_ras/r_e2 [4]),
        .I2(\u_ras/u_ras_line/_inferred__5_carry__0_n_6 ),
        .I3(\u_ras/r_e2 [5]),
        .O(result0_inferred__1_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result0_inferred__1_carry_i_7
       (.I0(\u_ras/u_ras_line/_inferred__5_carry_n_5 ),
        .I1(\u_ras/r_e2 [2]),
        .I2(\u_ras/u_ras_line/_inferred__5_carry_n_4 ),
        .I3(\u_ras/r_e2 [3]),
        .O(result0_inferred__1_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h09)) 
    result0_inferred__1_carry_i_8
       (.I0(\u_ras/u_ras_line/_inferred__5_carry_n_6 ),
        .I1(\u_ras/r_e2 [1]),
        .I2(\u_ras/u_ras_line/_inferred__5_carry_n_7 ),
        .O(result0_inferred__1_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    result3_carry__0_i_1
       (.I0(w_scr_w_m1[10]),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_[10] ),
        .I2(w_scr_w_m1[11]),
        .O(result3_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_carry__0_i_2
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[8] ),
        .I1(w_scr_w_m1[8]),
        .I2(w_scr_w_m1[9]),
        .I3(\u_ras/u_ras_state/r_v1_x_reg_n_0_[9] ),
        .O(result3_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    result3_carry__0_i_3
       (.I0(w_scr_w_m1[14]),
        .I1(w_scr_w_m1[15]),
        .O(result3_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    result3_carry__0_i_4
       (.I0(w_scr_w_m1[12]),
        .I1(w_scr_w_m1[13]),
        .O(result3_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h09)) 
    result3_carry__0_i_5
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[10] ),
        .I1(w_scr_w_m1[10]),
        .I2(w_scr_w_m1[11]),
        .O(result3_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_carry__0_i_6
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[8] ),
        .I1(w_scr_w_m1[8]),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[9] ),
        .I3(w_scr_w_m1[9]),
        .O(result3_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_carry_i_1
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[6] ),
        .I1(w_scr_w_m1[6]),
        .I2(w_scr_w_m1[7]),
        .I3(\u_ras/u_ras_state/r_v1_x_reg_n_0_[7] ),
        .O(result3_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_carry_i_2
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[4] ),
        .I1(w_scr_w_m1[4]),
        .I2(w_scr_w_m1[5]),
        .I3(\u_ras/u_ras_state/r_v1_x_reg_n_0_[5] ),
        .O(result3_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_carry_i_3
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[2] ),
        .I1(w_scr_w_m1[2]),
        .I2(w_scr_w_m1[3]),
        .I3(\u_ras/u_ras_state/r_v1_x_reg_n_0_[3] ),
        .O(result3_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_carry_i_4
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_ ),
        .I1(w_scr_w_m1[0]),
        .I2(w_scr_w_m1[1]),
        .I3(\u_ras/u_ras_state/r_v1_x_reg_n_0_[1] ),
        .O(result3_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_carry_i_5
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[6] ),
        .I1(w_scr_w_m1[6]),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[7] ),
        .I3(w_scr_w_m1[7]),
        .O(result3_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_carry_i_6
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[4] ),
        .I1(w_scr_w_m1[4]),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[5] ),
        .I3(w_scr_w_m1[5]),
        .O(result3_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_carry_i_7
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[2] ),
        .I1(w_scr_w_m1[2]),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[3] ),
        .I3(w_scr_w_m1[3]),
        .O(result3_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_carry_i_8
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_ ),
        .I1(w_scr_w_m1[0]),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[1] ),
        .I3(w_scr_w_m1[1]),
        .O(result3_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    result3_inferred__0_carry__0_i_1
       (.I0(w_scr_w_m1[10]),
        .I1(\u_ras/u_ras_state/r_v0_x_reg_n_0_[10] ),
        .I2(w_scr_w_m1[11]),
        .O(result3_inferred__0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__0_carry__0_i_2
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[8] ),
        .I1(w_scr_w_m1[8]),
        .I2(w_scr_w_m1[9]),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[9] ),
        .O(result3_inferred__0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    result3_inferred__0_carry__0_i_3
       (.I0(w_scr_w_m1[14]),
        .I1(w_scr_w_m1[15]),
        .O(result3_inferred__0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    result3_inferred__0_carry__0_i_4
       (.I0(w_scr_w_m1[12]),
        .I1(w_scr_w_m1[13]),
        .O(result3_inferred__0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h09)) 
    result3_inferred__0_carry__0_i_5
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[10] ),
        .I1(w_scr_w_m1[10]),
        .I2(w_scr_w_m1[11]),
        .O(result3_inferred__0_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__0_carry__0_i_6
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[8] ),
        .I1(w_scr_w_m1[8]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[9] ),
        .I3(w_scr_w_m1[9]),
        .O(result3_inferred__0_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__0_carry_i_1
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[6] ),
        .I1(w_scr_w_m1[6]),
        .I2(w_scr_w_m1[7]),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[7] ),
        .O(result3_inferred__0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__0_carry_i_2
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[4] ),
        .I1(w_scr_w_m1[4]),
        .I2(w_scr_w_m1[5]),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[5] ),
        .O(result3_inferred__0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__0_carry_i_3
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[2] ),
        .I1(w_scr_w_m1[2]),
        .I2(w_scr_w_m1[3]),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[3] ),
        .O(result3_inferred__0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__0_carry_i_4
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_ ),
        .I1(w_scr_w_m1[0]),
        .I2(w_scr_w_m1[1]),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[1] ),
        .O(result3_inferred__0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__0_carry_i_5
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[6] ),
        .I1(w_scr_w_m1[6]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[7] ),
        .I3(w_scr_w_m1[7]),
        .O(result3_inferred__0_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__0_carry_i_6
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[4] ),
        .I1(w_scr_w_m1[4]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[5] ),
        .I3(w_scr_w_m1[5]),
        .O(result3_inferred__0_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__0_carry_i_7
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[2] ),
        .I1(w_scr_w_m1[2]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[3] ),
        .I3(w_scr_w_m1[3]),
        .O(result3_inferred__0_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__0_carry_i_8
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_ ),
        .I1(w_scr_w_m1[0]),
        .I2(\u_ras/u_ras_state/r_v0_x_reg_n_0_[1] ),
        .I3(w_scr_w_m1[1]),
        .O(result3_inferred__0_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    result3_inferred__1_carry__0_i_1
       (.I0(w_scr_h_m1[10]),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[10] ),
        .I2(w_scr_h_m1[11]),
        .O(result3_inferred__1_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__1_carry__0_i_2
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[8] ),
        .I1(w_scr_h_m1[8]),
        .I2(w_scr_h_m1[9]),
        .I3(\u_ras/u_ras_state/r_v1_y_reg_n_0_[9] ),
        .O(result3_inferred__1_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    result3_inferred__1_carry__0_i_3
       (.I0(w_scr_h_m1[14]),
        .I1(w_scr_h_m1[15]),
        .O(result3_inferred__1_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    result3_inferred__1_carry__0_i_4
       (.I0(w_scr_h_m1[12]),
        .I1(w_scr_h_m1[13]),
        .O(result3_inferred__1_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h09)) 
    result3_inferred__1_carry__0_i_5
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[10] ),
        .I1(w_scr_h_m1[10]),
        .I2(w_scr_h_m1[11]),
        .O(result3_inferred__1_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__1_carry__0_i_6
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[8] ),
        .I1(w_scr_h_m1[8]),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[9] ),
        .I3(w_scr_h_m1[9]),
        .O(result3_inferred__1_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__1_carry_i_1
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[6] ),
        .I1(w_scr_h_m1[6]),
        .I2(w_scr_h_m1[7]),
        .I3(\u_ras/u_ras_state/r_v1_y_reg_n_0_[7] ),
        .O(result3_inferred__1_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__1_carry_i_2
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[4] ),
        .I1(w_scr_h_m1[4]),
        .I2(w_scr_h_m1[5]),
        .I3(\u_ras/u_ras_state/r_v1_y_reg_n_0_[5] ),
        .O(result3_inferred__1_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__1_carry_i_3
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[2] ),
        .I1(w_scr_h_m1[2]),
        .I2(w_scr_h_m1[3]),
        .I3(\u_ras/u_ras_state/r_v1_y_reg_n_0_[3] ),
        .O(result3_inferred__1_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__1_carry_i_4
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_ ),
        .I1(w_scr_h_m1[0]),
        .I2(w_scr_h_m1[1]),
        .I3(\u_ras/u_ras_state/r_v1_y_reg_n_0_[1] ),
        .O(result3_inferred__1_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__1_carry_i_5
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[6] ),
        .I1(w_scr_h_m1[6]),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[7] ),
        .I3(w_scr_h_m1[7]),
        .O(result3_inferred__1_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__1_carry_i_6
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[4] ),
        .I1(w_scr_h_m1[4]),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[5] ),
        .I3(w_scr_h_m1[5]),
        .O(result3_inferred__1_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__1_carry_i_7
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[2] ),
        .I1(w_scr_h_m1[2]),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[3] ),
        .I3(w_scr_h_m1[3]),
        .O(result3_inferred__1_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__1_carry_i_8
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_ ),
        .I1(w_scr_h_m1[0]),
        .I2(\u_ras/u_ras_state/r_v1_y_reg_n_0_[1] ),
        .I3(w_scr_h_m1[1]),
        .O(result3_inferred__1_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    result3_inferred__2_carry__0_i_1
       (.I0(w_scr_h_m1[10]),
        .I1(\u_ras/u_ras_state/r_v0_y_reg_n_0_[10] ),
        .I2(w_scr_h_m1[11]),
        .O(result3_inferred__2_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__2_carry__0_i_2
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[8] ),
        .I1(w_scr_h_m1[8]),
        .I2(w_scr_h_m1[9]),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[9] ),
        .O(result3_inferred__2_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    result3_inferred__2_carry__0_i_3
       (.I0(w_scr_h_m1[14]),
        .I1(w_scr_h_m1[15]),
        .O(result3_inferred__2_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    result3_inferred__2_carry__0_i_4
       (.I0(w_scr_h_m1[12]),
        .I1(w_scr_h_m1[13]),
        .O(result3_inferred__2_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h09)) 
    result3_inferred__2_carry__0_i_5
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[10] ),
        .I1(w_scr_h_m1[10]),
        .I2(w_scr_h_m1[11]),
        .O(result3_inferred__2_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__2_carry__0_i_6
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[8] ),
        .I1(w_scr_h_m1[8]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[9] ),
        .I3(w_scr_h_m1[9]),
        .O(result3_inferred__2_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__2_carry_i_1
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[6] ),
        .I1(w_scr_h_m1[6]),
        .I2(w_scr_h_m1[7]),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[7] ),
        .O(result3_inferred__2_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__2_carry_i_2
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[4] ),
        .I1(w_scr_h_m1[4]),
        .I2(w_scr_h_m1[5]),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[5] ),
        .O(result3_inferred__2_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__2_carry_i_3
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[2] ),
        .I1(w_scr_h_m1[2]),
        .I2(w_scr_h_m1[3]),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[3] ),
        .O(result3_inferred__2_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__2_carry_i_4
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_ ),
        .I1(w_scr_h_m1[0]),
        .I2(w_scr_h_m1[1]),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[1] ),
        .O(result3_inferred__2_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__2_carry_i_5
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[6] ),
        .I1(w_scr_h_m1[6]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[7] ),
        .I3(w_scr_h_m1[7]),
        .O(result3_inferred__2_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__2_carry_i_6
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[4] ),
        .I1(w_scr_h_m1[4]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[5] ),
        .I3(w_scr_h_m1[5]),
        .O(result3_inferred__2_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__2_carry_i_7
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[2] ),
        .I1(w_scr_h_m1[2]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[3] ),
        .I3(w_scr_h_m1[3]),
        .O(result3_inferred__2_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__2_carry_i_8
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_ ),
        .I1(w_scr_h_m1[0]),
        .I2(\u_ras/u_ras_state/r_v0_y_reg_n_0_[1] ),
        .I3(w_scr_h_m1[1]),
        .O(result3_inferred__2_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    result3_inferred__3_carry__0_i_1
       (.I0(w_scr_w_m1[10]),
        .I1(\u_ras/u_ras_state/r_v2_x_reg_n_0_[10] ),
        .I2(w_scr_w_m1[11]),
        .O(result3_inferred__3_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__3_carry__0_i_2
       (.I0(\u_ras/u_ras_state/r_v2_x_reg_n_0_[8] ),
        .I1(w_scr_w_m1[8]),
        .I2(w_scr_w_m1[9]),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[9] ),
        .O(result3_inferred__3_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    result3_inferred__3_carry__0_i_3
       (.I0(w_scr_w_m1[14]),
        .I1(w_scr_w_m1[15]),
        .O(result3_inferred__3_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    result3_inferred__3_carry__0_i_4
       (.I0(w_scr_w_m1[12]),
        .I1(w_scr_w_m1[13]),
        .O(result3_inferred__3_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h09)) 
    result3_inferred__3_carry__0_i_5
       (.I0(\u_ras/u_ras_state/r_v2_x_reg_n_0_[10] ),
        .I1(w_scr_w_m1[10]),
        .I2(w_scr_w_m1[11]),
        .O(result3_inferred__3_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__3_carry__0_i_6
       (.I0(\u_ras/u_ras_state/r_v2_x_reg_n_0_[8] ),
        .I1(w_scr_w_m1[8]),
        .I2(\u_ras/u_ras_state/r_v2_x_reg_n_0_[9] ),
        .I3(w_scr_w_m1[9]),
        .O(result3_inferred__3_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__3_carry_i_1
       (.I0(\u_ras/u_ras_state/r_v2_x_reg_n_0_[6] ),
        .I1(w_scr_w_m1[6]),
        .I2(w_scr_w_m1[7]),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[7] ),
        .O(result3_inferred__3_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__3_carry_i_2
       (.I0(\u_ras/u_ras_state/r_v2_x_reg_n_0_[4] ),
        .I1(w_scr_w_m1[4]),
        .I2(w_scr_w_m1[5]),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[5] ),
        .O(result3_inferred__3_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__3_carry_i_3
       (.I0(\u_ras/u_ras_state/r_v2_x_reg_n_0_[2] ),
        .I1(w_scr_w_m1[2]),
        .I2(w_scr_w_m1[3]),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[3] ),
        .O(result3_inferred__3_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__3_carry_i_4
       (.I0(\u_ras/u_ras_state/r_v2_x_reg_n_0_ ),
        .I1(w_scr_w_m1[0]),
        .I2(w_scr_w_m1[1]),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[1] ),
        .O(result3_inferred__3_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__3_carry_i_5
       (.I0(\u_ras/u_ras_state/r_v2_x_reg_n_0_[6] ),
        .I1(w_scr_w_m1[6]),
        .I2(\u_ras/u_ras_state/r_v2_x_reg_n_0_[7] ),
        .I3(w_scr_w_m1[7]),
        .O(result3_inferred__3_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__3_carry_i_6
       (.I0(\u_ras/u_ras_state/r_v2_x_reg_n_0_[4] ),
        .I1(w_scr_w_m1[4]),
        .I2(\u_ras/u_ras_state/r_v2_x_reg_n_0_[5] ),
        .I3(w_scr_w_m1[5]),
        .O(result3_inferred__3_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__3_carry_i_7
       (.I0(\u_ras/u_ras_state/r_v2_x_reg_n_0_[2] ),
        .I1(w_scr_w_m1[2]),
        .I2(\u_ras/u_ras_state/r_v2_x_reg_n_0_[3] ),
        .I3(w_scr_w_m1[3]),
        .O(result3_inferred__3_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__3_carry_i_8
       (.I0(\u_ras/u_ras_state/r_v2_x_reg_n_0_ ),
        .I1(w_scr_w_m1[0]),
        .I2(\u_ras/u_ras_state/r_v2_x_reg_n_0_[1] ),
        .I3(w_scr_w_m1[1]),
        .O(result3_inferred__3_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    result3_inferred__4_carry__0_i_1
       (.I0(w_scr_h_m1[10]),
        .I1(\u_ras/u_ras_state/r_v2_y_reg_n_0_[10] ),
        .I2(w_scr_h_m1[11]),
        .O(result3_inferred__4_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__4_carry__0_i_2
       (.I0(\u_ras/u_ras_state/r_v2_y_reg_n_0_[8] ),
        .I1(w_scr_h_m1[8]),
        .I2(w_scr_h_m1[9]),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[9] ),
        .O(result3_inferred__4_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    result3_inferred__4_carry__0_i_3
       (.I0(w_scr_h_m1[14]),
        .I1(w_scr_h_m1[15]),
        .O(result3_inferred__4_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    result3_inferred__4_carry__0_i_4
       (.I0(w_scr_h_m1[12]),
        .I1(w_scr_h_m1[13]),
        .O(result3_inferred__4_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h09)) 
    result3_inferred__4_carry__0_i_5
       (.I0(\u_ras/u_ras_state/r_v2_y_reg_n_0_[10] ),
        .I1(w_scr_h_m1[10]),
        .I2(w_scr_h_m1[11]),
        .O(result3_inferred__4_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__4_carry__0_i_6
       (.I0(\u_ras/u_ras_state/r_v2_y_reg_n_0_[8] ),
        .I1(w_scr_h_m1[8]),
        .I2(\u_ras/u_ras_state/r_v2_y_reg_n_0_[9] ),
        .I3(w_scr_h_m1[9]),
        .O(result3_inferred__4_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__4_carry_i_1
       (.I0(\u_ras/u_ras_state/r_v2_y_reg_n_0_[6] ),
        .I1(w_scr_h_m1[6]),
        .I2(w_scr_h_m1[7]),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[7] ),
        .O(result3_inferred__4_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__4_carry_i_2
       (.I0(\u_ras/u_ras_state/r_v2_y_reg_n_0_[4] ),
        .I1(w_scr_h_m1[4]),
        .I2(w_scr_h_m1[5]),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[5] ),
        .O(result3_inferred__4_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__4_carry_i_3
       (.I0(\u_ras/u_ras_state/r_v2_y_reg_n_0_[2] ),
        .I1(w_scr_h_m1[2]),
        .I2(w_scr_h_m1[3]),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[3] ),
        .O(result3_inferred__4_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    result3_inferred__4_carry_i_4
       (.I0(\u_ras/u_ras_state/r_v2_y_reg_n_0_ ),
        .I1(w_scr_h_m1[0]),
        .I2(w_scr_h_m1[1]),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[1] ),
        .O(result3_inferred__4_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__4_carry_i_5
       (.I0(\u_ras/u_ras_state/r_v2_y_reg_n_0_[6] ),
        .I1(w_scr_h_m1[6]),
        .I2(\u_ras/u_ras_state/r_v2_y_reg_n_0_[7] ),
        .I3(w_scr_h_m1[7]),
        .O(result3_inferred__4_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__4_carry_i_6
       (.I0(\u_ras/u_ras_state/r_v2_y_reg_n_0_[4] ),
        .I1(w_scr_h_m1[4]),
        .I2(\u_ras/u_ras_state/r_v2_y_reg_n_0_[5] ),
        .I3(w_scr_h_m1[5]),
        .O(result3_inferred__4_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__4_carry_i_7
       (.I0(\u_ras/u_ras_state/r_v2_y_reg_n_0_[2] ),
        .I1(w_scr_h_m1[2]),
        .I2(\u_ras/u_ras_state/r_v2_y_reg_n_0_[3] ),
        .I3(w_scr_h_m1[3]),
        .O(result3_inferred__4_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    result3_inferred__4_carry_i_8
       (.I0(\u_ras/u_ras_state/r_v2_y_reg_n_0_ ),
        .I1(w_scr_h_m1[0]),
        .I2(\u_ras/u_ras_state/r_v2_y_reg_n_0_[1] ),
        .I3(w_scr_h_m1[1]),
        .O(result3_inferred__4_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    s_wb_ack_o_INST_0
       (.I0(s_wb_stb_i),
        .I1(s_wb_we_i),
        .I2(\u_sys/r_rstr ),
        .O(s_wb_ack_o));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[11]_i_2 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[11] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [11]),
        .O(\u_fadd/r_mats[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[11]_i_2__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[11] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [11]),
        .O(\u_fadd/r_mats ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[11]_i_3 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[10] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [10]),
        .O(\u_fadd/r_mats[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[11]_i_3__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[10] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [10]),
        .O(\u_fadd/r_mats[11]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[11]_i_4 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[9] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [9]),
        .O(\u_fadd/r_mats[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[11]_i_4__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[9] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [9]),
        .O(\u_fadd/r_mats[11]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[11]_i_5 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[8] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [8]),
        .O(\u_fadd/r_mats[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[11]_i_5__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[8] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [8]),
        .O(\u_fadd/r_mats[11]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[15]_i_2 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[15] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [15]),
        .O(\u_fadd/r_mats[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[15]_i_2__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[15] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [15]),
        .O(\u_fadd/r_mats[15]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[15]_i_3 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[14] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [14]),
        .O(\u_fadd/r_mats[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[15]_i_3__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[14] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [14]),
        .O(\u_fadd/r_mats[15]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[15]_i_4 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[13] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [13]),
        .O(\u_fadd/r_mats[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[15]_i_4__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[13] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [13]),
        .O(\u_fadd/r_mats[15]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[15]_i_5 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[12] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [12]),
        .O(\u_fadd/r_mats[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[15]_i_5__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[12] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [12]),
        .O(\u_fadd/r_mats[15]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[3]_i_2 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [3]),
        .O(\u_fadd/r_mats[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[3]_i_2__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [3]),
        .O(\u_fadd/r_mats[3]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[3]_i_3 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[2] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [2]),
        .O(\u_fadd/r_mats[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[3]_i_3__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[2] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [2]),
        .O(\u_fadd/r_mats[3]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[3]_i_4 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[1] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [1]),
        .O(\u_fadd/r_mats[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[3]_i_4__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[1] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [1]),
        .O(\u_fadd/r_mats[3]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[7]_i_2 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[7] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [7]),
        .O(\u_fadd/r_mats[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[7]_i_2__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[7] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [7]),
        .O(\u_fadd/r_mats[7]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[7]_i_3 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[6] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [6]),
        .O(\u_fadd/r_mats[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[7]_i_3__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[6] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [6]),
        .O(\u_fadd/r_mats[7]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[7]_i_4 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[5] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [5]),
        .O(\u_fadd/r_mats[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[7]_i_4__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[5] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [5]),
        .O(\u_fadd/r_mats[7]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[7]_i_5 
       (.I0(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[4] ),
        .I1(\u_geo/u_geo_clip/r_sub ),
        .I2(\u_geo/u_geo_clip/r_f0 [4]),
        .O(\u_fadd/r_mats[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd/r_mats[7]_i_5__0 
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[4] ),
        .I1(\u_geo/u_geo_viewport/r_sub ),
        .I2(\u_geo/u_geo_viewport/r_f0 [4]),
        .O(\u_fadd/r_mats[7]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[11]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [11]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [11]),
        .O(\u_fadd_m01/r_mats ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[11]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [10]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [10]),
        .O(\u_fadd_m01/r_mats[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[11]_i_4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [9]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [9]),
        .O(\u_fadd_m01/r_mats[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[11]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [8]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [8]),
        .O(\u_fadd_m01/r_mats[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[15]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [15]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [15]),
        .O(\u_fadd_m01/r_mats[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[15]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [14]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [14]),
        .O(\u_fadd_m01/r_mats[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[15]_i_4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [13]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [13]),
        .O(\u_fadd_m01/r_mats[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[15]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [12]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [12]),
        .O(\u_fadd_m01/r_mats[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[3]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [3]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [3]),
        .O(\u_fadd_m01/r_mats[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[3]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [2]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [2]),
        .O(\u_fadd_m01/r_mats[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[3]_i_4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [1]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [1]),
        .O(\u_fadd_m01/r_mats[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[7]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [7]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [7]),
        .O(\u_fadd_m01/r_mats[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[7]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [6]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [6]),
        .O(\u_fadd_m01/r_mats[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[7]_i_4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [5]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [5]),
        .O(\u_fadd_m01/r_mats[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m01/r_mats[7]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [4]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [4]),
        .O(\u_fadd_m01/r_mats[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[11]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [11]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [11]),
        .O(\u_fadd_m0123/r_mats ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[11]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [10]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [10]),
        .O(\u_fadd_m0123/r_mats[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[11]_i_4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [9]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [9]),
        .O(\u_fadd_m0123/r_mats[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[11]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [8]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [8]),
        .O(\u_fadd_m0123/r_mats[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[15]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [15]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [15]),
        .O(\u_fadd_m0123/r_mats[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[15]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [14]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [14]),
        .O(\u_fadd_m0123/r_mats[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[15]_i_4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [13]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [13]),
        .O(\u_fadd_m0123/r_mats[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[15]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [12]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [12]),
        .O(\u_fadd_m0123/r_mats[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[3]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [3]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [3]),
        .O(\u_fadd_m0123/r_mats[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[3]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [2]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [2]),
        .O(\u_fadd_m0123/r_mats[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[3]_i_4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [1]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [1]),
        .O(\u_fadd_m0123/r_mats[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[7]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [7]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [7]),
        .O(\u_fadd_m0123/r_mats[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[7]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [6]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [6]),
        .O(\u_fadd_m0123/r_mats[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[7]_i_4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [5]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [5]),
        .O(\u_fadd_m0123/r_mats[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m0123/r_mats[7]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [4]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [4]),
        .O(\u_fadd_m0123/r_mats[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[11]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [11]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [11]),
        .O(\u_fadd_m23/r_mats ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[11]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [10]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [10]),
        .O(\u_fadd_m23/r_mats[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[11]_i_4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [9]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [9]),
        .O(\u_fadd_m23/r_mats[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[11]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [8]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [8]),
        .O(\u_fadd_m23/r_mats[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[15]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [15]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [15]),
        .O(\u_fadd_m23/r_mats[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[15]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [14]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [14]),
        .O(\u_fadd_m23/r_mats[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[15]_i_4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [13]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [13]),
        .O(\u_fadd_m23/r_mats[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[15]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [12]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [12]),
        .O(\u_fadd_m23/r_mats[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[3]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [3]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [3]),
        .O(\u_fadd_m23/r_mats[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[3]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [2]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [2]),
        .O(\u_fadd_m23/r_mats[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[3]_i_4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [1]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [1]),
        .O(\u_fadd_m23/r_mats[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[7]_i_2 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [7]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [7]),
        .O(\u_fadd_m23/r_mats[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[7]_i_3 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [6]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [6]),
        .O(\u_fadd_m23/r_mats[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[7]_i_4 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [5]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [5]),
        .O(\u_fadd_m23/r_mats[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \u_fadd_m23/r_mats[7]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [4]),
        .I1(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .I2(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [4]),
        .O(\u_fadd_m23/r_mats[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0F0F0F0F0F1)) 
    \u_fmul/r_c[21]_i_1 
       (.I0(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [3]),
        .I1(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [4]),
        .I2(\r_c[20]_i_2__7_n_0 ),
        .I3(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [1]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [2]),
        .I5(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [0]),
        .O(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0F0F0F0F0F1)) 
    \u_fmul/r_c[21]_i_1__0 
       (.I0(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [3]),
        .I1(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [4]),
        .I2(\r_c[20]_i_2__9_n_0 ),
        .I3(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [1]),
        .I4(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [2]),
        .I5(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [0]),
        .O(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFB847)) 
    \u_fmul/r_ce_tmp_1z[0]_i_1 
       (.I0(\u_geo/w_vx_pdiv [16]),
        .I1(\r_ce_tmp_1z[4]_i_3__2_n_0 ),
        .I2(\u_geo/w_vy_pdiv [16]),
        .I3(\u_geo/u_geo_persdiv/w_b_exp [0]),
        .I4(\u_geo/u_geo_persdiv/u_fmul/w_adder_out ),
        .O(\u_fmul/r_ce_tmp_1z[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFE41B)) 
    \u_fmul/r_ce_tmp_1z[0]_i_1__0 
       (.I0(\r_ce_tmp_1z[4]_i_3__3_n_0 ),
        .I1(w_vh[16]),
        .I2(w_vw[16]),
        .I3(\u_geo/u_geo_viewport/w_a_exp [0]),
        .I4(\u_geo/u_geo_viewport/u_fmul/w_adder_out ),
        .O(\u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFB84747B8)) 
    \u_fmul/r_ce_tmp_1z[1]_i_1 
       (.I0(\u_geo/w_vx_pdiv [17]),
        .I1(\r_ce_tmp_1z[4]_i_3__2_n_0 ),
        .I2(\u_geo/w_vy_pdiv [17]),
        .I3(\u_geo/u_geo_persdiv/w_b_exp [1]),
        .I4(\r_ce_tmp_1z[1]_i_2__3_n_0 ),
        .I5(\u_geo/u_geo_persdiv/u_fmul/w_adder_out ),
        .O(\u_fmul/r_ce_tmp_1z[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF665A99A5)) 
    \u_fmul/r_ce_tmp_1z[1]_i_1__0 
       (.I0(\u_geo/u_geo_viewport/w_a_exp [1]),
        .I1(w_vw[17]),
        .I2(w_vh[17]),
        .I3(\r_ce_tmp_1z[4]_i_3__3_n_0 ),
        .I4(\r_ce_tmp_1z[1]_i_2__4_n_0 ),
        .I5(\u_geo/u_geo_viewport/u_fmul/w_adder_out ),
        .O(\u_fmul/r_ce_tmp_1z[1]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF66699969)) 
    \u_fmul/r_ce_tmp_1z[2]_i_1 
       (.I0(\r_ce_tmp_1z[2]_i_2__3_n_0 ),
        .I1(\u_geo/u_geo_persdiv/w_b_exp [2]),
        .I2(\u_geo/w_vy_pdiv [18]),
        .I3(\r_ce_tmp_1z[4]_i_3__2_n_0 ),
        .I4(\u_geo/w_vx_pdiv [18]),
        .I5(\u_geo/u_geo_persdiv/u_fmul/w_adder_out ),
        .O(\u_fmul/r_ce_tmp_1z[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF99966966)) 
    \u_fmul/r_ce_tmp_1z[2]_i_1__0 
       (.I0(\r_ce_tmp_1z[2]_i_2__4_n_0 ),
        .I1(\u_geo/u_geo_viewport/w_a_exp [2]),
        .I2(\r_ce_tmp_1z[4]_i_3__3_n_0 ),
        .I3(w_vh[18]),
        .I4(w_vw[18]),
        .I5(\u_geo/u_geo_viewport/u_fmul/w_adder_out ),
        .O(\u_fmul/r_ce_tmp_1z[2]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF656A9A95)) 
    \u_fmul/r_ce_tmp_1z[3]_i_1 
       (.I0(\r_ce_tmp_1z[3]_i_2__3_n_0 ),
        .I1(\u_geo/w_vx_pdiv [19]),
        .I2(\r_ce_tmp_1z[4]_i_3__2_n_0 ),
        .I3(\u_geo/w_vy_pdiv [19]),
        .I4(\u_geo/u_geo_persdiv/w_b_exp [3]),
        .I5(\u_geo/u_geo_persdiv/u_fmul/w_adder_out ),
        .O(\u_fmul/r_ce_tmp_1z[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFA965569A)) 
    \u_fmul/r_ce_tmp_1z[3]_i_1__0 
       (.I0(\r_ce_tmp_1z[3]_i_2__4_n_0 ),
        .I1(\r_ce_tmp_1z[4]_i_3__3_n_0 ),
        .I2(w_vh[19]),
        .I3(w_vw[19]),
        .I4(\u_geo/u_geo_viewport/w_a_exp [3]),
        .I5(\u_geo/u_geo_viewport/u_fmul/w_adder_out ),
        .O(\u_fmul/r_ce_tmp_1z[3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hE21DFFE2)) 
    \u_fmul/r_ce_tmp_1z[4]_i_2 
       (.I0(\u_geo/w_vy_pdiv [20]),
        .I1(\r_ce_tmp_1z[4]_i_3__2_n_0 ),
        .I2(\u_geo/w_vx_pdiv [20]),
        .I3(\u_geo/u_geo_persdiv/w_b_exp [4]),
        .I4(\r_ce_tmp_1z[4]_i_4__2_n_0 ),
        .O(\u_fmul/r_ce_tmp_1z[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99A5EEFA)) 
    \u_fmul/r_ce_tmp_1z[4]_i_2__0 
       (.I0(\u_geo/u_geo_viewport/w_a_exp [4]),
        .I1(w_vw[20]),
        .I2(w_vh[20]),
        .I3(\r_ce_tmp_1z[4]_i_3__3_n_0 ),
        .I4(\r_ce_tmp_1z[4]_i_4__3_n_0 ),
        .O(\u_fmul/r_ce_tmp_1z[4]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \u_frcp/ 
       (.I0(\u_geo/w_vw_clip [20]),
        .I1(\u_geo/w_vw_clip [19]),
        .I2(\u_geo/w_vw_clip [16]),
        .I3(\u_geo/w_vw_clip [18]),
        .I4(\u_geo/w_vw_clip [17]),
        .O(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \u_frcp/frcp_rom/r_c[30]_i_1 
       (.I0(g0_b30_n_0),
        .I1(\u_geo/w_vw_clip [14]),
        .O(\u_frcp/frcp_rom/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFFFFFF)) 
    \u_geo/r_int_i_4 
       (.I0(\u_geo/u_geo_cull/r_state [0]),
        .I1(\u_geo/u_geo_cull/r_state [1]),
        .I2(\u_geo/w_state_clip ),
        .I3(\u_geo/w_state_mat ),
        .I4(\u_geo/w_dma_end ),
        .O(\u_geo/r_int_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \u_geo/r_int_i_5 
       (.I0(\u_geo/u_geo_viewport/r_state [3]),
        .I1(\u_geo/u_geo_viewport/r_state [0]),
        .I2(\u_geo/u_geo_viewport/r_state [1]),
        .I3(\u_geo/u_geo_viewport/r_state [2]),
        .I4(\u_geo/w_state_if ),
        .I5(\u_geo/w_state_pd ),
        .O(\u_geo/r_int_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/FSM_onehot_r_state_reg[0] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[9]_i_1_n_0 ),
        .D(\u_geo/w_en_clip ),
        .Q(\u_geo/w_state_clip ),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/FSM_onehot_r_state_reg[1] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[9]_i_1_n_0 ),
        .D(\u_geo/w_state_clip ),
        .Q(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/FSM_onehot_r_state_reg[2] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[9]_i_1_n_0 ),
        .D(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_ ),
        .Q(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/FSM_onehot_r_state_reg[3] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[9]_i_1_n_0 ),
        .D(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[2] ),
        .Q(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/FSM_onehot_r_state_reg[4] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[9]_i_1_n_0 ),
        .D(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[3] ),
        .Q(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/FSM_onehot_r_state_reg[5] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[9]_i_1_n_0 ),
        .D(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[4] ),
        .Q(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/FSM_onehot_r_state_reg[6] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[9]_i_1_n_0 ),
        .D(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[5] ),
        .Q(\u_geo/u_geo_clip/r_bc ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/FSM_onehot_r_state_reg[7] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[9]_i_1_n_0 ),
        .D(\u_geo/u_geo_clip/r_bc ),
        .Q(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[7] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/FSM_onehot_r_state_reg[8] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[9]_i_1_n_0 ),
        .D(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[7] ),
        .Q(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[8] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/FSM_onehot_r_state_reg[9] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[9]_i_1_n_0 ),
        .D(\u_geo/u_geo_clip/FSM_onehot_r_state_reg_n_0_[8] ),
        .Q(\u_geo/w_en_clip ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_bc_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_bc),
        .Q(\u_geo/w_outcode_clip [0]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_bc_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_bc[1]_i_1_n_0 ),
        .Q(\u_geo/w_outcode_clip [1]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_bc_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_bc[2]_i_1_n_0 ),
        .Q(\u_geo/w_outcode_clip [2]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_bc_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_bc[3]_i_1_n_0 ),
        .Q(\u_geo/w_outcode_clip [3]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_bc_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_bc[4]_i_1_n_0 ),
        .Q(\u_geo/w_outcode_clip [4]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_bc_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_bc[5]_i_1_n_0 ),
        .Q(\u_geo/w_outcode_clip [5]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[0] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [0]),
        .Q(\u_geo/w_vw_clip [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[10] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [10]),
        .Q(\u_geo/w_vw_clip [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[11] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [11]),
        .Q(\u_geo/w_vw_clip [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[12] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [12]),
        .Q(\u_geo/w_vw_clip [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[13] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [13]),
        .Q(\u_geo/w_vw_clip [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[14] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [14]),
        .Q(\u_geo/w_vw_clip [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[15] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [15]),
        .Q(\u_geo/u_geo_clip/r_vw_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[16] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [16]),
        .Q(\u_geo/w_vw_clip [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[17] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [17]),
        .Q(\u_geo/w_vw_clip [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[18] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [18]),
        .Q(\u_geo/w_vw_clip [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[19] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [19]),
        .Q(\u_geo/w_vw_clip [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[1] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [1]),
        .Q(\u_geo/w_vw_clip [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[20] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [20]),
        .Q(\u_geo/w_vw_clip [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[21] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [21]),
        .Q(\u_geo/w_vw_clip [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[2] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [2]),
        .Q(\u_geo/w_vw_clip [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[3] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [3]),
        .Q(\u_geo/w_vw_clip [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[4] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [4]),
        .Q(\u_geo/w_vw_clip [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[5] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [5]),
        .Q(\u_geo/w_vw_clip [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[6] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [6]),
        .Q(\u_geo/w_vw_clip [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[7] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [7]),
        .Q(\u_geo/w_vw_clip [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[8] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [8]),
        .Q(\u_geo/w_vw_clip [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vw_reg[9] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vw_mvp [9]),
        .Q(\u_geo/w_vw_clip [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[0] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [0]),
        .Q(\u_geo/w_vx_clip [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[10] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [10]),
        .Q(\u_geo/w_vx_clip [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[11] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [11]),
        .Q(\u_geo/w_vx_clip [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[12] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [12]),
        .Q(\u_geo/w_vx_clip [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[13] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [13]),
        .Q(\u_geo/w_vx_clip [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[14] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [14]),
        .Q(\u_geo/w_vx_clip [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[15] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [15]),
        .Q(\u_geo/w_vx_clip [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[16] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [16]),
        .Q(\u_geo/w_vx_clip [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[17] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [17]),
        .Q(\u_geo/w_vx_clip [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[18] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [18]),
        .Q(\u_geo/w_vx_clip [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[19] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [19]),
        .Q(\u_geo/w_vx_clip [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[1] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [1]),
        .Q(\u_geo/w_vx_clip [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[20] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [20]),
        .Q(\u_geo/w_vx_clip [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[21] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [21]),
        .Q(\u_geo/w_vx_clip [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[2] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [2]),
        .Q(\u_geo/w_vx_clip [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[3] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [3]),
        .Q(\u_geo/w_vx_clip [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[4] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [4]),
        .Q(\u_geo/w_vx_clip [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[5] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [5]),
        .Q(\u_geo/w_vx_clip [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[6] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [6]),
        .Q(\u_geo/w_vx_clip [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[7] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [7]),
        .Q(\u_geo/w_vx_clip [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[8] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [8]),
        .Q(\u_geo/w_vx_clip [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vx_reg[9] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vx_mvp [9]),
        .Q(\u_geo/w_vx_clip [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[0] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [0]),
        .Q(\u_geo/w_vy_clip [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[10] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [10]),
        .Q(\u_geo/w_vy_clip [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[11] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [11]),
        .Q(\u_geo/w_vy_clip [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[12] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [12]),
        .Q(\u_geo/w_vy_clip [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[13] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [13]),
        .Q(\u_geo/w_vy_clip [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[14] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [14]),
        .Q(\u_geo/w_vy_clip [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[15] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [15]),
        .Q(\u_geo/w_vy_clip [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[16] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [16]),
        .Q(\u_geo/w_vy_clip [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[17] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [17]),
        .Q(\u_geo/w_vy_clip [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[18] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [18]),
        .Q(\u_geo/w_vy_clip [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[19] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [19]),
        .Q(\u_geo/w_vy_clip [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[1] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [1]),
        .Q(\u_geo/w_vy_clip [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[20] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [20]),
        .Q(\u_geo/w_vy_clip [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[21] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [21]),
        .Q(\u_geo/w_vy_clip [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[2] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [2]),
        .Q(\u_geo/w_vy_clip [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[3] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [3]),
        .Q(\u_geo/w_vy_clip [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[4] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [4]),
        .Q(\u_geo/w_vy_clip [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[5] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [5]),
        .Q(\u_geo/w_vy_clip [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[6] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [6]),
        .Q(\u_geo/w_vy_clip [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[7] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [7]),
        .Q(\u_geo/w_vy_clip [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[8] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [8]),
        .Q(\u_geo/w_vy_clip [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vy_reg[9] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vy_mvp [9]),
        .Q(\u_geo/w_vy_clip [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[0] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [0]),
        .Q(\u_geo/u_geo_clip/r_vz [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[10] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [10]),
        .Q(\u_geo/u_geo_clip/r_vz [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[11] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [11]),
        .Q(\u_geo/u_geo_clip/r_vz [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[12] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [12]),
        .Q(\u_geo/u_geo_clip/r_vz [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[13] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [13]),
        .Q(\u_geo/u_geo_clip/r_vz [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[14] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [14]),
        .Q(\u_geo/u_geo_clip/r_vz [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[15] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [15]),
        .Q(\u_geo/u_geo_clip/r_vz [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[16] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [16]),
        .Q(\u_geo/u_geo_clip/r_vz [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[17] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [17]),
        .Q(\u_geo/u_geo_clip/r_vz [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[18] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [18]),
        .Q(\u_geo/u_geo_clip/r_vz [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[19] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [19]),
        .Q(\u_geo/u_geo_clip/r_vz [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[1] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [1]),
        .Q(\u_geo/u_geo_clip/r_vz [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[20] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [20]),
        .Q(\u_geo/u_geo_clip/r_vz [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[21] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [21]),
        .Q(\u_geo/u_geo_clip/r_vz [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[2] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [2]),
        .Q(\u_geo/u_geo_clip/r_vz [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[3] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [3]),
        .Q(\u_geo/u_geo_clip/r_vz [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[4] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [4]),
        .Q(\u_geo/u_geo_clip/r_vz [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[5] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [5]),
        .Q(\u_geo/u_geo_clip/r_vz [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[6] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [6]),
        .Q(\u_geo/u_geo_clip/r_vz [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[7] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [7]),
        .Q(\u_geo/u_geo_clip/r_vz [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[8] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [8]),
        .Q(\u_geo/u_geo_clip/r_vz [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/r_vz_reg[9] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1_n_0 ),
        .D(\u_geo/w_vz_mvp [9]),
        .Q(\u_geo/u_geo_clip/r_vz [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry_n_0 ,\u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry_n_1 ,\u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry_n_2 ,\u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry_n_3 }),
        .CYINIT(\u_geo/u_geo_clip/r_exp_2z [0]),
        .DI({\u_geo/u_geo_clip/r_exp_2z [3:1],_inferred__1_carry_i_1__14_n_0}),
        .O(\u_geo/u_geo_clip/u_fadd/norm/f_incdec_return [3:0]),
        .S({_inferred__1_carry_i_2__6_n_0,_inferred__1_carry_i_3__6_n_0,_inferred__1_carry_i_4__6_n_0,_inferred__1_carry_i_5__7_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry__0 
       (.CI(\u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_clip/u_fadd/r_mats [16]}),
        .O({\u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry__0_n_4 ,\u_geo/u_geo_clip/u_fadd/norm/_inferred__1_carry__0_n_5 ,\u_geo/u_geo_clip/u_fadd/norm/f_incdec_return [5:4]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,_inferred__1_carry_i_1__13_n_0,_inferred__1_carry_i_2__18_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/u_fadd/w_c ),
        .Q(\u_geo/u_geo_clip/p_0_in0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_exp_1z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/u_fadd/w_exp_l [0]),
        .Q(\u_geo/u_geo_clip/r_exp_1z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_exp_1z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/u_fadd/w_exp_l [1]),
        .Q(\u_geo/u_geo_clip/r_exp_1z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_exp_1z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/u_fadd/w_exp_l [2]),
        .Q(\u_geo/u_geo_clip/r_exp_1z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_exp_1z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/u_fadd/w_exp_l [3]),
        .Q(\u_geo/u_geo_clip/r_exp_1z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_exp_1z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/u_fadd/w_exp_l [4]),
        .Q(\u_geo/u_geo_clip/r_exp_1z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_exp_2z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/r_exp_1z [0]),
        .Q(\u_geo/u_geo_clip/r_exp_2z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_exp_2z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/r_exp_1z [1]),
        .Q(\u_geo/u_geo_clip/r_exp_2z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_exp_2z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/r_exp_1z [2]),
        .Q(\u_geo/u_geo_clip/r_exp_2z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_exp_2z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/r_exp_1z [3]),
        .Q(\u_geo/u_geo_clip/r_exp_2z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_exp_2z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/r_exp_1z [4]),
        .Q(\u_geo/u_geo_clip/r_exp_2z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [0]),
        .Q(\u_geo/u_geo_clip/r_f0 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [10]),
        .Q(\u_geo/u_geo_clip/r_f0 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [11]),
        .Q(\u_geo/u_geo_clip/r_f0 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [12]),
        .Q(\u_geo/u_geo_clip/r_f0 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [13]),
        .Q(\u_geo/u_geo_clip/r_f0 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [14]),
        .Q(\u_geo/u_geo_clip/r_f0 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [15]),
        .Q(\u_geo/u_geo_clip/r_f0 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [1]),
        .Q(\u_geo/u_geo_clip/r_f0 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [2]),
        .Q(\u_geo/u_geo_clip/r_f0 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [3]),
        .Q(\u_geo/u_geo_clip/r_f0 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [4]),
        .Q(\u_geo/u_geo_clip/r_f0 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [5]),
        .Q(\u_geo/u_geo_clip/r_f0 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [6]),
        .Q(\u_geo/u_geo_clip/r_f0 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [7]),
        .Q(\u_geo/u_geo_clip/r_f0 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [8]),
        .Q(\u_geo/u_geo_clip/r_f0 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f0_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f0 [9]),
        .Q(\u_geo/u_geo_clip/r_f0 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [0]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [10]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [11]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [12]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [13]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [14]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [15]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [1]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [2]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [3]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [4]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [5]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [6]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [7]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [8]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_f1t_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_f1t [9]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_f1t_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [0]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [10]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [11]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [12]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [13]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [14]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [15]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [16]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [1]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [2]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [3]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [4]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [5]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [6]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [7]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [8]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_mats_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/w_mats [9]),
        .Q(\u_geo/u_geo_clip/u_fadd/r_mats [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_sign_1z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/u_fadd/w_sign ),
        .Q(\u_geo/u_geo_clip/r_sign_1z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_sign_2z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_clip/r_sign_1z ),
        .Q(\u_geo/u_geo_clip/u_fadd/r_sign_2z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_clip/u_fadd/r_sub_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_sub_i_1__3_n_0),
        .Q(\u_geo/u_geo_clip/r_sub ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_clip/u_fadd/w_mag_frac_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_clip/u_fadd/w_mag_frac_carry_n_0 ,\u_geo/u_geo_clip/u_fadd/w_mag_frac_carry_n_1 ,\u_geo/u_geo_clip/u_fadd/w_mag_frac_carry_n_2 ,\u_geo/u_geo_clip/u_fadd/w_mag_frac_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({w_mag_frac_carry_i_1__5_n_0,w_mag_frac_carry_i_2__5_n_0,w_mag_frac_carry_i_3__5_n_0,w_mag_frac_carry_i_4__5_n_0}),
        .S({w_mag_frac_carry_i_5__5_n_0,w_mag_frac_carry_i_6__5_n_0,w_mag_frac_carry_i_7__5_n_0,w_mag_frac_carry_i_8__5_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_clip/u_fadd/w_mag_frac_carry__0 
       (.CI(\u_geo/u_geo_clip/u_fadd/w_mag_frac_carry_n_0 ),
        .CO({\u_geo/u_geo_clip/data0 ,\u_geo/u_geo_clip/u_fadd/w_mag_frac_carry__0_n_1 ,\u_geo/u_geo_clip/u_fadd/w_mag_frac_carry__0_n_2 ,\u_geo/u_geo_clip/u_fadd/w_mag_frac_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({w_mag_frac_carry_i_1__6_n_0,w_mag_frac_carry_i_2__6_n_0,w_mag_frac_carry_i_3__6_n_0,w_mag_frac_carry_i_4__6_n_0}),
        .S({w_mag_frac_carry_i_5__6_n_0,w_mag_frac_carry_i_6__6_n_0,w_mag_frac_carry_i_7__6_n_0,w_mag_frac_carry_i_8__6_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(0),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \u_geo/u_geo_cull/f_multi_return 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,f_multi_return_i_13_n_0,f_multi_return_i_14_n_0,f_multi_return_i_15_n_0,f_multi_return_i_16_n_0,f_multi_return_i_17_n_0,f_multi_return_i_18_n_0,f_multi_return_i_19_n_0,f_multi_return_i_20_n_0,f_multi_return_i_21_n_0,f_multi_return_i_22_n_0,f_multi_return_i_23_n_0,f_multi_return_i_24_n_0}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,f_multi_return_i_1_n_0,f_multi_return_i_2_n_0,f_multi_return_i_3_n_0,f_multi_return_i_4_n_0,f_multi_return_i_5_n_0,f_multi_return_i_6_n_0,f_multi_return_i_7_n_0,f_multi_return_i_8_n_0,f_multi_return_i_9_n_0,f_multi_return_i_10_n_0,f_multi_return_i_11_n_0,f_multi_return_i_12_n_0}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_cull/f_multi_return0_n_82 ,\u_geo/u_geo_cull/f_multi_return0_n_83 ,\u_geo/u_geo_cull/f_multi_return0_n_84 ,\u_geo/u_geo_cull/f_multi_return0_n_85 ,\u_geo/u_geo_cull/f_multi_return0_n_86 ,\u_geo/u_geo_cull/f_multi_return0_n_87 ,\u_geo/u_geo_cull/f_multi_return0_n_88 ,\u_geo/u_geo_cull/f_multi_return0_n_89 ,\u_geo/u_geo_cull/f_multi_return0_n_90 ,\u_geo/u_geo_cull/f_multi_return0_n_91 ,\u_geo/u_geo_cull/f_multi_return0_n_92 ,\u_geo/u_geo_cull/f_multi_return0_n_93 ,\u_geo/u_geo_cull/f_multi_return0_n_94 ,\u_geo/u_geo_cull/f_multi_return0_n_95 ,\u_geo/u_geo_cull/f_multi_return0_n_96 ,\u_geo/u_geo_cull/f_multi_return0_n_97 ,\u_geo/u_geo_cull/f_multi_return0_n_98 ,\u_geo/u_geo_cull/f_multi_return0_n_99 ,\u_geo/u_geo_cull/f_multi_return0_n_100 ,\u_geo/u_geo_cull/f_multi_return0_n_101 ,\u_geo/u_geo_cull/f_multi_return0_n_102 ,\u_geo/u_geo_cull/f_multi_return0_n_103 ,\u_geo/u_geo_cull/f_multi_return0_n_104 ,\u_geo/u_geo_cull/f_multi_return0_n_105 }),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const1>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\u_geo/u_geo_cull/f_multi_return_n_58 ,\u_geo/u_geo_cull/f_multi_return_n_59 ,\u_geo/u_geo_cull/f_multi_return_n_60 ,\u_geo/u_geo_cull/f_multi_return_n_61 ,\u_geo/u_geo_cull/f_multi_return_n_62 ,\u_geo/u_geo_cull/f_multi_return_n_63 ,\u_geo/u_geo_cull/f_multi_return_n_64 ,\u_geo/u_geo_cull/f_multi_return_n_65 ,\u_geo/u_geo_cull/f_multi_return_n_66 ,\u_geo/u_geo_cull/f_multi_return_n_67 ,\u_geo/u_geo_cull/f_multi_return_n_68 ,\u_geo/u_geo_cull/f_multi_return_n_69 ,\u_geo/u_geo_cull/f_multi_return_n_70 ,\u_geo/u_geo_cull/f_multi_return_n_71 ,\u_geo/u_geo_cull/f_multi_return_n_72 ,\u_geo/u_geo_cull/f_multi_return_n_73 ,\u_geo/u_geo_cull/f_multi_return_n_74 ,\u_geo/u_geo_cull/f_multi_return_n_75 ,\u_geo/u_geo_cull/f_multi_return_n_76 ,\u_geo/u_geo_cull/f_multi_return_n_77 ,\u_geo/u_geo_cull/f_multi_return_n_78 ,\u_geo/u_geo_cull/f_multi_return_n_79 ,\u_geo/u_geo_cull/f_multi_return_n_80 ,\u_geo/u_geo_cull/f_multi_return_n_81 ,\u_geo/u_geo_cull/f_multi_return_n_82 ,\u_geo/u_geo_cull/f_multi_return_n_83 ,\u_geo/u_geo_cull/f_multi_return_n_84 ,\u_geo/u_geo_cull/f_multi_return_n_85 ,\u_geo/u_geo_cull/f_multi_return_n_86 ,\u_geo/u_geo_cull/f_multi_return_n_87 ,\u_geo/u_geo_cull/f_multi_return_n_88 ,\u_geo/u_geo_cull/f_multi_return_n_89 ,\u_geo/u_geo_cull/f_multi_return_n_90 ,\u_geo/u_geo_cull/f_multi_return_n_91 ,\u_geo/u_geo_cull/f_multi_return_n_92 ,\u_geo/u_geo_cull/f_multi_return_n_93 ,\u_geo/u_geo_cull/f_multi_return_n_94 ,\u_geo/u_geo_cull/f_multi_return_n_95 ,\u_geo/u_geo_cull/f_multi_return_n_96 ,\u_geo/u_geo_cull/f_multi_return_n_97 ,\u_geo/u_geo_cull/f_multi_return_n_98 ,\u_geo/u_geo_cull/f_multi_return_n_99 ,\u_geo/u_geo_cull/f_multi_return_n_100 ,\u_geo/u_geo_cull/f_multi_return_n_101 ,\u_geo/u_geo_cull/f_multi_return_n_102 ,\u_geo/u_geo_cull/f_multi_return_n_103 ,\u_geo/u_geo_cull/f_multi_return_n_104 ,\u_geo/u_geo_cull/f_multi_return_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \u_geo/u_geo_cull/f_multi_return0 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_cull/A }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_cull/B }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\u_geo/u_geo_cull/f_multi_return0_n_58 ,\u_geo/u_geo_cull/f_multi_return0_n_59 ,\u_geo/u_geo_cull/f_multi_return0_n_60 ,\u_geo/u_geo_cull/f_multi_return0_n_61 ,\u_geo/u_geo_cull/f_multi_return0_n_62 ,\u_geo/u_geo_cull/f_multi_return0_n_63 ,\u_geo/u_geo_cull/f_multi_return0_n_64 ,\u_geo/u_geo_cull/f_multi_return0_n_65 ,\u_geo/u_geo_cull/f_multi_return0_n_66 ,\u_geo/u_geo_cull/f_multi_return0_n_67 ,\u_geo/u_geo_cull/f_multi_return0_n_68 ,\u_geo/u_geo_cull/f_multi_return0_n_69 ,\u_geo/u_geo_cull/f_multi_return0_n_70 ,\u_geo/u_geo_cull/f_multi_return0_n_71 ,\u_geo/u_geo_cull/f_multi_return0_n_72 ,\u_geo/u_geo_cull/f_multi_return0_n_73 ,\u_geo/u_geo_cull/f_multi_return0_n_74 ,\u_geo/u_geo_cull/f_multi_return0_n_75 ,\u_geo/u_geo_cull/f_multi_return0_n_76 ,\u_geo/u_geo_cull/f_multi_return0_n_77 ,\u_geo/u_geo_cull/f_multi_return0_n_78 ,\u_geo/u_geo_cull/f_multi_return0_n_79 ,\u_geo/u_geo_cull/f_multi_return0_n_80 ,\u_geo/u_geo_cull/f_multi_return0_n_81 ,\u_geo/u_geo_cull/f_multi_return0_n_82 ,\u_geo/u_geo_cull/f_multi_return0_n_83 ,\u_geo/u_geo_cull/f_multi_return0_n_84 ,\u_geo/u_geo_cull/f_multi_return0_n_85 ,\u_geo/u_geo_cull/f_multi_return0_n_86 ,\u_geo/u_geo_cull/f_multi_return0_n_87 ,\u_geo/u_geo_cull/f_multi_return0_n_88 ,\u_geo/u_geo_cull/f_multi_return0_n_89 ,\u_geo/u_geo_cull/f_multi_return0_n_90 ,\u_geo/u_geo_cull/f_multi_return0_n_91 ,\u_geo/u_geo_cull/f_multi_return0_n_92 ,\u_geo/u_geo_cull/f_multi_return0_n_93 ,\u_geo/u_geo_cull/f_multi_return0_n_94 ,\u_geo/u_geo_cull/f_multi_return0_n_95 ,\u_geo/u_geo_cull/f_multi_return0_n_96 ,\u_geo/u_geo_cull/f_multi_return0_n_97 ,\u_geo/u_geo_cull/f_multi_return0_n_98 ,\u_geo/u_geo_cull/f_multi_return0_n_99 ,\u_geo/u_geo_cull/f_multi_return0_n_100 ,\u_geo/u_geo_cull/f_multi_return0_n_101 ,\u_geo/u_geo_cull/f_multi_return0_n_102 ,\u_geo/u_geo_cull/f_multi_return0_n_103 ,\u_geo/u_geo_cull/f_multi_return0_n_104 ,\u_geo/u_geo_cull/f_multi_return0_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_x_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_x_tri [0]),
        .Q(w_v0_x[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_x_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_x_tri [10]),
        .Q(w_v0_x[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_x_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_x_tri [11]),
        .Q(w_v0_x[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_x_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_x_tri [1]),
        .Q(w_v0_x[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_x_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_x_tri [2]),
        .Q(w_v0_x[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_x_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_x_tri [3]),
        .Q(w_v0_x[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_x_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_x_tri [4]),
        .Q(w_v0_x[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_x_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_x_tri [5]),
        .Q(w_v0_x[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_x_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_x_tri [6]),
        .Q(w_v0_x[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_x_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_x_tri [7]),
        .Q(w_v0_x[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_x_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_x_tri [8]),
        .Q(w_v0_x[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_x_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_x_tri [9]),
        .Q(w_v0_x[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_y_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_y_tri [0]),
        .Q(w_v0_y[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_y_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_y_tri [10]),
        .Q(w_v0_y[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_y_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_y_tri [11]),
        .Q(w_v0_y[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_y_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_y_tri [1]),
        .Q(w_v0_y[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_y_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_y_tri [2]),
        .Q(w_v0_y[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_y_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_y_tri [3]),
        .Q(w_v0_y[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_y_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_y_tri [4]),
        .Q(w_v0_y[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_y_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_y_tri [5]),
        .Q(w_v0_y[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_y_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_y_tri [6]),
        .Q(w_v0_y[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_y_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_y_tri [7]),
        .Q(w_v0_y[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_y_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_y_tri [8]),
        .Q(w_v0_y[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v0_y_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v0_y_tri [9]),
        .Q(w_v0_y[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_x_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_x_tri [0]),
        .Q(w_v1_x[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_x_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_x_tri [10]),
        .Q(w_v1_x[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_x_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_x_tri [11]),
        .Q(w_v1_x[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_x_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_x_tri [1]),
        .Q(w_v1_x[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_x_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_x_tri [2]),
        .Q(w_v1_x[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_x_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_x_tri [3]),
        .Q(w_v1_x[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_x_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_x_tri [4]),
        .Q(w_v1_x[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_x_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_x_tri [5]),
        .Q(w_v1_x[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_x_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_x_tri [6]),
        .Q(w_v1_x[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_x_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_x_tri [7]),
        .Q(w_v1_x[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_x_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_x_tri [8]),
        .Q(w_v1_x[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_x_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_x_tri [9]),
        .Q(w_v1_x[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_y_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_y_tri [0]),
        .Q(w_v1_y[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_y_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_y_tri [10]),
        .Q(w_v1_y[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_y_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_y_tri [11]),
        .Q(w_v1_y[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_y_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_y_tri [1]),
        .Q(w_v1_y[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_y_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_y_tri [2]),
        .Q(w_v1_y[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_y_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_y_tri [3]),
        .Q(w_v1_y[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_y_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_y_tri [4]),
        .Q(w_v1_y[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_y_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_y_tri [5]),
        .Q(w_v1_y[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_y_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_y_tri [6]),
        .Q(w_v1_y[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_y_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_y_tri [7]),
        .Q(w_v1_y[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_y_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_y_tri [8]),
        .Q(w_v1_y[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v1_y_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v1_y_tri [9]),
        .Q(w_v1_y[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_x_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_x_tri [0]),
        .Q(w_v2_x[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_x_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_x_tri [10]),
        .Q(w_v2_x[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_x_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_x_tri [11]),
        .Q(w_v2_x[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_x_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_x_tri [1]),
        .Q(w_v2_x[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_x_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_x_tri [2]),
        .Q(w_v2_x[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_x_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_x_tri [3]),
        .Q(w_v2_x[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_x_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_x_tri [4]),
        .Q(w_v2_x[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_x_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_x_tri [5]),
        .Q(w_v2_x[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_x_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_x_tri [6]),
        .Q(w_v2_x[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_x_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_x_tri [7]),
        .Q(w_v2_x[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_x_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_x_tri [8]),
        .Q(w_v2_x[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_x_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_x_tri [9]),
        .Q(w_v2_x[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_y_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_y_tri [0]),
        .Q(w_v2_y[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_y_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_y_tri [10]),
        .Q(w_v2_y[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_y_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_y_tri [11]),
        .Q(w_v2_y[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_y_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_y_tri [1]),
        .Q(w_v2_y[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_y_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_y_tri [2]),
        .Q(w_v2_y[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_y_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_y_tri [3]),
        .Q(w_v2_y[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_y_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_y_tri [4]),
        .Q(w_v2_y[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_y_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_y_tri [5]),
        .Q(w_v2_y[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_y_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_y_tri [6]),
        .Q(w_v2_y[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_y_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_y_tri [7]),
        .Q(w_v2_y[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_y_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_y_tri [8]),
        .Q(w_v2_y[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/o_v2_y_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_cull/w_set_tri ),
        .D(\u_geo/w_v2_y_tri [9]),
        .Q(w_v2_y[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_state_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_state),
        .Q(\u_geo/u_geo_cull/r_state [0]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_state_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_state[1]_i_1_n_0 ),
        .Q(\u_geo/u_geo_cull/r_state [1]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[0] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [0]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_ ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[10] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [10]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[10] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[11] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [11]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[11] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[12] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [12]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[12] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[13] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [13]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[13] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[14] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [14]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[14] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[15] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [15]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[15] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[16] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [16]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[16] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[17] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [17]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[17] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[18] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [18]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[18] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[19] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [19]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[19] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[1] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [1]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[1] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[20] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [20]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[20] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[21] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [21]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[21] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[22] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [22]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[22] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[23] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [23]),
        .Q(\u_geo/u_geo_cull/p_0_in ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[2] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [2]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[2] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[3] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [3]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[3] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[4] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [4]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[4] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[5] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [5]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[5] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[6] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [6]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[6] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[7] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [7]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[7] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[8] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [8]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[8] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_cull/r_sum_reg[9] 
       (.C(clk_i),
        .CE(\r_sum[23]_i_1_n_0 ),
        .D(\u_geo/u_geo_cull/p_1_in [9]),
        .Q(\u_geo/u_geo_cull/r_sum_reg_n_0_[9] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/FSM_onehot_r_state_reg[0] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[5]_i_1__0_n_0 ),
        .D(\u_geo/w_en_mvp ),
        .Q(\u_geo/w_state_mat ),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/FSM_onehot_r_state_reg[1] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[5]_i_1__0_n_0 ),
        .D(\u_geo/w_state_mat ),
        .Q(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/FSM_onehot_r_state_reg[2] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[5]_i_1__0_n_0 ),
        .D(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .Q(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/FSM_onehot_r_state_reg[3] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[5]_i_1__0_n_0 ),
        .D(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .Q(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/FSM_onehot_r_state_reg[4] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[5]_i_1__0_n_0 ),
        .D(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .Q(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[4] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/FSM_onehot_r_state_reg[5] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[5]_i_1__0_n_0 ),
        .D(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[4] ),
        .Q(\u_geo/w_en_mvp ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_lat_cnt_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_lat_cnt ),
        .D(r_vz_in),
        .Q(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_ ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_lat_cnt_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_lat_cnt ),
        .D(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_ ),
        .Q(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[1] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_lat_cnt_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_lat_cnt ),
        .D(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[1] ),
        .Q(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[2] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_lat_cnt_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_lat_cnt ),
        .D(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[2] ),
        .Q(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[3] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_lat_cnt_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_lat_cnt ),
        .D(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[3] ),
        .Q(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[4] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_lat_cnt_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_lat_cnt ),
        .D(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[4] ),
        .Q(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[5] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_lat_cnt_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_lat_cnt ),
        .D(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[5] ),
        .Q(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[6] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_lat_cnt_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_lat_cnt ),
        .D(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[6] ),
        .Q(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[7] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_lat_cnt_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_lat_cnt ),
        .D(\u_geo/u_geo_matrix/r_lat_cnt_reg_n_0_[7] ),
        .Q(\u_geo/u_geo_matrix/w_wait_end ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [0]),
        .Q(\u_geo/w_vw_mvp [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [10]),
        .Q(\u_geo/w_vw_mvp [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [11]),
        .Q(\u_geo/w_vw_mvp [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[12] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [12]),
        .Q(\u_geo/w_vw_mvp [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[13] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [13]),
        .Q(\u_geo/w_vw_mvp [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[14] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [14]),
        .Q(\u_geo/w_vw_mvp [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[15] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [15]),
        .Q(\u_geo/w_vw_mvp [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[16] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [16]),
        .Q(\u_geo/w_vw_mvp [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[17] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [17]),
        .Q(\u_geo/w_vw_mvp [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[18] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [18]),
        .Q(\u_geo/w_vw_mvp [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[19] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [19]),
        .Q(\u_geo/w_vw_mvp [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [1]),
        .Q(\u_geo/w_vw_mvp [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[20] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [20]),
        .Q(\u_geo/w_vw_mvp [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[21] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [21]),
        .Q(\u_geo/w_vw_mvp [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [2]),
        .Q(\u_geo/w_vw_mvp [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [3]),
        .Q(\u_geo/w_vw_mvp [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [4]),
        .Q(\u_geo/w_vw_mvp [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [5]),
        .Q(\u_geo/w_vw_mvp [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [6]),
        .Q(\u_geo/w_vw_mvp [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [7]),
        .Q(\u_geo/w_vw_mvp [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [8]),
        .Q(\u_geo/w_vw_mvp [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vw_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [9]),
        .Q(\u_geo/w_vw_mvp [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[0] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [0]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[10] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [10]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[11] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [11]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[12] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [12]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[13] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [13]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[14] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [14]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[15] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [15]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[16] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [16]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[17] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [17]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[18] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [18]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[19] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [19]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[1] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [1]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[20] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [20]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[21] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [21]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[2] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [2]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[3] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [3]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[4] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [4]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[5] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [5]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[6] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [6]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[7] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [7]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[8] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [8]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_in_reg[9] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vx_dma [9]),
        .Q(\u_geo/u_geo_matrix/r_vx_in [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [0]),
        .Q(\u_geo/w_vx_mvp [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [10]),
        .Q(\u_geo/w_vx_mvp [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [11]),
        .Q(\u_geo/w_vx_mvp [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[12] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [12]),
        .Q(\u_geo/w_vx_mvp [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[13] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [13]),
        .Q(\u_geo/w_vx_mvp [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[14] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [14]),
        .Q(\u_geo/w_vx_mvp [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[15] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [15]),
        .Q(\u_geo/w_vx_mvp [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[16] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [16]),
        .Q(\u_geo/w_vx_mvp [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[17] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [17]),
        .Q(\u_geo/w_vx_mvp [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[18] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [18]),
        .Q(\u_geo/w_vx_mvp [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[19] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [19]),
        .Q(\u_geo/w_vx_mvp [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [1]),
        .Q(\u_geo/w_vx_mvp [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[20] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [20]),
        .Q(\u_geo/w_vx_mvp [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[21] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [21]),
        .Q(\u_geo/w_vx_mvp [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [2]),
        .Q(\u_geo/w_vx_mvp [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [3]),
        .Q(\u_geo/w_vx_mvp [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [4]),
        .Q(\u_geo/w_vx_mvp [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [5]),
        .Q(\u_geo/w_vx_mvp [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [6]),
        .Q(\u_geo/w_vx_mvp [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [7]),
        .Q(\u_geo/w_vx_mvp [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [8]),
        .Q(\u_geo/w_vx_mvp [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vx_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/w_wait_end ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [9]),
        .Q(\u_geo/w_vx_mvp [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[0] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [0]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[10] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [10]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[11] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [11]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[12] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [12]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[13] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [13]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[14] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [14]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[15] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [15]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[16] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [16]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[17] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [17]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[18] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [18]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[19] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [19]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[1] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [1]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[20] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [20]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[21] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [21]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[2] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [2]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[3] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [3]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[4] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [4]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[5] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [5]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[6] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [6]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[7] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [7]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[8] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [8]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_in_reg[9] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vy_dma [9]),
        .Q(\u_geo/u_geo_matrix/r_vy_in [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [0]),
        .Q(\u_geo/w_vy_mvp [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [10]),
        .Q(\u_geo/w_vy_mvp [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [11]),
        .Q(\u_geo/w_vy_mvp [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[12] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [12]),
        .Q(\u_geo/w_vy_mvp [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[13] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [13]),
        .Q(\u_geo/w_vy_mvp [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[14] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [14]),
        .Q(\u_geo/w_vy_mvp [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[15] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [15]),
        .Q(\u_geo/w_vy_mvp [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[16] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [16]),
        .Q(\u_geo/w_vy_mvp [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[17] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [17]),
        .Q(\u_geo/w_vy_mvp [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[18] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [18]),
        .Q(\u_geo/w_vy_mvp [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[19] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [19]),
        .Q(\u_geo/w_vy_mvp [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [1]),
        .Q(\u_geo/w_vy_mvp [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[20] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [20]),
        .Q(\u_geo/w_vy_mvp [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[21] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [21]),
        .Q(\u_geo/w_vy_mvp [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [2]),
        .Q(\u_geo/w_vy_mvp [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [3]),
        .Q(\u_geo/w_vy_mvp [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [4]),
        .Q(\u_geo/w_vy_mvp [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [5]),
        .Q(\u_geo/w_vy_mvp [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [6]),
        .Q(\u_geo/w_vy_mvp [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [7]),
        .Q(\u_geo/w_vy_mvp [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [8]),
        .Q(\u_geo/w_vy_mvp [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vy_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [9]),
        .Q(\u_geo/w_vy_mvp [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[0] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [0]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[10] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [10]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[11] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [11]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[12] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [12]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[13] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [13]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[14] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [14]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[15] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [15]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[16] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [16]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[17] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [17]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[18] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [18]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[19] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [19]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[1] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [1]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[20] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [20]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[21] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [21]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[2] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [2]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[3] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [3]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[4] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [4]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[5] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [5]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[6] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [6]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[7] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [7]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[8] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [8]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_in_reg[9] 
       (.C(clk_i),
        .CE(r_vz_in),
        .D(\u_geo/w_vz_dma [9]),
        .Q(\u_geo/u_geo_matrix/r_vz_in [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [0]),
        .Q(\u_geo/w_vz_mvp [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [10]),
        .Q(\u_geo/w_vz_mvp [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [11]),
        .Q(\u_geo/w_vz_mvp [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[12] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [12]),
        .Q(\u_geo/w_vz_mvp [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[13] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [13]),
        .Q(\u_geo/w_vz_mvp [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[14] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [14]),
        .Q(\u_geo/w_vz_mvp [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[15] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [15]),
        .Q(\u_geo/w_vz_mvp [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[16] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [16]),
        .Q(\u_geo/w_vz_mvp [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[17] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [17]),
        .Q(\u_geo/w_vz_mvp [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[18] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [18]),
        .Q(\u_geo/w_vz_mvp [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[19] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [19]),
        .Q(\u_geo/w_vz_mvp [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [1]),
        .Q(\u_geo/w_vz_mvp [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[20] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [20]),
        .Q(\u_geo/w_vz_mvp [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[21] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [21]),
        .Q(\u_geo/w_vz_mvp [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [2]),
        .Q(\u_geo/w_vz_mvp [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [3]),
        .Q(\u_geo/w_vz_mvp [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [4]),
        .Q(\u_geo/w_vz_mvp [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [5]),
        .Q(\u_geo/w_vz_mvp [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [6]),
        .Q(\u_geo/w_vz_mvp [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [7]),
        .Q(\u_geo/w_vz_mvp [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [8]),
        .Q(\u_geo/w_vz_mvp [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_vz_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .D(\u_geo/u_geo_matrix/w_add0123_out [9]),
        .Q(\u_geo/w_vz_mvp [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_wait_end_1z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/w_wait_end ),
        .Q(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_wait_end_2z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/r_wait_end_1z ),
        .Q(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/r_wait_end_3z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/r_wait_end_2z ),
        .Q(\u_geo/u_geo_matrix/r_wait_end_3z ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry_n_0 ,\u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry_n_1 ,\u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry_n_2 ,\u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry_n_3 }),
        .CYINIT(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [0]),
        .DI({\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [3:1],_inferred__1_carry_i_1__8_n_0}),
        .O(\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [3:0]),
        .S({_inferred__1_carry_i_2__3_n_0,_inferred__1_carry_i_3__3_n_0,_inferred__1_carry_i_4__3_n_0,_inferred__1_carry_i_5__4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry__0 
       (.CI(\u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]}),
        .O({\u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry__0_n_4 ,\u_geo/u_geo_matrix/u_fadd_m01/norm/_inferred__1_carry__0_n_5 ,\u_geo/u_geo_matrix/u_fadd_m01/norm/f_incdec_return [5:4]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,_inferred__1_carry_i_1__7_n_0,_inferred__1_carry_i_2__15_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[0]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [0]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[10]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [10]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[11]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [11]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[12]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [12]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[13]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [13]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[14]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [14]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_c ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/norm/w_c_exp [0]),
        .Q(\u_geo/u_geo_matrix/w_add01_out [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/norm/w_c_exp [1]),
        .Q(\u_geo/u_geo_matrix/w_add01_out [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/norm/w_c_exp [2]),
        .Q(\u_geo/u_geo_matrix/w_add01_out [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/norm/w_c_exp [3]),
        .Q(\u_geo/u_geo_matrix/w_add01_out [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[1]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [1]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/norm/w_c_exp [4]),
        .Q(\u_geo/u_geo_matrix/w_add01_out [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/r_sign_2z ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [21]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[2]_i_1__6_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [2]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[3]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [3]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[4]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [4]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[5]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [5]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[6]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [6]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[7]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [7]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[8]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [8]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_c_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[9]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add01_out [9]),
        .R(\r_c[21]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_exp_l [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_exp_l [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_exp_l [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_exp_l [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_exp_l [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_1z [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_exp_2z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [10]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [11]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [12]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [13]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [14]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [15]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [5]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [6]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [7]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [8]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f0_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f0 [9]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f0 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [10]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [11]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [12]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [13]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [14]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [15]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [5]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [6]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [7]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [8]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_f1t_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_f1t [9]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_f1t [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [10]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [11]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [12]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [13]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [14]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [15]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [16]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [5]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [6]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [7]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [8]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_mats_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_mats [9]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_mats [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_sign_1z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_sign ),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_sign_1z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_sign_2z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/r_sign_1z ),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_sign_2z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m01/r_sub_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m01/w_sub11_in ),
        .Q(\u_geo/u_geo_matrix/u_fadd_m01/r_sub ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry_n_0 ,\u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry_n_1 ,\u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry_n_2 ,\u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({w_mag_frac_carry_i_1_n_0,w_mag_frac_carry_i_2_n_0,w_mag_frac_carry_i_3_n_0,w_mag_frac_carry_i_4_n_0}),
        .S({w_mag_frac_carry_i_5_n_0,w_mag_frac_carry_i_6_n_0,w_mag_frac_carry_i_7_n_0,w_mag_frac_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry__0 
       (.CI(\u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry_n_0 ),
        .CO({\u_geo/u_geo_matrix/u_fadd_m01/data0 ,\u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry__0_n_1 ,\u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry__0_n_2 ,\u_geo/u_geo_matrix/u_fadd_m01/w_mag_frac_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({w_mag_frac_carry_i_1__0_n_0,w_mag_frac_carry_i_2__0_n_0,w_mag_frac_carry_i_3__0_n_0,w_mag_frac_carry_i_4__0_n_0}),
        .S({w_mag_frac_carry_i_5__0_n_0,w_mag_frac_carry_i_6__0_n_0,w_mag_frac_carry_i_7__0_n_0,w_mag_frac_carry_i_8__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry_n_0 ,\u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry_n_1 ,\u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry_n_2 ,\u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry_n_3 }),
        .CYINIT(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [0]),
        .DI({\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [3:1],_inferred__1_carry_i_1__12_n_0}),
        .O(\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [3:0]),
        .S({_inferred__1_carry_i_2__5_n_0,_inferred__1_carry_i_3__5_n_0,_inferred__1_carry_i_4__5_n_0,_inferred__1_carry_i_5__6_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry__0 
       (.CI(\u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]}),
        .O({\u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry__0_n_4 ,\u_geo/u_geo_matrix/u_fadd_m0123/norm/_inferred__1_carry__0_n_5 ,\u_geo/u_geo_matrix/u_fadd_m0123/norm/f_incdec_return [5:4]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,_inferred__1_carry_i_1__11_n_0,_inferred__1_carry_i_2__17_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[0]_i_1__6_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [0]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[10]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [10]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[11]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [11]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[12]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [12]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[13]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [13]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[14]_i_1__6_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [14]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_c ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/norm/w_c_exp [0]),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/norm/w_c_exp [1]),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/norm/w_c_exp [2]),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/norm/w_c_exp [3]),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[1]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [1]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/norm/w_c_exp [4]),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/r_sign_2z ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [21]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[2]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [2]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[3]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [3]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[4]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [4]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[5]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [5]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[6]_i_1__6_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [6]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[7]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [7]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[8]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [8]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_c_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[9]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add0123_out [9]),
        .R(\r_c[21]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_exp_l [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_exp_l [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_exp_l [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_exp_l [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_exp_l [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_1z [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_exp_2z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [10]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [11]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [12]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [13]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [14]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [15]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [5]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [6]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [7]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [8]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f0_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f0 [9]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f0 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [10]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [11]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [12]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [13]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [14]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [15]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [5]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [6]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [7]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [8]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_f1t_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_f1t [9]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_f1t [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [10]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [11]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [12]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [13]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [14]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [15]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [16]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [5]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [6]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [7]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [8]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_mats_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_mats [9]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_mats [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_sign_1z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_sign ),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_sign_1z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_sign_2z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/r_sign_1z ),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_sign_2z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m0123/r_sub_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m0123/w_sub11_in ),
        .Q(\u_geo/u_geo_matrix/u_fadd_m0123/r_sub ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry_n_0 ,\u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry_n_1 ,\u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry_n_2 ,\u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({w_mag_frac_carry_i_1__3_n_0,w_mag_frac_carry_i_2__3_n_0,w_mag_frac_carry_i_3__3_n_0,w_mag_frac_carry_i_4__3_n_0}),
        .S({w_mag_frac_carry_i_5__3_n_0,w_mag_frac_carry_i_6__3_n_0,w_mag_frac_carry_i_7__3_n_0,w_mag_frac_carry_i_8__3_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry__0 
       (.CI(\u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry_n_0 ),
        .CO({\u_geo/u_geo_matrix/u_fadd_m0123/data0 ,\u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry__0_n_1 ,\u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry__0_n_2 ,\u_geo/u_geo_matrix/u_fadd_m0123/w_mag_frac_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({w_mag_frac_carry_i_1__4_n_0,w_mag_frac_carry_i_2__4_n_0,w_mag_frac_carry_i_3__4_n_0,w_mag_frac_carry_i_4__4_n_0}),
        .S({w_mag_frac_carry_i_5__4_n_0,w_mag_frac_carry_i_6__4_n_0,w_mag_frac_carry_i_7__4_n_0,w_mag_frac_carry_i_8__4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry_n_0 ,\u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry_n_1 ,\u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry_n_2 ,\u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry_n_3 }),
        .CYINIT(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [0]),
        .DI({\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [3:1],_inferred__1_carry_i_1__10_n_0}),
        .O(\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [3:0]),
        .S({_inferred__1_carry_i_2__4_n_0,_inferred__1_carry_i_3__4_n_0,_inferred__1_carry_i_4__4_n_0,_inferred__1_carry_i_5__5_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry__0 
       (.CI(\u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]}),
        .O({\u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry__0_n_4 ,\u_geo/u_geo_matrix/u_fadd_m23/norm/_inferred__1_carry__0_n_5 ,\u_geo/u_geo_matrix/u_fadd_m23/norm/f_incdec_return [5:4]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,_inferred__1_carry_i_1__9_n_0,_inferred__1_carry_i_2__16_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[0]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [0]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[10]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [10]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[11]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [11]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[12]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [12]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[13]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [13]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[14]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [14]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_c ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/norm/w_c_exp [0]),
        .Q(\u_geo/u_geo_matrix/w_add23_out [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/norm/w_c_exp [1]),
        .Q(\u_geo/u_geo_matrix/w_add23_out [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/norm/w_c_exp [2]),
        .Q(\u_geo/u_geo_matrix/w_add23_out [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/norm/w_c_exp [3]),
        .Q(\u_geo/u_geo_matrix/w_add23_out [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[1]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [1]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/norm/w_c_exp [4]),
        .Q(\u_geo/u_geo_matrix/w_add23_out [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/r_sign_2z ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [21]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[2]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [2]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[3]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [3]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[4]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [4]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[5]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [5]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[6]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [6]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[7]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [7]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[8]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [8]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_c_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[9]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_add23_out [9]),
        .R(\r_c[21]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_exp_l [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_exp_l [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_exp_l [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_exp_l [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_exp_l [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_1z [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_exp_2z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [10]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [11]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [12]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [13]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [14]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [15]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [5]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [6]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [7]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [8]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f0_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f0 [9]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f0 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [10]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [11]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [12]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [13]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [14]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [15]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [5]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [6]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [7]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [8]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_f1t_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_f1t [9]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_f1t [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [0]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [10]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [11]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [12]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [13]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [14]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [15]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [16]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [1]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [2]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [3]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [4]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [5]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [6]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [7]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [8]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_mats_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_mats [9]),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_mats [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_sign_1z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_sign ),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_sign_1z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_sign_2z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/r_sign_1z ),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_sign_2z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fadd_m23/r_sub_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fadd_m23/w_sub11_in ),
        .Q(\u_geo/u_geo_matrix/u_fadd_m23/r_sub ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry_n_0 ,\u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry_n_1 ,\u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry_n_2 ,\u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({w_mag_frac_carry_i_1__1_n_0,w_mag_frac_carry_i_2__1_n_0,w_mag_frac_carry_i_3__1_n_0,w_mag_frac_carry_i_4__1_n_0}),
        .S({w_mag_frac_carry_i_5__1_n_0,w_mag_frac_carry_i_6__1_n_0,w_mag_frac_carry_i_7__1_n_0,w_mag_frac_carry_i_8__1_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry__0 
       (.CI(\u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry_n_0 ),
        .CO({\u_geo/u_geo_matrix/u_fadd_m23/data0 ,\u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry__0_n_1 ,\u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry__0_n_2 ,\u_geo/u_geo_matrix/u_fadd_m23/w_mag_frac_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({w_mag_frac_carry_i_1__2_n_0,w_mag_frac_carry_i_2__2_n_0,w_mag_frac_carry_i_3__2_n_0,w_mag_frac_carry_i_4__2_n_0}),
        .S({w_mag_frac_carry_i_5__2_n_0,w_mag_frac_carry_i_6__2_n_0,w_mag_frac_carry_i_7__2_n_0,w_mag_frac_carry_i_8__2_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry_n_0 ,\u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry_n_1 ,\u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry_n_2 ,\u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry_n_3 }),
        .CYINIT(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [0]),
        .DI({\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [3:1],_inferred__1_carry_i_1__0_n_0}),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [3:0]),
        .S({_inferred__1_carry_i_2_n_0,_inferred__1_carry_i_3_n_0,_inferred__1_carry_i_4_n_0,_inferred__1_carry_i_5__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry__0 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]}),
        .O({\u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry__0_n_4 ,\u_geo/u_geo_matrix/u_fmul_m0/norm/_inferred__1_carry__0_n_5 ,\u_geo/u_geo_matrix/u_fmul_m0/norm/f_incdec_return [5:4]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,_inferred__1_carry_i_1_n_0,_inferred__1_carry_i_2__11_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_c),
        .Q(\u_geo/u_geo_matrix/w_m0_out [0]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[10]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [10]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[11]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [11]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[12]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [12]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[13]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [13]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[14]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [14]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_c ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/norm/w_c_exp [0]),
        .Q(\u_geo/u_geo_matrix/w_m0_out [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/norm/w_c_exp [1]),
        .Q(\u_geo/u_geo_matrix/w_m0_out [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/norm/w_c_exp [2]),
        .Q(\u_geo/u_geo_matrix/w_m0_out [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/norm/w_c_exp [3]),
        .Q(\u_geo/u_geo_matrix/w_m0_out [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[1]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [1]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/norm/w_c_exp [4]),
        .Q(\u_geo/u_geo_matrix/w_m0_out [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/r_sign_2z ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [21]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[2]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [2]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[3]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [3]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[4]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [4]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[5]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [5]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[6]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [6]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[7]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [7]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[8]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [8]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_c_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[9]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m0_out [9]),
        .R(\r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[0]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_ ),
        .R(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[1]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_[1] ),
        .R(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[2]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_[2] ),
        .R(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[3]_i_1_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_[3] ),
        .R(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[4]_i_2_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_[4] ),
        .R(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_ ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_[1] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_[2] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_[3] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_1z_reg_n_0_[4] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_ce_tmp_2z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2[3]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m0/p_0_in [1]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m0/p_0_in [0]),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [0]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [10]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [11]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[11]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[7]_i_1_n_0 ),
        .CO(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [11:8]),
        .S(\u_geo/u_geo_matrix/u_fmul_m0/p_0_in [12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [12]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [13]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [14]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [15]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[15]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg [3]),
        .CO({\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[15]_i_1_n_0 ,\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[15]_i_1_n_1 ,\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[15]_i_1_n_2 ,\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [15:12]),
        .S(\u_geo/u_geo_matrix/u_fmul_m0/p_0_in [16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [16]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[16]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[15]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[16]_i_1_n_4 ,\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[16]_i_1_n_5 ,\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[16]_i_1_n_6 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [16]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fmul_m0/p_0_in [17]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [1]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [2]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [3]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[3]_i_1_n_0 ,\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[3]_i_1_n_1 ,\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[3]_i_1_n_2 ,\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fmul_m0/p_0_in [1]}),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [3:0]),
        .S({\u_geo/u_geo_matrix/u_fmul_m0/p_0_in [4:2],\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2[3]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [4]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [5]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [6]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [7]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[7]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[3]_i_1_n_0 ),
        .CO({\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[7]_i_1_n_0 ,\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[7]_i_1_n_1 ,\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[7]_i_1_n_2 ,\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [7:4]),
        .S(\u_geo/u_geo_matrix/u_fmul_m0/p_0_in [8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [8]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp2 [9]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_cf_tmp2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_sign_1z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/w_sign ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_sign_1z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m0/r_sign_2z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m0/r_sign_1z ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m0/r_sign_2z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/w_vx_in }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,w_cf_tmp_i_1_n_0,w_cf_tmp_i_2_n_0,w_cf_tmp_i_3_n_0,w_cf_tmp_i_4_n_0,w_cf_tmp_i_5_n_0,w_cf_tmp_i_6_n_0,w_cf_tmp_i_7_n_0,w_cf_tmp_i_8_n_0,w_cf_tmp_i_9_n_0,w_cf_tmp_i_10_n_0,w_cf_tmp_i_11_n_0,w_cf_tmp_i_12_n_0,w_cf_tmp_i_13_n_0,w_cf_tmp_i_14_n_0,w_cf_tmp_i_15_n_0,w_cf_tmp_i_16_n_0}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const1>__0__0 ),
        .CLK(clk_i),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_58 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_59 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_60 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_61 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_62 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_63 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_64 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_65 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_66 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_67 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_68 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_69 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_70 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_71 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_72 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_73 ,\u_geo/u_geo_matrix/u_fmul_m0/p_0_in ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_92 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_93 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_94 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_95 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_96 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_97 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_98 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_99 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_100 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_101 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_102 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_103 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_104 ,\u_geo/u_geo_matrix/u_fmul_m0/w_cf_tmp_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry_n_0 ,\u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry_n_1 ,\u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry_n_2 ,\u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry_n_3 }),
        .CYINIT(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [0]),
        .DI({\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [3:1],_inferred__1_carry_i_1__2_n_0}),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [3:0]),
        .S({_inferred__1_carry_i_2__0_n_0,_inferred__1_carry_i_3__0_n_0,_inferred__1_carry_i_4__0_n_0,_inferred__1_carry_i_5__1_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry__0 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]}),
        .O({\u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry__0_n_4 ,\u_geo/u_geo_matrix/u_fmul_m1/norm/_inferred__1_carry__0_n_5 ,\u_geo/u_geo_matrix/u_fmul_m1/norm/f_incdec_return [5:4]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,_inferred__1_carry_i_1__1_n_0,_inferred__1_carry_i_2__12_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[0]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [0]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[10]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [10]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[11]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [11]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[12]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [12]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[13]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [13]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[14]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [14]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_c ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/norm/w_c_exp [0]),
        .Q(\u_geo/u_geo_matrix/w_m1_out [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/norm/w_c_exp [1]),
        .Q(\u_geo/u_geo_matrix/w_m1_out [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/norm/w_c_exp [2]),
        .Q(\u_geo/u_geo_matrix/w_m1_out [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/norm/w_c_exp [3]),
        .Q(\u_geo/u_geo_matrix/w_m1_out [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[1]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [1]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/norm/w_c_exp [4]),
        .Q(\u_geo/u_geo_matrix/w_m1_out [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/r_sign_2z ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [21]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[2]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [2]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[3]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [3]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[4]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [4]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[5]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [5]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[6]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [6]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[7]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [7]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[8]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [8]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_c_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[9]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m1_out [9]),
        .R(\r_c[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_ce_tmp_1z),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_ ),
        .R(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[1]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_[1] ),
        .R(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[2]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_[2] ),
        .R(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[3]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_[3] ),
        .R(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[4]_i_2__0_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_[4] ),
        .R(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_ ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_[1] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_[2] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_[3] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_1z_reg_n_0_[4] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_ce_tmp_2z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2[3]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m1/p_0_in [1]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m1/p_0_in [0]),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [0]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [10]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [11]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[11]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[7]_i_1_n_0 ),
        .CO(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [11:8]),
        .S(\u_geo/u_geo_matrix/u_fmul_m1/p_0_in [12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [12]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [13]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [14]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [15]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[15]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg [3]),
        .CO({\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[15]_i_1_n_0 ,\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[15]_i_1_n_1 ,\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[15]_i_1_n_2 ,\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [15:12]),
        .S(\u_geo/u_geo_matrix/u_fmul_m1/p_0_in [16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [16]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[16]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[15]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[16]_i_1_n_4 ,\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[16]_i_1_n_5 ,\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[16]_i_1_n_6 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [16]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fmul_m1/p_0_in [17]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [1]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [2]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [3]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[3]_i_1_n_0 ,\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[3]_i_1_n_1 ,\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[3]_i_1_n_2 ,\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fmul_m1/p_0_in [1]}),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [3:0]),
        .S({\u_geo/u_geo_matrix/u_fmul_m1/p_0_in [4:2],\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2[3]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [4]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [5]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [6]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [7]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[7]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[3]_i_1_n_0 ),
        .CO({\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[7]_i_1_n_0 ,\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[7]_i_1_n_1 ,\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[7]_i_1_n_2 ,\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [7:4]),
        .S(\u_geo/u_geo_matrix/u_fmul_m1/p_0_in [8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [8]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp2 [9]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_cf_tmp2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_sign_1z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/w_sign ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_sign_1z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m1/r_sign_2z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m1/r_sign_1z ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m1/r_sign_2z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/w_vy_in }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,w_cf_tmp_i_1__0_n_0,w_cf_tmp_i_2__0_n_0,w_cf_tmp_i_3__0_n_0,w_cf_tmp_i_4__0_n_0,w_cf_tmp_i_5__0_n_0,w_cf_tmp_i_6__0_n_0,w_cf_tmp_i_7__0_n_0,w_cf_tmp_i_8__0_n_0,w_cf_tmp_i_9__0_n_0,w_cf_tmp_i_10__0_n_0,w_cf_tmp_i_11__0_n_0,w_cf_tmp_i_12__0_n_0,w_cf_tmp_i_13__0_n_0,w_cf_tmp_i_14__0_n_0,w_cf_tmp_i_15__0_n_0,w_cf_tmp_i_16__0_n_0}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const1>__0__0 ),
        .CLK(clk_i),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_58 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_59 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_60 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_61 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_62 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_63 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_64 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_65 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_66 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_67 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_68 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_69 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_70 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_71 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_72 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_73 ,\u_geo/u_geo_matrix/u_fmul_m1/p_0_in ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_92 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_93 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_94 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_95 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_96 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_97 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_98 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_99 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_100 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_101 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_102 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_103 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_104 ,\u_geo/u_geo_matrix/u_fmul_m1/w_cf_tmp_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry_n_0 ,\u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry_n_1 ,\u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry_n_2 ,\u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry_n_3 }),
        .CYINIT(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [0]),
        .DI({\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [3:1],_inferred__1_carry_i_1__4_n_0}),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [3:0]),
        .S({_inferred__1_carry_i_2__1_n_0,_inferred__1_carry_i_3__1_n_0,_inferred__1_carry_i_4__1_n_0,_inferred__1_carry_i_5__2_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry__0 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]}),
        .O({\u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry__0_n_4 ,\u_geo/u_geo_matrix/u_fmul_m2/norm/_inferred__1_carry__0_n_5 ,\u_geo/u_geo_matrix/u_fmul_m2/norm/f_incdec_return [5:4]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,_inferred__1_carry_i_1__3_n_0,_inferred__1_carry_i_2__13_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[0]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [0]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[10]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [10]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[11]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [11]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[12]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [12]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[13]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [13]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[14]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [14]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_c ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/norm/w_c_exp [0]),
        .Q(\u_geo/u_geo_matrix/w_m2_out [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/norm/w_c_exp [1]),
        .Q(\u_geo/u_geo_matrix/w_m2_out [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/norm/w_c_exp [2]),
        .Q(\u_geo/u_geo_matrix/w_m2_out [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/norm/w_c_exp [3]),
        .Q(\u_geo/u_geo_matrix/w_m2_out [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[1]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [1]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/norm/w_c_exp [4]),
        .Q(\u_geo/u_geo_matrix/w_m2_out [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/r_sign_2z ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [21]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[2]_i_1__4_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [2]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[3]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [3]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[4]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [4]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[5]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [5]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[6]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [6]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[7]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [7]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[8]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [8]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_c_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[9]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m2_out [9]),
        .R(\r_c[21]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[0]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_ ),
        .R(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[1]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_[1] ),
        .R(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[2]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_[2] ),
        .R(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[3]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_[3] ),
        .R(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[4]_i_2__1_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_[4] ),
        .R(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_ ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_[1] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_[2] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_[3] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_1z_reg_n_0_[4] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_ce_tmp_2z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2[3]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m2/p_0_in [1]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m2/p_0_in [0]),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [0]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [10]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [11]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[11]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[7]_i_1_n_0 ),
        .CO(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [11:8]),
        .S(\u_geo/u_geo_matrix/u_fmul_m2/p_0_in [12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [12]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [13]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [14]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [15]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[15]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg [3]),
        .CO({\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[15]_i_1_n_0 ,\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[15]_i_1_n_1 ,\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[15]_i_1_n_2 ,\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [15:12]),
        .S(\u_geo/u_geo_matrix/u_fmul_m2/p_0_in [16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [16]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[16]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[15]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[16]_i_1_n_4 ,\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[16]_i_1_n_5 ,\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[16]_i_1_n_6 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [16]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fmul_m2/p_0_in [17]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [1]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [2]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [3]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[3]_i_1_n_0 ,\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[3]_i_1_n_1 ,\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[3]_i_1_n_2 ,\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fmul_m2/p_0_in [1]}),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [3:0]),
        .S({\u_geo/u_geo_matrix/u_fmul_m2/p_0_in [4:2],\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2[3]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [4]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [5]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [6]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [7]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[7]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[3]_i_1_n_0 ),
        .CO({\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[7]_i_1_n_0 ,\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[7]_i_1_n_1 ,\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[7]_i_1_n_2 ,\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [7:4]),
        .S(\u_geo/u_geo_matrix/u_fmul_m2/p_0_in [8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [8]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp2 [9]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_cf_tmp2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_sign_1z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/w_sign ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_sign_1z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m2/r_sign_2z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m2/r_sign_1z ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m2/r_sign_2z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/w_vz_in }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,w_cf_tmp_i_1__1_n_0,w_cf_tmp_i_2__1_n_0,w_cf_tmp_i_3__1_n_0,w_cf_tmp_i_4__1_n_0,w_cf_tmp_i_5__1_n_0,w_cf_tmp_i_6__1_n_0,w_cf_tmp_i_7__1_n_0,w_cf_tmp_i_8__1_n_0,w_cf_tmp_i_9__1_n_0,w_cf_tmp_i_10__1_n_0,w_cf_tmp_i_11__1_n_0,w_cf_tmp_i_12__1_n_0,w_cf_tmp_i_13__1_n_0,w_cf_tmp_i_14__1_n_0,w_cf_tmp_i_15__1_n_0,w_cf_tmp_i_16__1_n_0}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const1>__0__0 ),
        .CLK(clk_i),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_58 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_59 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_60 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_61 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_62 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_63 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_64 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_65 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_66 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_67 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_68 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_69 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_70 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_71 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_72 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_73 ,\u_geo/u_geo_matrix/u_fmul_m2/p_0_in ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_92 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_93 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_94 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_95 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_96 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_97 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_98 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_99 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_100 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_101 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_102 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_103 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_104 ,\u_geo/u_geo_matrix/u_fmul_m2/w_cf_tmp_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry_n_0 ,\u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry_n_1 ,\u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry_n_2 ,\u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry_n_3 }),
        .CYINIT(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [0]),
        .DI({\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [3:1],_inferred__1_carry_i_1__6_n_0}),
        .O(\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [3:0]),
        .S({_inferred__1_carry_i_2__2_n_0,_inferred__1_carry_i_3__2_n_0,_inferred__1_carry_i_4__2_n_0,_inferred__1_carry_i_5__3_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry__0 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]}),
        .O({\u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry__0_n_4 ,\u_geo/u_geo_matrix/u_fmul_m3/norm/_inferred__1_carry__0_n_5 ,\u_geo/u_geo_matrix/u_fmul_m3/norm/f_incdec_return [5:4]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,_inferred__1_carry_i_1__5_n_0,_inferred__1_carry_i_2__14_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[0]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [0]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[10]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [10]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[11]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [11]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[12]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [12]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[13]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [13]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[14]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [14]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_c ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/norm/w_c_exp [0]),
        .Q(\u_geo/u_geo_matrix/w_m3_out [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/norm/w_c_exp [1]),
        .Q(\u_geo/u_geo_matrix/w_m3_out [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/norm/w_c_exp [2]),
        .Q(\u_geo/u_geo_matrix/w_m3_out [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/norm/w_c_exp [3]),
        .Q(\u_geo/u_geo_matrix/w_m3_out [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[1]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [1]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/norm/w_c_exp [4]),
        .Q(\u_geo/u_geo_matrix/w_m3_out [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/r_sign_2z ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [21]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[2]_i_1__5_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [2]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[3]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [3]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[4]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [4]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[5]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [5]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[6]_i_1__3_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [6]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[7]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [7]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[8]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [8]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_c_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[9]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/w_m3_out [9]),
        .R(\r_c[21]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[0]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[1]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[2]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[3]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp_1z[4]_i_1__2_n_0 ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_ ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_[1] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_[2] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_[3] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_1z_reg_n_0_[4] ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_ce_tmp_2z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2[3]_i_5 
       (.I0(\u_geo/u_geo_matrix/u_fmul_m3/p_0_in [1]),
        .I1(\u_geo/u_geo_matrix/u_fmul_m3/p_0_in [0]),
        .O(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [0]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [10]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [11]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[11]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[7]_i_1_n_0 ),
        .CO(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [11:8]),
        .S(\u_geo/u_geo_matrix/u_fmul_m3/p_0_in [12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [12]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [13]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [14]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [15]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[15]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg [3]),
        .CO({\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[15]_i_1_n_0 ,\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[15]_i_1_n_1 ,\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[15]_i_1_n_2 ,\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [15:12]),
        .S(\u_geo/u_geo_matrix/u_fmul_m3/p_0_in [16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [16]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[16]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[15]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[16]_i_1_n_4 ,\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[16]_i_1_n_5 ,\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[16]_i_1_n_6 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [16]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fmul_m3/p_0_in [17]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [1]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [2]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [3]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[3]_i_1_n_0 ,\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[3]_i_1_n_1 ,\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[3]_i_1_n_2 ,\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_matrix/u_fmul_m3/p_0_in [1]}),
        .O(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [3:0]),
        .S({\u_geo/u_geo_matrix/u_fmul_m3/p_0_in [4:2],\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2[3]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [4]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [5]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [6]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [7]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[7]_i_1 
       (.CI(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[3]_i_1_n_0 ),
        .CO({\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[7]_i_1_n_0 ,\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[7]_i_1_n_1 ,\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[7]_i_1_n_2 ,\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [7:4]),
        .S(\u_geo/u_geo_matrix/u_fmul_m3/p_0_in [8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [8]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp2 [9]),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_cf_tmp2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_sign_1z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_sign_1z_i_1__5_n_0),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_sign_1z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_matrix/u_fmul_m3/r_sign_2z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_matrix/u_fmul_m3/r_sign_1z ),
        .Q(\u_geo/u_geo_matrix/u_fmul_m3/r_sign_2z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,w_cf_tmp_i_1__2_n_0,w_cf_tmp_i_2__2_n_0,w_cf_tmp_i_3__2_n_0,w_cf_tmp_i_4__2_n_0,w_cf_tmp_i_5__2_n_0,w_cf_tmp_i_6__2_n_0,w_cf_tmp_i_7__2_n_0,w_cf_tmp_i_8__2_n_0,w_cf_tmp_i_9__2_n_0,w_cf_tmp_i_10__2_n_0,w_cf_tmp_i_11__2_n_0,w_cf_tmp_i_12__2_n_0,w_cf_tmp_i_13__2_n_0,w_cf_tmp_i_14__2_n_0,w_cf_tmp_i_15__2_n_0,w_cf_tmp_i_16__2_n_0}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const1>__0__0 ),
        .CLK(clk_i),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_58 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_59 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_60 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_61 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_62 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_63 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_64 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_65 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_66 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_67 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_68 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_69 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_70 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_71 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_72 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_73 ,\u_geo/u_geo_matrix/u_fmul_m3/p_0_in ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_92 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_93 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_94 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_95 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_96 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_97 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_98 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_99 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_100 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_101 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_102 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_103 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_104 ,\u_geo/u_geo_matrix/u_fmul_m3/w_cf_tmp_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/FSM_onehot_r_state_reg[0] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[5]_i_1_n_0 ),
        .D(\FSM_onehot_r_state[0]_i_1_n_0 ),
        .Q(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_ ),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/FSM_onehot_r_state_reg[1] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[5]_i_1_n_0 ),
        .D(\FSM_onehot_r_state[1]_i_1_n_0 ),
        .Q(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/FSM_onehot_r_state_reg[2] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[5]_i_1_n_0 ),
        .D(\FSM_onehot_r_state[2]_i_1_n_0 ),
        .Q(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/FSM_onehot_r_state_reg[3] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[5]_i_1_n_0 ),
        .D(\FSM_onehot_r_state[3]_i_1_n_0 ),
        .Q(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/FSM_onehot_r_state_reg[4] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[5]_i_1_n_0 ),
        .D(\FSM_onehot_r_state[4]_i_1_n_0 ),
        .Q(\u_geo/w_en_dma ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/FSM_onehot_r_state_reg[5] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[5]_i_1_n_0 ),
        .D(\FSM_onehot_r_state[5]_i_2_n_0 ),
        .Q(\u_geo/w_dma_end ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \u_geo/u_geo_mem/o_req_m 
       (.I0(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[1] ),
        .I2(\u_geo/u_geo_mem/FSM_onehot_r_state_reg_n_0_[2] ),
        .O(w_req_geo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[0] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [0]),
        .Q(w_adrs_geo[2]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[10] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [10]),
        .Q(w_adrs_geo[12]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[11] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [11]),
        .Q(w_adrs_geo[13]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[12] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [12]),
        .Q(w_adrs_geo[14]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2 
       (.CI(\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_0 ),
        .CO(\u_geo/u_geo_mem/r_cur_adrs_reg ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2_n_4 ,\u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2_n_5 ,\u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2_n_6 ,\u_geo/u_geo_mem/r_cur_adrs_reg[12]_i_2_n_7 }),
        .S(w_adrs_geo[14:11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[13] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [13]),
        .Q(w_adrs_geo[15]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[14] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [14]),
        .Q(w_adrs_geo[16]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[15] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [15]),
        .Q(w_adrs_geo[17]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[16] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [16]),
        .Q(w_adrs_geo[18]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2 
       (.CI(\u_geo/u_geo_mem/r_cur_adrs_reg [3]),
        .CO({\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_0 ,\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_1 ,\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_2 ,\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_4 ,\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_5 ,\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_6 ,\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_7 }),
        .S(w_adrs_geo[18:15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[17] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [17]),
        .Q(w_adrs_geo[19]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[18] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [18]),
        .Q(w_adrs_geo[20]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[19] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [19]),
        .Q(w_adrs_geo[21]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[1] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [1]),
        .Q(w_adrs_geo[3]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[20] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [20]),
        .Q(w_adrs_geo[22]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2 
       (.CI(\u_geo/u_geo_mem/r_cur_adrs_reg[16]_i_2_n_0 ),
        .CO({\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_0 ,\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_1 ,\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_2 ,\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_4 ,\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_5 ,\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_6 ,\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_7 }),
        .S(w_adrs_geo[22:19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[21] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [21]),
        .Q(w_adrs_geo[23]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[22] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [22]),
        .Q(w_adrs_geo[24]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[23] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [23]),
        .Q(w_adrs_geo[25]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[24] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [24]),
        .Q(w_adrs_geo[26]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2 
       (.CI(\u_geo/u_geo_mem/r_cur_adrs_reg[20]_i_2_n_0 ),
        .CO({\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_0 ,\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_1 ,\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_2 ,\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_4 ,\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_5 ,\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_6 ,\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_7 }),
        .S(w_adrs_geo[26:23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[25] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [25]),
        .Q(w_adrs_geo[27]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[26] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [26]),
        .Q(w_adrs_geo[28]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[27] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [27]),
        .Q(w_adrs_geo[29]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[28] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [28]),
        .Q(w_adrs_geo[30]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2 
       (.CI(\u_geo/u_geo_mem/r_cur_adrs_reg[24]_i_2_n_0 ),
        .CO({\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_0 ,\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_1 ,\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_2 ,\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_4 ,\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_5 ,\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_6 ,\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_7 }),
        .S(w_adrs_geo[30:27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[29] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [29]),
        .Q(w_adrs_geo[31]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_mem/r_cur_adrs_reg[29]_i_2 
       (.CI(\u_geo/u_geo_mem/r_cur_adrs_reg[28]_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_mem/r_cur_adrs_reg[29]_i_2_n_4 ,\u_geo/u_geo_mem/r_cur_adrs_reg[29]_i_2_n_5 ,\u_geo/u_geo_mem/r_cur_adrs_reg[29]_i_2_n_6 ,\u_geo/u_geo_mem/r_cur_adrs_reg[29]_i_2_n_7 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,w_adrs_geo[31]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[2] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [2]),
        .Q(w_adrs_geo[4]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[3] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [3]),
        .Q(w_adrs_geo[5]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[4] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [4]),
        .Q(w_adrs_geo[6]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_0 ,\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_1 ,\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_2 ,\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_3 }),
        .CYINIT(w_adrs_geo[2]),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_4 ,\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_5 ,\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_6 ,\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_7 }),
        .S(w_adrs_geo[6:3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[5] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [5]),
        .Q(w_adrs_geo[7]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[6] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [6]),
        .Q(w_adrs_geo[8]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[7] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [7]),
        .Q(w_adrs_geo[9]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[8] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [8]),
        .Q(w_adrs_geo[10]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2 
       (.CI(\u_geo/u_geo_mem/r_cur_adrs_reg[4]_i_2_n_0 ),
        .CO({\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_0 ,\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_1 ,\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_2 ,\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_4 ,\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_5 ,\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_6 ,\u_geo/u_geo_mem/r_cur_adrs_reg[8]_i_2_n_7 }),
        .S(w_adrs_geo[10:7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_cur_adrs_reg[9] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_cur_adrs [9]),
        .Q(w_adrs_geo[11]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[0] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(r_size),
        .Q(\u_geo/u_geo_mem/r_size__0 [0]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[10] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [10]),
        .Q(\u_geo/u_geo_mem/r_size__0 [10]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[11] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [11]),
        .Q(\u_geo/u_geo_mem/r_size__0 [11]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[12] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [12]),
        .Q(\u_geo/u_geo_mem/r_size__0 [12]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[13] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [13]),
        .Q(\u_geo/u_geo_mem/r_size__0 [13]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[14] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [14]),
        .Q(\u_geo/u_geo_mem/r_size__0 [14]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[15] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [15]),
        .Q(\u_geo/u_geo_mem/r_size__0 [15]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[1] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [1]),
        .Q(\u_geo/u_geo_mem/r_size__0 [1]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[2] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [2]),
        .Q(\u_geo/u_geo_mem/r_size__0 [2]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[3] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [3]),
        .Q(\u_geo/u_geo_mem/r_size__0 [3]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[4] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [4]),
        .Q(\u_geo/u_geo_mem/r_size__0 [4]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[5] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [5]),
        .Q(\u_geo/u_geo_mem/r_size__0 [5]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[6] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [6]),
        .Q(\u_geo/u_geo_mem/r_size__0 [6]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[7] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [7]),
        .Q(\u_geo/u_geo_mem/r_size__0 [7]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[8] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [8]),
        .Q(\u_geo/u_geo_mem/r_size__0 [8]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_size_reg[9] 
       (.C(clk_i),
        .CE(\r_size[15]_i_1_n_0 ),
        .D(\u_geo/u_geo_mem/r_size [9]),
        .Q(\u_geo/u_geo_mem/r_size__0 [9]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[3]_i_1_n_7 ),
        .Q(\u_geo/w_vx_dma [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[11]_i_1_n_5 ),
        .Q(\u_geo/w_vx_dma [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[11]_i_1_n_4 ),
        .Q(\u_geo/w_vx_dma [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[12] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[14]_i_1_n_7 ),
        .Q(\u_geo/w_vx_dma [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[13] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[14]_i_1_n_6 ),
        .Q(\u_geo/w_vx_dma [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[14] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[14]_i_1_n_5 ),
        .Q(\u_geo/w_vx_dma [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[15] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\u_geo/u_geo_mem/w_f22 [15]),
        .Q(\u_geo/w_vx_dma [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[16] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\u_geo/u_geo_mem/w_f22 [16]),
        .Q(\u_geo/w_vx_dma [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[17] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\u_geo/u_geo_mem/w_f22 [17]),
        .Q(\u_geo/w_vx_dma [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[18] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\u_geo/u_geo_mem/w_f22 [18]),
        .Q(\u_geo/w_vx_dma [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[19] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\u_geo/u_geo_mem/w_f22 [19]),
        .Q(\u_geo/w_vx_dma [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[3]_i_1_n_6 ),
        .Q(\u_geo/w_vx_dma [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[20] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\u_geo/u_geo_mem/w_f22 [20]),
        .Q(\u_geo/w_vx_dma [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[21] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(m_wb_dat_i[31]),
        .Q(\u_geo/w_vx_dma [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[3]_i_1_n_5 ),
        .Q(\u_geo/w_vx_dma [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[3]_i_1_n_4 ),
        .Q(\u_geo/w_vx_dma [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[7]_i_1_n_7 ),
        .Q(\u_geo/w_vx_dma [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[7]_i_1_n_6 ),
        .Q(\u_geo/w_vx_dma [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[7]_i_1_n_5 ),
        .Q(\u_geo/w_vx_dma [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[7]_i_1_n_4 ),
        .Q(\u_geo/w_vx_dma [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[11]_i_1_n_7 ),
        .Q(\u_geo/w_vx_dma [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vx_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vx ),
        .D(\r_vx_reg[11]_i_1_n_6 ),
        .Q(\u_geo/w_vx_dma [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[3]_i_1_n_7 ),
        .Q(\u_geo/w_vy_dma [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[11]_i_1_n_5 ),
        .Q(\u_geo/w_vy_dma [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[11]_i_1_n_4 ),
        .Q(\u_geo/w_vy_dma [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[12] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[14]_i_1_n_7 ),
        .Q(\u_geo/w_vy_dma [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[13] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[14]_i_1_n_6 ),
        .Q(\u_geo/w_vy_dma [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[14] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[14]_i_1_n_5 ),
        .Q(\u_geo/w_vy_dma [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[15] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\u_geo/u_geo_mem/w_f22 [15]),
        .Q(\u_geo/w_vy_dma [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[16] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\u_geo/u_geo_mem/w_f22 [16]),
        .Q(\u_geo/w_vy_dma [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[17] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\u_geo/u_geo_mem/w_f22 [17]),
        .Q(\u_geo/w_vy_dma [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[18] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\u_geo/u_geo_mem/w_f22 [18]),
        .Q(\u_geo/w_vy_dma [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[19] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\u_geo/u_geo_mem/w_f22 [19]),
        .Q(\u_geo/w_vy_dma [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[3]_i_1_n_6 ),
        .Q(\u_geo/w_vy_dma [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[20] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\u_geo/u_geo_mem/w_f22 [20]),
        .Q(\u_geo/w_vy_dma [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[21] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(m_wb_dat_i[31]),
        .Q(\u_geo/w_vy_dma [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[3]_i_1_n_5 ),
        .Q(\u_geo/w_vy_dma [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[3]_i_1_n_4 ),
        .Q(\u_geo/w_vy_dma [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[7]_i_1_n_7 ),
        .Q(\u_geo/w_vy_dma [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[7]_i_1_n_6 ),
        .Q(\u_geo/w_vy_dma [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[7]_i_1_n_5 ),
        .Q(\u_geo/w_vy_dma [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[7]_i_1_n_4 ),
        .Q(\u_geo/w_vy_dma [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[11]_i_1_n_7 ),
        .Q(\u_geo/w_vy_dma [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vy_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vy ),
        .D(\r_vx_reg[11]_i_1_n_6 ),
        .Q(\u_geo/w_vy_dma [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[3]_i_1_n_7 ),
        .Q(\u_geo/w_vz_dma [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[11]_i_1_n_5 ),
        .Q(\u_geo/w_vz_dma [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[11]_i_1_n_4 ),
        .Q(\u_geo/w_vz_dma [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[12] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[14]_i_1_n_7 ),
        .Q(\u_geo/w_vz_dma [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[13] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[14]_i_1_n_6 ),
        .Q(\u_geo/w_vz_dma [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[14] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[14]_i_1_n_5 ),
        .Q(\u_geo/w_vz_dma [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[15] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\u_geo/u_geo_mem/w_f22 [15]),
        .Q(\u_geo/w_vz_dma [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[16] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\u_geo/u_geo_mem/w_f22 [16]),
        .Q(\u_geo/w_vz_dma [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[17] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\u_geo/u_geo_mem/w_f22 [17]),
        .Q(\u_geo/w_vz_dma [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[18] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\u_geo/u_geo_mem/w_f22 [18]),
        .Q(\u_geo/w_vz_dma [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[19] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\u_geo/u_geo_mem/w_f22 [19]),
        .Q(\u_geo/w_vz_dma [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[3]_i_1_n_6 ),
        .Q(\u_geo/w_vz_dma [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[20] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\u_geo/u_geo_mem/w_f22 [20]),
        .Q(\u_geo/w_vz_dma [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[21] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(m_wb_dat_i[31]),
        .Q(\u_geo/w_vz_dma [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[3]_i_1_n_5 ),
        .Q(\u_geo/w_vz_dma [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[3]_i_1_n_4 ),
        .Q(\u_geo/w_vz_dma [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[7]_i_1_n_7 ),
        .Q(\u_geo/w_vz_dma [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[7]_i_1_n_6 ),
        .Q(\u_geo/w_vz_dma [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[7]_i_1_n_5 ),
        .Q(\u_geo/w_vz_dma [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[7]_i_1_n_4 ),
        .Q(\u_geo/w_vz_dma [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[11]_i_1_n_7 ),
        .Q(\u_geo/w_vz_dma [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_mem/r_vz_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_mem/r_vz ),
        .D(\r_vx_reg[11]_i_1_n_6 ),
        .Q(\u_geo/w_vz_dma [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/FSM_sequential_r_state_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[0]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/r_state [0]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/FSM_sequential_r_state_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[1]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/r_state [1]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/FSM_sequential_r_state_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[2]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/r_state [2]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[0] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_ ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[10] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[10] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[11] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[11] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[12] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[12] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[13] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[13] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[14] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[14] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[15] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[15] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_b_exp [0]),
        .Q(\u_geo/u_geo_persdiv/r_ivw [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_b_exp [1]),
        .Q(\u_geo/u_geo_persdiv/r_ivw [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_b_exp [2]),
        .Q(\u_geo/u_geo_persdiv/r_ivw [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_b_exp [3]),
        .Q(\u_geo/u_geo_persdiv/r_ivw [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[1] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[1] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_b_exp [4]),
        .Q(\u_geo/u_geo_persdiv/r_ivw [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ivw[21]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[2] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[2] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[3] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[3] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[4] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[4] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[5] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[5] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[6] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[6] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[7] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[7] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[8] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[8] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_ivw_reg[9] 
       (.C(clk_i),
        .CE(r_ivw),
        .D(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[9] ),
        .Q(\u_geo/u_geo_persdiv/r_ivw [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_outcode_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/w_state_pd ),
        .D(\u_geo/w_outcode_clip [0]),
        .Q(\u_geo/w_outcode_pdiv [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_outcode_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/w_state_pd ),
        .D(\u_geo/w_outcode_clip [1]),
        .Q(\u_geo/w_outcode_pdiv [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_outcode_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/w_state_pd ),
        .D(\u_geo/w_outcode_clip [2]),
        .Q(\u_geo/w_outcode_pdiv [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_outcode_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/w_state_pd ),
        .D(\u_geo/w_outcode_clip [3]),
        .Q(\u_geo/w_outcode_pdiv [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_outcode_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/w_state_pd ),
        .D(\u_geo/w_outcode_clip [4]),
        .Q(\u_geo/w_outcode_pdiv [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_outcode_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/w_state_pd ),
        .D(\u_geo/w_outcode_clip [5]),
        .Q(\u_geo/w_outcode_pdiv [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[0] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(r_vx),
        .Q(\u_geo/w_vx_pdiv [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[10] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[10]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[11] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[11]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[12] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[12]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[13] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[13]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[14] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[14]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[15] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[15]_i_1__0_n_0 ),
        .Q(\u_geo/w_vx_pdiv [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[16] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[16]_i_1__0_n_0 ),
        .Q(\u_geo/w_vx_pdiv [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[17] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[17]_i_1__0_n_0 ),
        .Q(\u_geo/w_vx_pdiv [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[18] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[18]_i_1__0_n_0 ),
        .Q(\u_geo/w_vx_pdiv [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[19] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[19]_i_1__0_n_0 ),
        .Q(\u_geo/w_vx_pdiv [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[1] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[1]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[20] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[20]_i_1__0_n_0 ),
        .Q(\u_geo/w_vx_pdiv [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[21] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[21]_i_2_n_0 ),
        .Q(\u_geo/w_vx_pdiv [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[2] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[2]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[3] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[3]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[4] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[4]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[5] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[5]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[6] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[6]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[7] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[7]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[8] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[8]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vx_reg[9] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__0_n_0 ),
        .D(\r_vx[9]_i_1_n_0 ),
        .Q(\u_geo/w_vx_pdiv [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[0] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(r_vy),
        .Q(\u_geo/w_vy_pdiv [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[10] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[10]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[11] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[11]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[12] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[12]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[13] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[13]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[14] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[14]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[15] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[15]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[16] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[16]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[17] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[17]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[18] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[18]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[19] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[19]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[1] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[1]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[20] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[20]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[21] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[21]_i_2_n_0 ),
        .Q(\u_geo/w_vy_pdiv [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[2] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[2]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[3] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[3]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[4] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[4]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[5] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[5]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[6] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[6]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[7] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[7]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[8] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[8]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/r_vy_reg[9] 
       (.C(clk_i),
        .CE(\r_vy[21]_i_1__0_n_0 ),
        .D(\r_vy[9]_i_1_n_0 ),
        .Q(\u_geo/w_vy_pdiv [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry_n_0 ,\u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry_n_1 ,\u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry_n_2 ,\u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry_n_3 }),
        .CYINIT(\u_geo/u_geo_persdiv/r_ce_tmp_2z [0]),
        .DI({\u_geo/u_geo_persdiv/r_ce_tmp_2z [3:1],_inferred__1_carry_i_1__16_n_0}),
        .O(\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [3:0]),
        .S({_inferred__1_carry_i_2__7_n_0,_inferred__1_carry_i_3__7_n_0,_inferred__1_carry_i_4__7_n_0,_inferred__1_carry_i_5__8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry__0 
       (.CI(\u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]}),
        .O({\u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry__0_n_4 ,\u_geo/u_geo_persdiv/u_fmul/norm/_inferred__1_carry__0_n_5 ,\u_geo/u_geo_persdiv/u_fmul/norm/f_incdec_return [5:4]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,_inferred__1_carry_i_1__15_n_0,_inferred__1_carry_i_2__19_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[0]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_ ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[10]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[10] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[11]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[11] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[12]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[12] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[13]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[13] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[14]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[14] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_fmul/w_c ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_fmul/norm/w_c_exp [0]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_fmul/norm/w_c_exp [1]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_fmul/norm/w_c_exp [2]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_fmul/norm/w_c_exp [3]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[1]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[1] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_fmul/norm/w_c_exp [4]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_fmul/r_sign_2z ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[21] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[2]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[2] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[3]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[3] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[4]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[4] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[5]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[5] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[6]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[6] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[7]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[7] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[8]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[8] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_c_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[9]_i_1__7_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_c_reg_n_0_[9] ),
        .R(\u_fmul/r_c[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_1z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_fmul/r_ce_tmp_1z[0]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp_1z [0]),
        .R(\u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_1z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_fmul/r_ce_tmp_1z[1]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp_1z [1]),
        .R(\u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_1z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_fmul/r_ce_tmp_1z[2]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp_1z [2]),
        .R(\u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_1z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_fmul/r_ce_tmp_1z[3]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp_1z [3]),
        .R(\u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_1z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_fmul/r_ce_tmp_1z[4]_i_2_n_0 ),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp_1z [4]),
        .R(\u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_2z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/r_ce_tmp_1z [0]),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp_2z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_2z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/r_ce_tmp_1z [1]),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp_2z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_2z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/r_ce_tmp_1z [2]),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp_2z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_2z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/r_ce_tmp_1z [3]),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp_2z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_ce_tmp_2z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/r_ce_tmp_1z [4]),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp_2z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2[3]_i_5 
       (.I0(\u_geo/u_geo_persdiv/p_0_in [1]),
        .I1(\u_geo/u_geo_persdiv/p_0_in [0]),
        .O(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [0]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [10]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [11]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[11]_i_1 
       (.CI(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[7]_i_1_n_0 ),
        .CO(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_persdiv/w_cf_tmp2 [11:8]),
        .S(\u_geo/u_geo_persdiv/p_0_in [12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [12]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [13]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [14]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [15]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[15]_i_1 
       (.CI(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg [3]),
        .CO({\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[15]_i_1_n_0 ,\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[15]_i_1_n_1 ,\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[15]_i_1_n_2 ,\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_persdiv/w_cf_tmp2 [15:12]),
        .S(\u_geo/u_geo_persdiv/p_0_in [16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [16]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[16]_i_1 
       (.CI(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[15]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[16]_i_1_n_4 ,\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[16]_i_1_n_5 ,\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[16]_i_1_n_6 ,\u_geo/u_geo_persdiv/w_cf_tmp2 [16]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_persdiv/p_0_in [17]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [1]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [2]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [3]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[3]_i_1_n_0 ,\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[3]_i_1_n_1 ,\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[3]_i_1_n_2 ,\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_persdiv/p_0_in [1]}),
        .O(\u_geo/u_geo_persdiv/w_cf_tmp2 [3:0]),
        .S({\u_geo/u_geo_persdiv/p_0_in [4:2],\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2[3]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [4]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [5]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [6]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [7]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[7]_i_1 
       (.CI(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[3]_i_1_n_0 ),
        .CO({\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[7]_i_1_n_0 ,\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[7]_i_1_n_1 ,\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[7]_i_1_n_2 ,\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_persdiv/w_cf_tmp2 [7:4]),
        .S(\u_geo/u_geo_persdiv/p_0_in [8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [8]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/w_cf_tmp2 [9]),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_cf_tmp2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_sign_1z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_fmul/w_sign ),
        .Q(\u_geo/u_geo_persdiv/r_sign_1z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_fmul/r_sign_2z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/r_sign_1z ),
        .Q(\u_geo/u_geo_persdiv/u_fmul/r_sign_2z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \u_geo/u_geo_persdiv/u_fmul/w_cf_tmp 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_persdiv/w_fmul_a }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,w_cf_tmp_i_1__3_n_0,w_cf_tmp_i_2__3_n_0,w_cf_tmp_i_3__3_n_0,w_cf_tmp_i_4__3_n_0,w_cf_tmp_i_5__3_n_0,w_cf_tmp_i_6__3_n_0,w_cf_tmp_i_7__3_n_0,w_cf_tmp_i_8__3_n_0,w_cf_tmp_i_9__3_n_0,w_cf_tmp_i_10__3_n_0,w_cf_tmp_i_11__3_n_0,w_cf_tmp_i_12__3_n_0,w_cf_tmp_i_13__3_n_0,w_cf_tmp_i_14__3_n_0,w_cf_tmp_i_15__3_n_0,w_cf_tmp_i_16__3_n_0}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const1>__0__0 ),
        .CLK(clk_i),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_58 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_59 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_60 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_61 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_62 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_63 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_64 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_65 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_66 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_67 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_68 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_69 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_70 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_71 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_72 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_73 ,\u_geo/u_geo_persdiv/p_0_in ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_92 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_93 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_94 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_95 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_96 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_97 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_98 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_99 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_100 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_101 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_102 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_103 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_104 ,\u_geo/u_geo_persdiv/u_fmul/w_cf_tmp_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[16]_i_1 
       (.I0(g0_b16_n_0),
        .I1(g1_b16_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[17]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[17]_i_1 
       (.I0(g0_b17_n_0),
        .I1(g1_b17_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[17]_i_1_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[18]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[18]_i_1 
       (.I0(g0_b18_n_0),
        .I1(g1_b18_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[18]_i_1_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[19]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[19]_i_1 
       (.I0(g0_b19_n_0),
        .I1(g1_b19_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[19]_i_1_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[20]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[20]_i_1 
       (.I0(g0_b20_n_0),
        .I1(g1_b20_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[20]_i_1_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[21]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[21]_i_1 
       (.I0(g0_b21_n_0),
        .I1(g1_b21_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[21]_i_1_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[22] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[22]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[22]_i_1 
       (.I0(g0_b22_n_0),
        .I1(g1_b22_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[22]_i_1_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[23] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[23]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[23]_i_1 
       (.I0(g0_b23_n_0),
        .I1(g1_b23_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[23]_i_1_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[24] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[24]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[24]_i_1 
       (.I0(g0_b24_n_0),
        .I1(g1_b24_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[24]_i_1_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[25] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[25]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[25]_i_1 
       (.I0(g0_b25_n_0),
        .I1(g1_b25_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[25]_i_1_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[26] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[26]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[26]_i_1 
       (.I0(g0_b26_n_0),
        .I1(g1_b26_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[26]_i_1_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[27] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[27]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[27]_i_1 
       (.I0(g0_b27_n_0),
        .I1(g1_b27_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[27]_i_1_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[28] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[28]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[28]_i_1 
       (.I0(g0_b28_n_0),
        .I1(g1_b28_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[28]_i_1_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[29] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[29]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[30] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_frcp/frcp_rom/r_c ),
        .Q(\u_geo/u_geo_persdiv/w_rom_base [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[31]_inv 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[31]_inv_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[31]_inv_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_2 
       (.I0(\u_geo/w_vw_clip [14]),
        .I1(g0_b7_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_3 
       (.I0(g0_b6_n_0),
        .I1(g1_b6_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_3_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_4 
       (.I0(g0_b5_n_0),
        .I1(g1_b5_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_4_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_5 
       (.I0(g0_b4_n_0),
        .I1(g1_b4_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_5_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_6 
       (.I0(g0_b3_n_0),
        .I1(g1_b3_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_6_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_7 
       (.I0(g0_b2_n_0),
        .I1(g1_b2_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_7_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_8 
       (.I0(g0_b1_n_0),
        .I1(g1_b1_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_8_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_9 
       (.I0(g0_b0_n_0),
        .I1(g1_b0_n_0),
        .O(\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_9_n_0 ),
        .S(\u_geo/w_vw_clip [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_a_sign_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/w_vw_clip [21]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_a_sign ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [0]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_ ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [10]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[10] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [11]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[11] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [12]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[12] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [13]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[13] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [14]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[14] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [15]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[15] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [0]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[16] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [1]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[17] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [2]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[18] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [3]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[19] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [1]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[1] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/norm/w_c_exp [4]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[20] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [21]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[21] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [2]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[2] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [3]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[3] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [4]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[4] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [5]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[5] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [6]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[6] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [7]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[7] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [8]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[8] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_c_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_persdiv/u_frcp/w_c [9]),
        .Q(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[9] ),
        .R(\u_geo/u_geo_persdiv/u_frcp/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_ce_tmp_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/w_vw_clip [16]),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_ce_tmp_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_ce_tmp),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_ce_tmp_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp[2]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_ce_tmp_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp[3]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_persdiv/u_frcp/r_ce_tmp_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_ce_tmp[4]_i_1_n_0 ),
        .Q(\u_geo/u_geo_persdiv/r_ce_tmp [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry_n_0 ,\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry_n_1 ,\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry_n_2 ,\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI(\u_geo/u_geo_persdiv/w_rom_base [3:0]),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [3:0]),
        .S({w_cf_tmp_carry_i_1__2_n_0,w_cf_tmp_carry_i_2__2_n_0,w_cf_tmp_carry_i_3__2_n_0,w_cf_tmp_carry_i_4__1_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__0 
       (.CI(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry_n_0 ),
        .CO({\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__0_n_0 ,\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__0_n_1 ,\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__0_n_2 ,\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_persdiv/w_rom_base [7:4]),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [7:4]),
        .S({w_cf_tmp_carry_i_1__1_n_0,w_cf_tmp_carry_i_2__1_n_0,w_cf_tmp_carry_i_3__1_n_0,w_cf_tmp_carry_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__1 
       (.CI(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__0_n_0 ),
        .CO({\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__1_n_0 ,\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__1_n_1 ,\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__1_n_2 ,\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_geo/u_geo_persdiv/w_rom_base [11:8]),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [11:8]),
        .S({w_cf_tmp_carry_i_1__0_n_0,w_cf_tmp_carry_i_2__0_n_0,w_cf_tmp_carry_i_3__0_n_0,w_cf_tmp_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__2 
       (.CI(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp_carry__1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\u_geo/u_geo_persdiv/w_rom_base [14:12]}),
        .O(\u_geo/u_geo_persdiv/u_frcp/w_cf_tmp__45 [15:12]),
        .S({\u_geo/u_geo_persdiv/u_frcp/frcp_rom/r_c_reg[31]_inv_n_0 ,w_cf_tmp_carry_i_1_n_0,w_cf_tmp_carry_i_2_n_0,w_cf_tmp_carry_i_3_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(1),
    .BREG(1),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \u_geo/u_geo_persdiv/u_frcp/w_rom_correct 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,w_rom_correct_i_1_n_0,\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_2_n_0 ,\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_3_n_0 ,\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_4_n_0 ,\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_5_n_0 ,\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_6_n_0 ,\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_7_n_0 ,\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_8_n_0 ,\u_geo/u_geo_persdiv/u_frcp/frcp_rom/w_rom_correct_i_9_n_0 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/w_vw_clip [7:0]}),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const1>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(clk_i),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_58 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_59 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_60 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_61 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_62 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_63 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_64 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_65 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_66 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_67 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_68 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_69 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_70 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_71 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_72 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_73 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_74 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_75 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_76 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_77 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_78 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_79 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_80 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_81 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_82 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_83 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_84 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_85 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_86 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_87 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_88 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_89 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_90 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_91 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_92 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_93 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_94 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_95 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_96 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_97 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_98 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_99 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_100 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_101 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_102 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_103 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_104 ,\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/FSM_onehot_r_state_reg[0] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[6]_i_1_n_0 ),
        .D(FSM_onehot_r_state),
        .Q(\u_geo/w_state_if ),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/FSM_onehot_r_state_reg[1] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[6]_i_1_n_0 ),
        .D(\u_geo/w_state_if ),
        .Q(\u_geo/u_geo_tri/w_set_v0_y ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/FSM_onehot_r_state_reg[2] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[6]_i_1_n_0 ),
        .D(\FSM_onehot_r_state[2]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_tri/p_0_in0_in ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/FSM_onehot_r_state_reg[3] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[6]_i_1_n_0 ),
        .D(\FSM_onehot_r_state[3]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_tri/w_set_v1_y ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/FSM_onehot_r_state_reg[4] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[6]_i_1_n_0 ),
        .D(\FSM_onehot_r_state[4]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_tri/p_0_in ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/FSM_onehot_r_state_reg[5] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[6]_i_1_n_0 ),
        .D(\FSM_onehot_r_state[5]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_tri/w_set_v2_y ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/FSM_onehot_r_state_reg[6] 
       (.C(clk_i),
        .CE(\FSM_onehot_r_state[6]_i_1_n_0 ),
        .D(\FSM_onehot_r_state[6]_i_2_n_0 ),
        .Q(\u_geo/w_en_tri ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_outcode_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/w_outcode_view [0]),
        .Q(\u_geo/u_geo_tri/r_v0_outcode [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_outcode_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/w_outcode_view [1]),
        .Q(\u_geo/u_geo_tri/r_v0_outcode [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_outcode_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/w_outcode_view [2]),
        .Q(\u_geo/u_geo_tri/r_v0_outcode [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_outcode_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/w_outcode_view [3]),
        .Q(\u_geo/u_geo_tri/r_v0_outcode [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_outcode_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/w_outcode_view [4]),
        .Q(\u_geo/u_geo_tri/r_v0_outcode [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_outcode_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/w_outcode_view [5]),
        .Q(\u_geo/u_geo_tri/r_v0_outcode [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_x_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [0]),
        .Q(\u_geo/w_v0_x_tri [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_x_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [10]),
        .Q(\u_geo/w_v0_x_tri [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_x_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [11]),
        .Q(\u_geo/w_v0_x_tri [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_x_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [1]),
        .Q(\u_geo/w_v0_x_tri [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_x_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [2]),
        .Q(\u_geo/w_v0_x_tri [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_x_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [3]),
        .Q(\u_geo/w_v0_x_tri [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_x_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [4]),
        .Q(\u_geo/w_v0_x_tri [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_x_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [5]),
        .Q(\u_geo/w_v0_x_tri [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_x_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [6]),
        .Q(\u_geo/w_v0_x_tri [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_x_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [7]),
        .Q(\u_geo/w_v0_x_tri [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_x_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [8]),
        .Q(\u_geo/w_v0_x_tri [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_x_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [9]),
        .Q(\u_geo/w_v0_x_tri [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_y_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [0]),
        .Q(\u_geo/w_v0_y_tri [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_y_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [10]),
        .Q(\u_geo/w_v0_y_tri [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_y_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [11]),
        .Q(\u_geo/w_v0_y_tri [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_y_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [1]),
        .Q(\u_geo/w_v0_y_tri [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_y_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [2]),
        .Q(\u_geo/w_v0_y_tri [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_y_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [3]),
        .Q(\u_geo/w_v0_y_tri [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_y_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [4]),
        .Q(\u_geo/w_v0_y_tri [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_y_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [5]),
        .Q(\u_geo/w_v0_y_tri [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_y_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [6]),
        .Q(\u_geo/w_v0_y_tri [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_y_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [7]),
        .Q(\u_geo/w_v0_y_tri [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_y_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [8]),
        .Q(\u_geo/w_v0_y_tri [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v0_y_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v0_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [9]),
        .Q(\u_geo/w_v0_y_tri [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_outcode_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/w_outcode_view [0]),
        .Q(\u_geo/u_geo_tri/r_v1_outcode [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_outcode_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/w_outcode_view [1]),
        .Q(\u_geo/u_geo_tri/r_v1_outcode [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_outcode_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/w_outcode_view [2]),
        .Q(\u_geo/u_geo_tri/r_v1_outcode [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_outcode_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/w_outcode_view [3]),
        .Q(\u_geo/u_geo_tri/r_v1_outcode [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_outcode_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/w_outcode_view [4]),
        .Q(\u_geo/u_geo_tri/r_v1_outcode [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_outcode_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/w_outcode_view [5]),
        .Q(\u_geo/u_geo_tri/r_v1_outcode [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_x_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [0]),
        .Q(\u_geo/w_v1_x_tri [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_x_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [10]),
        .Q(\u_geo/w_v1_x_tri [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_x_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [11]),
        .Q(\u_geo/w_v1_x_tri [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_x_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [1]),
        .Q(\u_geo/w_v1_x_tri [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_x_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [2]),
        .Q(\u_geo/w_v1_x_tri [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_x_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [3]),
        .Q(\u_geo/w_v1_x_tri [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_x_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [4]),
        .Q(\u_geo/w_v1_x_tri [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_x_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [5]),
        .Q(\u_geo/w_v1_x_tri [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_x_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [6]),
        .Q(\u_geo/w_v1_x_tri [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_x_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [7]),
        .Q(\u_geo/w_v1_x_tri [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_x_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [8]),
        .Q(\u_geo/w_v1_x_tri [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_x_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [9]),
        .Q(\u_geo/w_v1_x_tri [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_y_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [0]),
        .Q(\u_geo/w_v1_y_tri [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_y_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [10]),
        .Q(\u_geo/w_v1_y_tri [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_y_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [11]),
        .Q(\u_geo/w_v1_y_tri [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_y_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [1]),
        .Q(\u_geo/w_v1_y_tri [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_y_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [2]),
        .Q(\u_geo/w_v1_y_tri [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_y_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [3]),
        .Q(\u_geo/w_v1_y_tri [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_y_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [4]),
        .Q(\u_geo/w_v1_y_tri [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_y_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [5]),
        .Q(\u_geo/w_v1_y_tri [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_y_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [6]),
        .Q(\u_geo/w_v1_y_tri [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_y_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [7]),
        .Q(\u_geo/w_v1_y_tri [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_y_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [8]),
        .Q(\u_geo/w_v1_y_tri [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v1_y_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v1_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [9]),
        .Q(\u_geo/w_v1_y_tri [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_outcode_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/w_outcode_view [0]),
        .Q(\u_geo/u_geo_tri/r_v2_outcode [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_outcode_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/w_outcode_view [1]),
        .Q(\u_geo/u_geo_tri/r_v2_outcode [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_outcode_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/w_outcode_view [2]),
        .Q(\u_geo/u_geo_tri/r_v2_outcode [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_outcode_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/w_outcode_view [3]),
        .Q(\u_geo/u_geo_tri/r_v2_outcode [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_outcode_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/w_outcode_view [4]),
        .Q(\u_geo/u_geo_tri/r_v2_outcode [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_outcode_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/w_outcode_view [5]),
        .Q(\u_geo/u_geo_tri/r_v2_outcode [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_x_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [0]),
        .Q(\u_geo/w_v2_x_tri [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_x_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [10]),
        .Q(\u_geo/w_v2_x_tri [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_x_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [11]),
        .Q(\u_geo/w_v2_x_tri [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_x_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [1]),
        .Q(\u_geo/w_v2_x_tri [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_x_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [2]),
        .Q(\u_geo/w_v2_x_tri [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_x_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [3]),
        .Q(\u_geo/w_v2_x_tri [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_x_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [4]),
        .Q(\u_geo/w_v2_x_tri [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_x_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [5]),
        .Q(\u_geo/w_v2_x_tri [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_x_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [6]),
        .Q(\u_geo/w_v2_x_tri [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_x_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [7]),
        .Q(\u_geo/w_v2_x_tri [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_x_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [8]),
        .Q(\u_geo/w_v2_x_tri [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_x_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_x ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [9]),
        .Q(\u_geo/w_v2_x_tri [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_y_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [0]),
        .Q(\u_geo/w_v2_y_tri [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_y_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [10]),
        .Q(\u_geo/w_v2_y_tri [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_y_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [11]),
        .Q(\u_geo/w_v2_y_tri [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_y_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [1]),
        .Q(\u_geo/w_v2_y_tri [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_y_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [2]),
        .Q(\u_geo/w_v2_y_tri [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_y_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [3]),
        .Q(\u_geo/w_v2_y_tri [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_y_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [4]),
        .Q(\u_geo/w_v2_y_tri [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_y_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [5]),
        .Q(\u_geo/w_v2_y_tri [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_y_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [6]),
        .Q(\u_geo/w_v2_y_tri [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_y_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [7]),
        .Q(\u_geo/w_v2_y_tri [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_y_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [8]),
        .Q(\u_geo/w_v2_y_tri [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_v2_y_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_v2_y ),
        .D(\u_geo/u_geo_tri/p_0_in__0 [9]),
        .Q(\u_geo/w_v2_y_tri [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [0]),
        .Q(\u_geo/u_geo_tri/r_vy [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [10]),
        .Q(\u_geo/u_geo_tri/r_vy [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [11]),
        .Q(\u_geo/u_geo_tri/r_vy [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[12] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [12]),
        .Q(\u_geo/u_geo_tri/r_vy [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[13] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [13]),
        .Q(\u_geo/u_geo_tri/r_vy [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[14] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [14]),
        .Q(\u_geo/u_geo_tri/r_vy [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[15] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [15]),
        .Q(\u_geo/u_geo_tri/r_vy [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[16] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [16]),
        .Q(\u_geo/u_geo_tri/r_vy [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[17] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [17]),
        .Q(\u_geo/u_geo_tri/r_vy [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[18] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [18]),
        .Q(\u_geo/u_geo_tri/r_vy [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[19] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [19]),
        .Q(\u_geo/u_geo_tri/r_vy [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [1]),
        .Q(\u_geo/u_geo_tri/r_vy [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[20] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [20]),
        .Q(\u_geo/u_geo_tri/r_vy [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[21] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [21]),
        .Q(\u_geo/u_geo_tri/r_vy [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [2]),
        .Q(\u_geo/u_geo_tri/r_vy [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [3]),
        .Q(\u_geo/u_geo_tri/r_vy [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [4]),
        .Q(\u_geo/u_geo_tri/r_vy [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [5]),
        .Q(\u_geo/u_geo_tri/r_vy [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [6]),
        .Q(\u_geo/u_geo_tri/r_vy [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [7]),
        .Q(\u_geo/u_geo_tri/r_vy [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [8]),
        .Q(\u_geo/u_geo_tri/r_vy [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_tri/r_vy_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_tri/w_set_y ),
        .D(\u_geo/w_vy_view [9]),
        .Q(\u_geo/u_geo_tri/r_vy [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/FSM_sequential_r_state_reg[0] 
       (.C(clk_i),
        .CE(FSM_sequential_r_state_reg),
        .D(FSM_sequential_r_state),
        .Q(\u_geo/u_geo_viewport/r_state [0]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/FSM_sequential_r_state_reg[1] 
       (.C(clk_i),
        .CE(FSM_sequential_r_state_reg),
        .D(\FSM_sequential_r_state[1]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_viewport/r_state [1]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/FSM_sequential_r_state_reg[2] 
       (.C(clk_i),
        .CE(FSM_sequential_r_state_reg),
        .D(\FSM_sequential_r_state[2]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_viewport/r_state [2]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/FSM_sequential_r_state_reg[3] 
       (.C(clk_i),
        .CE(FSM_sequential_r_state_reg),
        .D(\FSM_sequential_r_state[3]_i_2_n_0 ),
        .Q(\u_geo/u_geo_viewport/r_state [3]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_outcode_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/w_state_view ),
        .D(\u_geo/w_outcode_pdiv [0]),
        .Q(\u_geo/w_outcode_view [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_outcode_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/w_state_view ),
        .D(\u_geo/w_outcode_pdiv [1]),
        .Q(\u_geo/w_outcode_view [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_outcode_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/w_state_view ),
        .D(\u_geo/w_outcode_pdiv [2]),
        .Q(\u_geo/w_outcode_view [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_outcode_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/w_state_view ),
        .D(\u_geo/w_outcode_pdiv [3]),
        .Q(\u_geo/w_outcode_view [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_outcode_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/w_state_view ),
        .D(\u_geo/w_outcode_pdiv [4]),
        .Q(\u_geo/w_outcode_view [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_outcode_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/w_state_view ),
        .D(\u_geo/w_outcode_pdiv [5]),
        .Q(\u_geo/w_outcode_view [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[0] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_ ),
        .Q(\u_geo/w_vx_view [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[10] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[10] ),
        .Q(\u_geo/w_vx_view [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[11] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[11] ),
        .Q(\u_geo/w_vx_view [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[12] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[12] ),
        .Q(\u_geo/w_vx_view [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[13] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[13] ),
        .Q(\u_geo/w_vx_view [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[14] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[14] ),
        .Q(\u_geo/w_vx_view [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[15] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[15] ),
        .Q(\u_geo/w_vx_view [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[16] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[16] ),
        .Q(\u_geo/w_vx_view [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[17] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[17] ),
        .Q(\u_geo/w_vx_view [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[18] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[18] ),
        .Q(\u_geo/w_vx_view [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[19] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[19] ),
        .Q(\u_geo/w_vx_view [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[1] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[1] ),
        .Q(\u_geo/w_vx_view [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[20] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[20] ),
        .Q(\u_geo/w_vx_view [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[21] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[21] ),
        .Q(\u_geo/w_vx_view [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[2] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[2] ),
        .Q(\u_geo/w_vx_view [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[3] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[3] ),
        .Q(\u_geo/w_vx_view [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[4] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[4] ),
        .Q(\u_geo/w_vx_view [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[5] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[5] ),
        .Q(\u_geo/w_vx_view [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[6] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[6] ),
        .Q(\u_geo/w_vx_view [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[7] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[7] ),
        .Q(\u_geo/w_vx_view [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[8] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[8] ),
        .Q(\u_geo/w_vx_view [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vx_reg[9] 
       (.C(clk_i),
        .CE(\r_vx[21]_i_1__1_n_0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[9] ),
        .Q(\u_geo/w_vx_view [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[0] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_ ),
        .Q(\u_geo/w_vy_view [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[10] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[10] ),
        .Q(\u_geo/w_vy_view [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[11] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[11] ),
        .Q(\u_geo/w_vy_view [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[12] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[12] ),
        .Q(\u_geo/w_vy_view [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[13] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[13] ),
        .Q(\u_geo/w_vy_view [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[14] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[14] ),
        .Q(\u_geo/w_vy_view [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[15] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[15] ),
        .Q(\u_geo/w_vy_view [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[16] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[16] ),
        .Q(\u_geo/w_vy_view [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[17] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[17] ),
        .Q(\u_geo/w_vy_view [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[18] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[18] ),
        .Q(\u_geo/w_vy_view [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[19] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[19] ),
        .Q(\u_geo/w_vy_view [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[1] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[1] ),
        .Q(\u_geo/w_vy_view [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[20] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[20] ),
        .Q(\u_geo/w_vy_view [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[21] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[21] ),
        .Q(\u_geo/w_vy_view [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[2] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[2] ),
        .Q(\u_geo/w_vy_view [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[3] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[3] ),
        .Q(\u_geo/w_vy_view [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[4] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[4] ),
        .Q(\u_geo/w_vy_view [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[5] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[5] ),
        .Q(\u_geo/w_vy_view [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[6] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[6] ),
        .Q(\u_geo/w_vy_view [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[7] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[7] ),
        .Q(\u_geo/w_vy_view [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[8] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[8] ),
        .Q(\u_geo/w_vy_view [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/r_vy_reg[9] 
       (.C(clk_i),
        .CE(\u_geo/u_geo_viewport/w_set_vy ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[9] ),
        .Q(\u_geo/w_vy_view [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry_n_0 ,\u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry_n_1 ,\u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry_n_2 ,\u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry_n_3 }),
        .CYINIT(\u_geo/u_geo_viewport/r_exp_2z [0]),
        .DI({\u_geo/u_geo_viewport/r_exp_2z [3:1],_inferred__1_carry_i_1__18_n_0}),
        .O(\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [3:0]),
        .S({_inferred__1_carry_i_2__8_n_0,_inferred__1_carry_i_3__8_n_0,_inferred__1_carry_i_4__8_n_0,_inferred__1_carry_i_5__10_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry__0 
       (.CI(\u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_viewport/u_fadd/r_mats [16]}),
        .O({\u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry__0_n_4 ,\u_geo/u_geo_viewport/u_fadd/norm/_inferred__1_carry__0_n_5 ,\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [5:4]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,_inferred__1_carry_i_1__17_n_0,_inferred__1_carry_i_2__20_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_c_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fadd/norm/w_c_exp [0]),
        .Q(\u_geo/u_geo_viewport/w_a_exp [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_c_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fadd/norm/w_c_exp [1]),
        .Q(\u_geo/u_geo_viewport/w_a_exp [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_c_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fadd/norm/w_c_exp [2]),
        .Q(\u_geo/u_geo_viewport/w_a_exp [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_c_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fadd/norm/w_c_exp [3]),
        .Q(\u_geo/u_geo_viewport/w_a_exp [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_c_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fadd/norm/w_c_exp [4]),
        .Q(\u_geo/u_geo_viewport/w_a_exp [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fadd/w_c [21]),
        .Q(\u_geo/u_geo_viewport/w_fadd_out ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_exp_1z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fadd/w_exp_l [0]),
        .Q(\u_geo/u_geo_viewport/r_exp_1z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_exp_1z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fadd/w_exp_l [1]),
        .Q(\u_geo/u_geo_viewport/r_exp_1z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_exp_1z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fadd/w_exp_l [2]),
        .Q(\u_geo/u_geo_viewport/r_exp_1z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_exp_1z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fadd/w_exp_l [3]),
        .Q(\u_geo/u_geo_viewport/r_exp_1z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_exp_1z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [20]),
        .Q(\u_geo/u_geo_viewport/r_exp_1z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_exp_2z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/r_exp_1z [0]),
        .Q(\u_geo/u_geo_viewport/r_exp_2z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_exp_2z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/r_exp_1z [1]),
        .Q(\u_geo/u_geo_viewport/r_exp_2z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_exp_2z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/r_exp_1z [2]),
        .Q(\u_geo/u_geo_viewport/r_exp_2z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_exp_2z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/r_exp_1z [3]),
        .Q(\u_geo/u_geo_viewport/r_exp_2z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_exp_2z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/r_exp_1z [4]),
        .Q(\u_geo/u_geo_viewport/r_exp_2z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [0]),
        .Q(\u_geo/u_geo_viewport/r_f0 [0]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [10]),
        .Q(\u_geo/u_geo_viewport/r_f0 [10]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [11]),
        .Q(\u_geo/u_geo_viewport/r_f0 [11]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [12]),
        .Q(\u_geo/u_geo_viewport/r_f0 [12]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [13]),
        .Q(\u_geo/u_geo_viewport/r_f0 [13]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [14]),
        .Q(\u_geo/u_geo_viewport/r_f0 [14]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f0 ),
        .Q(\u_geo/u_geo_viewport/r_f0 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [1]),
        .Q(\u_geo/u_geo_viewport/r_f0 [1]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [2]),
        .Q(\u_geo/u_geo_viewport/r_f0 [2]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [3]),
        .Q(\u_geo/u_geo_viewport/r_f0 [3]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [4]),
        .Q(\u_geo/u_geo_viewport/r_f0 [4]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [5]),
        .Q(\u_geo/u_geo_viewport/r_f0 [5]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [6]),
        .Q(\u_geo/u_geo_viewport/r_f0 [6]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [7]),
        .Q(\u_geo/u_geo_viewport/r_f0 [7]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [8]),
        .Q(\u_geo/u_geo_viewport/r_f0 [8]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f0_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [9]),
        .Q(\u_geo/u_geo_viewport/r_f0 [9]),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [0]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [10]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [11]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [12]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [13]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [14]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [15]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [1]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [2]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [3]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [4]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [5]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [6]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [7]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [8]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_f1t_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_f1t [9]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_f1t_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [0]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [10]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [11]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [12]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [13]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [14]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [15]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [16]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [1]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [2]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [3]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [4]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [5]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [6]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [7]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [8]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_mats_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_mats [9]),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_mats [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_sign_1z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [21]),
        .Q(\u_geo/u_geo_viewport/r_sign_1z ),
        .R(\u_geo/u_geo_viewport/u_fadd/w_mag__7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_sign_2z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/r_sign_1z ),
        .Q(\u_geo/u_geo_viewport/u_fadd/r_sign_2z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fadd/r_sub_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_fadd_a [21]),
        .Q(\u_geo/u_geo_viewport/r_sub ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry_n_0 ,\u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry_n_1 ,\u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry_n_2 ,\u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry_n_3 }),
        .CYINIT(\u_geo/u_geo_viewport/r_ce_tmp_2z [0]),
        .DI({\u_geo/u_geo_viewport/r_ce_tmp_2z [3:1],_inferred__1_carry_i_1__20_n_0}),
        .O(\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [3:0]),
        .S({_inferred__1_carry_i_2__9_n_0,_inferred__1_carry_i_3__9_n_0,_inferred__1_carry_i_4__9_n_0,_inferred__1_carry_i_5__9_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry__0 
       (.CI(\u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]}),
        .O({\u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry__0_n_4 ,\u_geo/u_geo_viewport/u_fmul/norm/_inferred__1_carry__0_n_5 ,\u_geo/u_geo_viewport/u_fmul/norm/f_incdec_return [5:4]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,_inferred__1_carry_i_1__19_n_0,_inferred__1_carry_i_2__21_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[0]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_ ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[10]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[10] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[11]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[11] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[12]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[12] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[13]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[13] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[14]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[14] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/w_c ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/norm/w_c_exp [0]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/norm/w_c_exp [1]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/norm/w_c_exp [2]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/norm/w_c_exp [3]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[1]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[1] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/norm/w_c_exp [4]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_sign_2z ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[21] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[2]_i_1__1_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[2] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[3]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[3] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[4]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[4] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[5]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[5] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[6]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[6] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[7]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[7] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[8]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[8] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_c_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_c[9]_i_1__8_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_c_reg_n_0_[9] ),
        .R(\u_fmul/r_c ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_ce_tmp_1z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_fmul/r_ce_tmp_1z ),
        .Q(\u_geo/u_geo_viewport/r_ce_tmp_1z [0]),
        .R(\u_geo/u_geo_viewport/u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_ce_tmp_1z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_fmul/r_ce_tmp_1z[1]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_viewport/r_ce_tmp_1z [1]),
        .R(\u_geo/u_geo_viewport/u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_ce_tmp_1z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_fmul/r_ce_tmp_1z[2]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_viewport/r_ce_tmp_1z [2]),
        .R(\u_geo/u_geo_viewport/u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_ce_tmp_1z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_fmul/r_ce_tmp_1z[3]_i_1__0_n_0 ),
        .Q(\u_geo/u_geo_viewport/r_ce_tmp_1z [3]),
        .R(\u_geo/u_geo_viewport/u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_ce_tmp_1z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_fmul/r_ce_tmp_1z[4]_i_2__0_n_0 ),
        .Q(\u_geo/u_geo_viewport/r_ce_tmp_1z [4]),
        .R(\u_geo/u_geo_viewport/u_fmul/r_ce_tmp_1z ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_ce_tmp_2z_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/r_ce_tmp_1z [0]),
        .Q(\u_geo/u_geo_viewport/r_ce_tmp_2z [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_ce_tmp_2z_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/r_ce_tmp_1z [1]),
        .Q(\u_geo/u_geo_viewport/r_ce_tmp_2z [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_ce_tmp_2z_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/r_ce_tmp_1z [2]),
        .Q(\u_geo/u_geo_viewport/r_ce_tmp_2z [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_ce_tmp_2z_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/r_ce_tmp_1z [3]),
        .Q(\u_geo/u_geo_viewport/r_ce_tmp_2z [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_ce_tmp_2z_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/r_ce_tmp_1z [4]),
        .Q(\u_geo/u_geo_viewport/r_ce_tmp_2z [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2[3]_i_5 
       (.I0(\u_geo/u_geo_viewport/p_0_in [1]),
        .I1(\u_geo/u_geo_viewport/p_0_in [0]),
        .O(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [0]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [10]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [11]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[11]_i_1 
       (.CI(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[7]_i_1_n_0 ),
        .CO(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_viewport/w_cf_tmp2 [11:8]),
        .S(\u_geo/u_geo_viewport/p_0_in [12:9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [12]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [13]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [14]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [15]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[15]_i_1 
       (.CI(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg [3]),
        .CO({\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[15]_i_1_n_0 ,\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[15]_i_1_n_1 ,\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[15]_i_1_n_2 ,\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_viewport/w_cf_tmp2 [15:12]),
        .S(\u_geo/u_geo_viewport/p_0_in [16:13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [16]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[16]_i_1 
       (.CI(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[15]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[16]_i_1_n_4 ,\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[16]_i_1_n_5 ,\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[16]_i_1_n_6 ,\u_geo/u_geo_viewport/w_cf_tmp2 [16]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_viewport/p_0_in [17]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [1]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [2]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [3]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[3]_i_1_n_0 ,\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[3]_i_1_n_1 ,\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[3]_i_1_n_2 ,\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_viewport/p_0_in [1]}),
        .O(\u_geo/u_geo_viewport/w_cf_tmp2 [3:0]),
        .S({\u_geo/u_geo_viewport/p_0_in [4:2],\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2[3]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [4]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [5]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [6]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [7]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[7]_i_1 
       (.CI(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[3]_i_1_n_0 ),
        .CO({\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[7]_i_1_n_0 ,\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[7]_i_1_n_1 ,\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[7]_i_1_n_2 ,\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\u_geo/u_geo_viewport/w_cf_tmp2 [7:4]),
        .S(\u_geo/u_geo_viewport/p_0_in [8:5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [8]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_cf_tmp2_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/w_cf_tmp2 [9]),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_cf_tmp2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_sign_1z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/w_sign ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_sign_1z_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_geo/u_geo_viewport/u_fmul/r_sign_2z_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_geo/u_geo_viewport/u_fmul/r_sign_1z_reg_n_0 ),
        .Q(\u_geo/u_geo_viewport/u_fmul/r_sign_2z ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \u_geo/u_geo_viewport/u_fmul/w_cf_tmp 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_viewport/u_fadd/w_c [15:0]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\u_geo/u_geo_viewport/w_fmul_b }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const1>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const1>__0__0 ),
        .CLK(clk_i),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_58 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_59 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_60 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_61 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_62 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_63 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_64 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_65 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_66 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_67 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_68 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_69 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_70 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_71 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_72 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_73 ,\u_geo/u_geo_viewport/p_0_in ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_92 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_93 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_94 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_95 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_96 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_97 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_98 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_99 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_100 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_101 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_102 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_103 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_104 ,\u_geo/u_geo_viewport/u_fmul/w_cf_tmp_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_mem_arb/r_req_geo_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_req_geo_i_1_n_0),
        .Q(\u_mem_arb/r_req_geo ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_mem_arb/r_state_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_state_i_1__0_n_0),
        .Q(\u_mem_arb/r_state ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/_inferred__1_carry_n_0 ,\u_ras/u_ras_line/_inferred__1_carry_n_1 ,\u_ras/u_ras_line/_inferred__1_carry_n_2 ,\u_ras/u_ras_line/_inferred__1_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI(\u_ras/p_1_in [3:0]),
        .O(\u_ras/w_dy [3:0]),
        .S({_inferred__1_carry_i_5_n_0,_inferred__1_carry_i_6__10_n_0,_inferred__1_carry_i_7__10_n_0,_inferred__1_carry_i_8__10_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/_inferred__1_carry__0 
       (.CI(\u_ras/u_ras_line/_inferred__1_carry_n_0 ),
        .CO({\u_ras/u_ras_line/_inferred__1_carry__0_n_0 ,\u_ras/u_ras_line/_inferred__1_carry__0_n_1 ,\u_ras/u_ras_line/_inferred__1_carry__0_n_2 ,\u_ras/u_ras_line/_inferred__1_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_ras/p_1_in [7:4]),
        .O(\u_ras/w_dy [7:4]),
        .S({_inferred__1_carry__0_i_5_n_0,_inferred__1_carry__0_i_6_n_0,_inferred__1_carry__0_i_7_n_0,_inferred__1_carry__0_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/_inferred__1_carry__1 
       (.CI(\u_ras/u_ras_line/_inferred__1_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\u_ras/p_1_in [10:8]}),
        .O(\u_ras/w_dy [11:8]),
        .S({_inferred__1_carry__1_i_4_n_0,_inferred__1_carry__1_i_5_n_0,_inferred__1_carry__1_i_6_n_0,_inferred__1_carry__1_i_7_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/_inferred__5_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/_inferred__5_carry_n_0 ,\u_ras/u_ras_line/_inferred__5_carry_n_1 ,\u_ras/u_ras_line/_inferred__5_carry_n_2 ,\u_ras/u_ras_line/_inferred__5_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI(\u_ras/p_2_in [3:0]),
        .O({\u_ras/u_ras_line/_inferred__5_carry_n_4 ,\u_ras/u_ras_line/_inferred__5_carry_n_5 ,\u_ras/u_ras_line/_inferred__5_carry_n_6 ,\u_ras/u_ras_line/_inferred__5_carry_n_7 }),
        .S({_inferred__5_carry_i_5_n_0,_inferred__5_carry_i_6_n_0,_inferred__5_carry_i_7_n_0,_inferred__5_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/_inferred__5_carry__0 
       (.CI(\u_ras/u_ras_line/_inferred__5_carry_n_0 ),
        .CO({\u_ras/u_ras_line/_inferred__5_carry__0_n_0 ,\u_ras/u_ras_line/_inferred__5_carry__0_n_1 ,\u_ras/u_ras_line/_inferred__5_carry__0_n_2 ,\u_ras/u_ras_line/_inferred__5_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\u_ras/p_2_in[7]_repN ,\u_ras/p_2_in [6:4]}),
        .O({\u_ras/u_ras_line/_inferred__5_carry__0_n_4 ,\u_ras/u_ras_line/_inferred__5_carry__0_n_5 ,\u_ras/u_ras_line/_inferred__5_carry__0_n_6 ,\u_ras/u_ras_line/_inferred__5_carry__0_n_7 }),
        .S({_inferred__5_carry__0_i_5_n_0,_inferred__5_carry__0_i_6_n_0,_inferred__5_carry__0_i_7_n_0,_inferred__5_carry__0_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/_inferred__5_carry__1 
       (.CI(\u_ras/u_ras_line/_inferred__5_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\u_ras/p_2_in [10:8]}),
        .O({\u_ras/u_ras_line/w_dx ,\u_ras/u_ras_line/_inferred__5_carry__1_n_5 ,\u_ras/u_ras_line/_inferred__5_carry__1_n_6 ,\u_ras/u_ras_line/_inferred__5_carry__1_n_7 }),
        .S({_inferred__5_carry__1_i_4_n_0,_inferred__5_carry__1_i_5_n_0,_inferred__5_carry__1_i_6_n_0,_inferred__5_carry__1_i_7_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/_inferred__8__0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/_inferred__8__0_carry_n_0 ,\u_ras/u_ras_line/_inferred__8__0_carry_n_1 ,\u_ras/u_ras_line/_inferred__8__0_carry_n_2 ,\u_ras/u_ras_line/_inferred__8__0_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({_inferred__8__0_carry_i_1_n_0,_inferred__8__0_carry_i_2_n_0,_inferred__8__0_carry_i_3_n_0,\<const0>__0__0 }),
        .O(\u_ras/r_err [3:0]),
        .S({_inferred__8__0_carry_i_4_n_0,_inferred__8__0_carry_i_5_n_0,_inferred__8__0_carry_i_6_n_0,_inferred__8__0_carry_i_7_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/_inferred__8__0_carry__0 
       (.CI(\u_ras/u_ras_line/_inferred__8__0_carry_n_0 ),
        .CO({\u_ras/u_ras_line/_inferred__8__0_carry__0_n_0 ,\u_ras/u_ras_line/_inferred__8__0_carry__0_n_1 ,\u_ras/u_ras_line/_inferred__8__0_carry__0_n_2 ,\u_ras/u_ras_line/_inferred__8__0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({_inferred__8__0_carry__0_i_1_n_0,_inferred__8__0_carry__0_i_2_n_0,_inferred__8__0_carry__0_i_3_n_0,_inferred__8__0_carry__0_i_4_n_0}),
        .O(\u_ras/r_err [7:4]),
        .S({_inferred__8__0_carry__0_i_5_n_0,_inferred__8__0_carry__0_i_6_n_0,_inferred__8__0_carry__0_i_7_n_0,_inferred__8__0_carry__0_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/_inferred__8__0_carry__1 
       (.CI(\u_ras/u_ras_line/_inferred__8__0_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,_inferred__8__0_carry__1_i_1_n_0,_inferred__8__0_carry__1_i_2_n_0}),
        .O({\u_ras/u_ras_line/_inferred__8__0_carry__1_n_4 ,\u_ras/r_err [10:8]}),
        .S({\<const0>__0__0 ,_inferred__8__0_carry__1_i_3_n_0,_inferred__8__0_carry__1_i_4_n_0,_inferred__8__0_carry__1_i_5_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_e2_reg[10] 
       (.C(clk_i),
        .CE(r_e2),
        .D(\u_ras/w_e2 [10]),
        .Q(\u_ras/r_e2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_e2_reg[11] 
       (.C(clk_i),
        .CE(r_e2),
        .D(\u_ras/w_e2 [11]),
        .Q(\u_ras/u_ras_line/r_e2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_e2_reg[1] 
       (.C(clk_i),
        .CE(r_e2),
        .D(\u_ras/w_e2 [1]),
        .Q(\u_ras/r_e2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_e2_reg[2] 
       (.C(clk_i),
        .CE(r_e2),
        .D(\u_ras/w_e2 [2]),
        .Q(\u_ras/r_e2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_e2_reg[3] 
       (.C(clk_i),
        .CE(r_e2),
        .D(\u_ras/w_e2 [3]),
        .Q(\u_ras/r_e2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_e2_reg[4] 
       (.C(clk_i),
        .CE(r_e2),
        .D(\u_ras/w_e2 [4]),
        .Q(\u_ras/r_e2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_e2_reg[5] 
       (.C(clk_i),
        .CE(r_e2),
        .D(\u_ras/w_e2 [5]),
        .Q(\u_ras/r_e2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_e2_reg[6] 
       (.C(clk_i),
        .CE(r_e2),
        .D(\u_ras/w_e2 [6]),
        .Q(\u_ras/r_e2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_e2_reg[7] 
       (.C(clk_i),
        .CE(r_e2),
        .D(\u_ras/w_e2 [7]),
        .Q(\u_ras/r_e2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_e2_reg[8] 
       (.C(clk_i),
        .CE(r_e2),
        .D(\u_ras/w_e2 [8]),
        .Q(\u_ras/r_e2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_e2_reg[9] 
       (.C(clk_i),
        .CE(r_e2),
        .D(\u_ras/w_e2 [9]),
        .Q(\u_ras/r_e2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_err_reg[0] 
       (.C(clk_i),
        .CE(\r_err[10]_i_1_n_0 ),
        .D(r_err),
        .Q(\u_ras/w_e2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_err_reg[10] 
       (.C(clk_i),
        .CE(\r_err[10]_i_1_n_0 ),
        .D(\r_err[10]_i_2_n_0 ),
        .Q(\u_ras/w_e2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_err_reg[1] 
       (.C(clk_i),
        .CE(\r_err[10]_i_1_n_0 ),
        .D(\r_err[1]_i_1_n_0 ),
        .Q(\u_ras/w_e2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_err_reg[2] 
       (.C(clk_i),
        .CE(\r_err[10]_i_1_n_0 ),
        .D(\r_err[2]_i_1_n_0 ),
        .Q(\u_ras/w_e2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_err_reg[3] 
       (.C(clk_i),
        .CE(\r_err[10]_i_1_n_0 ),
        .D(\r_err[3]_i_1_n_0 ),
        .Q(\u_ras/w_e2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_err_reg[4] 
       (.C(clk_i),
        .CE(\r_err[10]_i_1_n_0 ),
        .D(\r_err[4]_i_1_n_0 ),
        .Q(\u_ras/w_e2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_err_reg[5] 
       (.C(clk_i),
        .CE(\r_err[10]_i_1_n_0 ),
        .D(\r_err[5]_i_1_n_0 ),
        .Q(\u_ras/w_e2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_err_reg[6] 
       (.C(clk_i),
        .CE(\r_err[10]_i_1_n_0 ),
        .D(\r_err[6]_i_1_n_0 ),
        .Q(\u_ras/w_e2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_err_reg[7] 
       (.C(clk_i),
        .CE(\r_err[10]_i_1_n_0 ),
        .D(\r_err[7]_i_1_n_0 ),
        .Q(\u_ras/w_e2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_err_reg[8] 
       (.C(clk_i),
        .CE(\r_err[10]_i_1_n_0 ),
        .D(\r_err[8]_i_1_n_0 ),
        .Q(\u_ras/w_e2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_err_reg[9] 
       (.C(clk_i),
        .CE(\r_err[10]_i_1_n_0 ),
        .D(\r_err[9]_i_1_n_0 ),
        .Q(\u_ras/w_e2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_state_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_ras_line/r_state ),
        .Q(\u_ras/u_ras_line/r_state_reg_n_0_ ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_state_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_ras_line/r_state[1]_i_1_n_0 ),
        .Q(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x0_reg[0] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_x [0]),
        .Q(\u_ras/u_ras_line/r_x0 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x0_reg[10] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_x [10]),
        .Q(\u_ras/u_ras_line/r_x0 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x0_reg[11] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_x [11]),
        .Q(\u_ras/u_ras_line/r_x0 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x0_reg[1] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_x [1]),
        .Q(\u_ras/u_ras_line/r_x0 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x0_reg[2] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_x [2]),
        .Q(\u_ras/u_ras_line/r_x0 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x0_reg[3] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_x [3]),
        .Q(\u_ras/u_ras_line/r_x0 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x0_reg[4] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_x [4]),
        .Q(\u_ras/u_ras_line/r_x0 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x0_reg[5] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_x [5]),
        .Q(\u_ras/u_ras_line/r_x0 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x0_reg[6] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_x [6]),
        .Q(\u_ras/u_ras_line/r_x0 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x0_reg[7] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_x [7]),
        .Q(\u_ras/u_ras_line/r_x0 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x0_reg[8] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_x [8]),
        .Q(\u_ras/u_ras_line/r_x0 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x0_reg[9] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_x [9]),
        .Q(\u_ras/u_ras_line/r_x0 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x1_reg[0] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_x [0]),
        .Q(\u_ras/u_ras_line/r_x1 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x1_reg[10] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_x [10]),
        .Q(\u_ras/u_ras_line/r_x1 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x1_reg[11] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_x [11]),
        .Q(\u_ras/u_ras_line/r_x1 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x1_reg[1] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_x [1]),
        .Q(\u_ras/u_ras_line/r_x1 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x1_reg[2] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_x [2]),
        .Q(\u_ras/u_ras_line/r_x1 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x1_reg[3] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_x [3]),
        .Q(\u_ras/u_ras_line/r_x1 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x1_reg[4] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_x [4]),
        .Q(\u_ras/u_ras_line/r_x1 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x1_reg[5] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_x [5]),
        .Q(\u_ras/u_ras_line/r_x1 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x1_reg[6] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_x [6]),
        .Q(\u_ras/u_ras_line/r_x1 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x1_reg[7] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_x [7]),
        .Q(\u_ras/u_ras_line/r_x1 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x1_reg[8] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_x [8]),
        .Q(\u_ras/u_ras_line/r_x1 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x1_reg[9] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_x [9]),
        .Q(\u_ras/u_ras_line/r_x1 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x_reg[0] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_x ),
        .D(r_x),
        .Q(\u_ras/u_ras_line/r_x_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x_reg[10] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_x ),
        .D(\r_x[10]_i_1_n_0 ),
        .Q(\u_ras/u_ras_line/r_x_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x_reg[11] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_x ),
        .D(\r_x[11]_i_2_n_0 ),
        .Q(\u_ras/w_x ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x_reg[1] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_x ),
        .D(\r_x[1]_i_1_n_0 ),
        .Q(\u_ras/u_ras_line/r_x_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x_reg[2] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_x ),
        .D(\r_x[2]_i_1_n_0 ),
        .Q(\u_ras/u_ras_line/r_x_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x_reg[3] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_x ),
        .D(\r_x[3]_i_1_n_0 ),
        .Q(\u_ras/u_ras_line/r_x_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x_reg[4] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_x ),
        .D(\r_x[4]_i_1_n_0 ),
        .Q(\u_ras/u_ras_line/r_x_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x_reg[5] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_x ),
        .D(\r_x[5]_i_1_n_0 ),
        .Q(\u_ras/u_ras_line/r_x_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x_reg[6] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_x ),
        .D(\r_x[6]_i_1_n_0 ),
        .Q(\u_ras/u_ras_line/r_x_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x_reg[7] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_x ),
        .D(\r_x[7]_i_1_n_0 ),
        .Q(\u_ras/u_ras_line/r_x_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x_reg[8] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_x ),
        .D(\r_x[8]_i_1_n_0 ),
        .Q(\u_ras/u_ras_line/r_x_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_x_reg[9] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_x ),
        .D(\r_x[9]_i_1_n_0 ),
        .Q(\u_ras/u_ras_line/r_x_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y0_reg[0] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_y [0]),
        .Q(\u_ras/u_ras_line/r_y0 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y0_reg[10] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_y [10]),
        .Q(\u_ras/u_ras_line/r_y0 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y0_reg[11] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_y [11]),
        .Q(\u_ras/u_ras_line/r_y0 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y0_reg[1] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_y [1]),
        .Q(\u_ras/u_ras_line/r_y0 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y0_reg[2] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_y [2]),
        .Q(\u_ras/u_ras_line/r_y0 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y0_reg[3] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_y [3]),
        .Q(\u_ras/u_ras_line/r_y0 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y0_reg[4] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_y [4]),
        .Q(\u_ras/u_ras_line/r_y0 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y0_reg[5] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_y [5]),
        .Q(\u_ras/u_ras_line/r_y0 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y0_reg[6] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_y [6]),
        .Q(\u_ras/u_ras_line/r_y0 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y0_reg[7] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_y [7]),
        .Q(\u_ras/u_ras_line/r_y0 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y0_reg[8] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_y [8]),
        .Q(\u_ras/u_ras_line/r_y0 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y0_reg[9] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v0_y [9]),
        .Q(\u_ras/u_ras_line/r_y0 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y1_reg[0] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_y [0]),
        .Q(\u_ras/u_ras_line/r_y1_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y1_reg[10] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_y [10]),
        .Q(\u_ras/u_ras_line/r_y1_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y1_reg[11] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_y [11]),
        .Q(\u_ras/u_ras_line/r_y1_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y1_reg[1] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_y [1]),
        .Q(\u_ras/u_ras_line/r_y1_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y1_reg[2] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_y [2]),
        .Q(\u_ras/u_ras_line/r_y1_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y1_reg[3] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_y [3]),
        .Q(\u_ras/u_ras_line/r_y1_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y1_reg[4] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_y [4]),
        .Q(\u_ras/u_ras_line/r_y1_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y1_reg[5] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_y [5]),
        .Q(\u_ras/u_ras_line/r_y1_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y1_reg[6] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_y [6]),
        .Q(\u_ras/u_ras_line/r_y1_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y1_reg[7] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_y [7]),
        .Q(\u_ras/u_ras_line/r_y1_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y1_reg[8] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_y [8]),
        .Q(\u_ras/u_ras_line/r_y1_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y1_reg[9] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y1 ),
        .D(\u_ras/w_v1_y [9]),
        .Q(\u_ras/u_ras_line/r_y1_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y_reg[0] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y ),
        .D(r_y),
        .Q(\u_ras/r_y [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y_reg[10] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y ),
        .D(\r_y[10]_i_1_n_0 ),
        .Q(\u_ras/r_y [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y_reg[11] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y ),
        .D(\r_y[11]_i_2_n_0 ),
        .Q(\u_ras/w_y ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y_reg[1] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y ),
        .D(\r_y[1]_i_1_n_0 ),
        .Q(\u_ras/r_y [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y_reg[2] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y ),
        .D(\r_y[2]_i_1_n_0 ),
        .Q(\u_ras/r_y [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y_reg[3] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y ),
        .D(\r_y[3]_i_1_n_0 ),
        .Q(\u_ras/r_y [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y_reg[4] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y ),
        .D(\r_y[4]_i_1_n_0 ),
        .Q(\u_ras/r_y [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y_reg[5] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y ),
        .D(\r_y[5]_i_1_n_0 ),
        .Q(\u_ras/r_y [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y_reg[6] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y ),
        .D(\r_y[6]_i_1_n_0 ),
        .Q(\u_ras/r_y [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y_reg[7] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y ),
        .D(\r_y[7]_i_1_n_0 ),
        .Q(\u_ras/r_y [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y_reg[8] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y ),
        .D(\r_y[8]_i_1_n_0 ),
        .Q(\u_ras/r_y [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_line/r_y_reg[9] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_line/r_y ),
        .D(\r_y[9]_i_1_n_0 ),
        .Q(\u_ras/r_y [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/result0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/result0_carry_n_0 ,\u_ras/u_ras_line/result0_carry_n_1 ,\u_ras/u_ras_line/result0_carry_n_2 ,\u_ras/u_ras_line/result0_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({result0_carry_i_1_n_0,result0_carry_i_2_n_0,result0_carry_i_3_n_0,result0_carry_i_4_n_0}),
        .S({result0_carry_i_5_n_0,result0_carry_i_6_n_0,result0_carry_i_7_n_0,result0_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/result0_carry__0 
       (.CI(\u_ras/u_ras_line/result0_carry_n_0 ),
        .CO({\u_ras/u_ras_line/result0_carry__0_n_0 ,\u_ras/u_ras_line/result0_carry__0_n_1 ,\u_ras/u_ras_line/result0_carry__0_n_2 ,\u_ras/u_ras_line/result0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,result0_carry__0_i_1_n_0,result0_carry__0_i_2_n_0}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,result0_carry__0_i_3_n_0,result0_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/result0_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/result0_inferred__1_carry_n_0 ,\u_ras/u_ras_line/result0_inferred__1_carry_n_1 ,\u_ras/u_ras_line/result0_inferred__1_carry_n_2 ,\u_ras/u_ras_line/result0_inferred__1_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({result0_inferred__1_carry_i_1_n_0,result0_inferred__1_carry_i_2_n_0,result0_inferred__1_carry_i_3_n_0,result0_inferred__1_carry_i_4_n_0}),
        .S({result0_inferred__1_carry_i_5_n_0,result0_inferred__1_carry_i_6_n_0,result0_inferred__1_carry_i_7_n_0,result0_inferred__1_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/result0_inferred__1_carry__0 
       (.CI(\u_ras/u_ras_line/result0_inferred__1_carry_n_0 ),
        .CO({\u_ras/u_ras_line/result0_inferred__1_carry__0_n_0 ,\u_ras/u_ras_line/result0_inferred__1_carry__0_n_1 ,\u_ras/u_ras_line/result0_inferred__1_carry__0_n_2 ,\u_ras/u_ras_line/result0_inferred__1_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,result0_inferred__1_carry__0_i_1_n_0,result0_inferred__1_carry__0_i_2_n_0}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,result0_inferred__1_carry__0_i_3_n_0,result0_inferred__1_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_dym_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/w_dym_carry_n_0 ,\u_ras/u_ras_line/w_dym_carry_n_1 ,\u_ras/u_ras_line/w_dym_carry_n_2 ,\u_ras/u_ras_line/w_dym_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\u_ras/u_ras_line/w_dym_carry_n_4 ,\u_ras/u_ras_line/w_dym_carry_n_5 ,\u_ras/u_ras_line/w_dym_carry_n_6 ,\u_ras/u_ras_line/w_dym_carry_n_7 }),
        .S({w_dym_carry_i_1_n_0,w_dym_carry_i_2_n_0,w_dym_carry_i_3_n_0,\u_ras/w_dy [0]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_dym_carry__0 
       (.CI(\u_ras/u_ras_line/w_dym_carry_n_0 ),
        .CO({\u_ras/u_ras_line/w_dym_carry__0_n_0 ,\u_ras/u_ras_line/w_dym_carry__0_n_1 ,\u_ras/u_ras_line/w_dym_carry__0_n_2 ,\u_ras/u_ras_line/w_dym_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_ras/u_ras_line/w_dym_carry__0_n_4 ,\u_ras/u_ras_line/w_dym_carry__0_n_5 ,\u_ras/u_ras_line/w_dym_carry__0_n_6 ,\u_ras/u_ras_line/w_dym_carry__0_n_7 }),
        .S({w_dym_carry__0_i_1_n_0,w_dym_carry__0_i_2_n_0,w_dym_carry__0_i_3_n_0,w_dym_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_dym_carry__1 
       (.CI(\u_ras/u_ras_line/w_dym_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\u_ras/u_ras_line/w_dym__22 ,\u_ras/u_ras_line/w_dym_carry__1_n_5 ,\u_ras/u_ras_line/w_dym_carry__1_n_6 ,\u_ras/u_ras_line/w_dym_carry__1_n_7 }),
        .S({w_dym_carry__1_i_1_n_0,w_dym_carry__1_i_2_n_0,w_dym_carry__1_i_3_n_0,w_dym_carry__1_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_end0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/w_end0__3 ,\u_ras/u_ras_line/w_end0_carry_n_1 ,\u_ras/u_ras_line/w_end0_carry_n_2 ,\u_ras/u_ras_line/w_end0_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({w_end0_carry_i_1_n_0,w_end0_carry_i_2_n_0,w_end0_carry_i_3_n_0,w_end0_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_end0_inferred__0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/w_end00_out ,\u_ras/u_ras_line/w_end0_inferred__0_carry_n_1 ,\u_ras/u_ras_line/w_end0_inferred__0_carry_n_2 ,\u_ras/u_ras_line/w_end0_inferred__0_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({w_end0_inferred__0_carry_i_1_n_0,w_end0_inferred__0_carry_i_2_n_0,w_end0_inferred__0_carry_i_3_n_0,w_end0_inferred__0_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_err__0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/w_err__0_carry_n_0 ,\u_ras/u_ras_line/w_err__0_carry_n_1 ,\u_ras/u_ras_line/w_err__0_carry_n_2 ,\u_ras/u_ras_line/w_err__0_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({w_err__0_carry_i_1_n_0,w_err__0_carry_i_2_n_0,w_err__0_carry_i_3_n_0,\<const1>__0__0 }),
        .O(\u_ras/w_err [3:0]),
        .S({w_err__0_carry_i_4_n_0,w_err__0_carry_i_5_n_0,w_err__0_carry_i_6_n_0,w_err__0_carry_i_7_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_err__0_carry__0 
       (.CI(\u_ras/u_ras_line/w_err__0_carry_n_0 ),
        .CO({\u_ras/u_ras_line/w_err__0_carry__0_n_0 ,\u_ras/u_ras_line/w_err__0_carry__0_n_1 ,\u_ras/u_ras_line/w_err__0_carry__0_n_2 ,\u_ras/u_ras_line/w_err__0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({w_err__0_carry__0_i_1_n_0,w_err__0_carry__0_i_2_n_0,w_err__0_carry__0_i_3_n_0,w_err__0_carry__0_i_4_n_0}),
        .O(\u_ras/w_err [7:4]),
        .S({w_err__0_carry__0_i_5_n_0,w_err__0_carry__0_i_6_n_0,w_err__0_carry__0_i_7_n_0,w_err__0_carry__0_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_err__0_carry__1 
       (.CI(\u_ras/u_ras_line/w_err__0_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,w_err__0_carry__1_i_1_n_0,w_err__0_carry__1_i_2_n_0}),
        .O({\u_ras/u_ras_line/w_err__0_carry__1_n_4 ,\u_ras/w_err [10:8]}),
        .S({\<const0>__0__0 ,w_err__0_carry__1_i_3_n_0,w_err__0_carry__1_i_4_n_0,w_err__0_carry__1_i_5_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_reject0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/w_reject0_carry_n_0 ,\u_ras/u_ras_line/w_reject0_carry_n_1 ,\u_ras/u_ras_line/w_reject0_carry_n_2 ,\u_ras/u_ras_line/w_reject0_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({w_reject0_carry_i_1_n_0,w_reject0_carry_i_2_n_0,w_reject0_carry_i_3_n_0,w_reject0_carry_i_4_n_0}),
        .S({w_reject0_carry_i_5_n_0,w_reject0_carry_i_6_n_0,w_reject0_carry_i_7_n_0,w_reject0_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_reject0_carry__0 
       (.CI(\u_ras/u_ras_line/w_reject0_carry_n_0 ),
        .CO({\u_ras/u_ras_line/w_reject0__7 ,\u_ras/u_ras_line/w_reject0_carry__0_n_1 ,\u_ras/u_ras_line/w_reject0_carry__0_n_2 ,\u_ras/u_ras_line/w_reject0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,w_reject0_carry__0_i_1_n_0,w_reject0_carry__0_i_2_n_0}),
        .S({w_reject0_carry__0_i_3_n_0,w_reject0_carry__0_i_4_n_0,w_reject0_carry__0_i_5_n_0,w_reject0_carry__0_i_6_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_reject1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/w_reject1_carry_n_0 ,\u_ras/u_ras_line/w_reject1_carry_n_1 ,\u_ras/u_ras_line/w_reject1_carry_n_2 ,\u_ras/u_ras_line/w_reject1_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({w_reject1_carry_i_1_n_0,w_reject1_carry_i_2_n_0,w_reject1_carry_i_3_n_0,w_reject1_carry_i_4_n_0}),
        .S({w_reject1_carry_i_5_n_0,w_reject1_carry_i_6_n_0,w_reject1_carry_i_7_n_0,w_reject1_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_reject1_carry__0 
       (.CI(\u_ras/u_ras_line/w_reject1_carry_n_0 ),
        .CO({\u_ras/u_ras_line/w_reject1__7 ,\u_ras/u_ras_line/w_reject1_carry__0_n_1 ,\u_ras/u_ras_line/w_reject1_carry__0_n_2 ,\u_ras/u_ras_line/w_reject1_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,w_reject1_carry__0_i_1_n_0,w_reject1_carry__0_i_2_n_0}),
        .S({w_reject1_carry__0_i_3_n_0,w_reject1_carry__0_i_4_n_0,w_reject1_carry__0_i_5_n_0,w_reject1_carry__0_i_6_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_sx_flag1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/w_sx_flag1_carry_n_0 ,\u_ras/u_ras_line/w_sx_flag1_carry_n_1 ,\u_ras/u_ras_line/w_sx_flag1_carry_n_2 ,\u_ras/u_ras_line/w_sx_flag1_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({w_sx_flag1_carry_i_1_n_0,w_sx_flag1_carry_i_2_n_0,w_sx_flag1_carry_i_3_n_0,w_sx_flag1_carry_i_4_n_0}),
        .S({w_sx_flag1_carry_i_5_n_0,w_sx_flag1_carry_i_6_n_0,w_sx_flag1_carry_i_7_n_0,w_sx_flag1_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_line/w_sx_flag1_carry__0 
       (.CI(\u_ras/u_ras_line/w_sx_flag1_carry_n_0 ),
        .CO({\u_ras/u_ras_line/w_sx_flag1_carry__0_n_0 ,\u_ras/u_ras_line/w_sx_flag1_carry__0_n_1 ,\u_ras/u_ras_line/w_sx_flag1__5 ,\u_ras/u_ras_line/w_sx_flag1_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,w_sx_flag1_carry__0_i_1_n_0,w_sx_flag1_carry__0_i_2_n_0}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,w_sx_flag1_carry__0_i_3_n_0,w_sx_flag1_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_line/w_sy_flag1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_line/w_sy_flag1_carry_n_0 ,\u_ras/u_ras_line/w_sy_flag1_carry_n_1 ,\u_ras/u_ras_line/w_sy_flag1_carry_n_2 ,\u_ras/u_ras_line/w_sy_flag1_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({w_sy_flag1_carry_i_1_n_0,w_sy_flag1_carry_i_2_n_0,w_sy_flag1_carry_i_3_n_0,w_sy_flag1_carry_i_4_n_0}),
        .S({w_sy_flag1_carry_i_5_n_0,w_sy_flag1_carry_i_6_n_0,w_sy_flag1_carry_i_7_n_0,w_sy_flag1_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_line/w_sy_flag1_carry__0 
       (.CI(\u_ras/u_ras_line/w_sy_flag1_carry_n_0 ),
        .CO({\u_ras/u_ras_line/w_sy_flag1_carry__0_n_0 ,\u_ras/u_ras_line/w_sy_flag1_carry__0_n_1 ,\u_ras/u_ras_line/w_sy_flag1__5 ,\u_ras/u_ras_line/w_sy_flag1_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,w_sy_flag1_carry__0_i_1_n_0,w_sy_flag1_carry__0_i_2_n_0}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,w_sy_flag1_carry__0_i_3_n_0,w_sy_flag1_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_2 
       (.I0(w_pixel_top_address[11]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_94 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_3 
       (.I0(w_pixel_top_address[10]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_95 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_4 
       (.I0(w_pixel_top_address[9]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_96 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_5 
       (.I0(w_pixel_top_address[8]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_97 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[13]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_2 
       (.I0(w_pixel_top_address[15]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_90 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_3 
       (.I0(w_pixel_top_address[14]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_91 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_4 
       (.I0(w_pixel_top_address[13]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_92 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_5 
       (.I0(w_pixel_top_address[12]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_93 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[17]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_2 
       (.I0(w_pixel_top_address[19]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_86 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_3 
       (.I0(w_pixel_top_address[18]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_87 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_4 
       (.I0(w_pixel_top_address[17]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_88 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_5 
       (.I0(w_pixel_top_address[16]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_89 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[21]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[25]_INST_0_i_3 
       (.I0(w_pixel_top_address[22]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_83 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[25]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[25]_INST_0_i_4 
       (.I0(w_pixel_top_address[21]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_84 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[25]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[25]_INST_0_i_5 
       (.I0(w_pixel_top_address[20]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_85 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[25]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_2 
       (.I0(w_pixel_top_address[3]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_102 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_3 
       (.I0(w_pixel_top_address[2]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_103 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_4 
       (.I0(w_pixel_top_address[1]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_104 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_5 
       (.I0(w_pixel_top_address[0]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_105 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[5]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_2 
       (.I0(w_pixel_top_address[7]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_98 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_3 
       (.I0(w_pixel_top_address[6]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_99 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_4 
       (.I0(w_pixel_top_address[5]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_100 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_5 
       (.I0(w_pixel_top_address[4]),
        .I1(\u_ras/u_ras_mem/r_adrs_m_reg_n_101 ),
        .O(\u_ras/u_ras_mem/m_wb_adr_o[9]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \u_ras/u_ras_mem/m_wb_sel_o[0]_INST_0 
       (.I0(\u_ras/u_ras_mem/r_x [0]),
        .I1(\u_ras/u_ras_mem/r_x [1]),
        .O(m_wb_sel_o[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \u_ras/u_ras_mem/m_wb_sel_o[3]_INST_0 
       (.I0(\u_ras/u_ras_mem/r_x [0]),
        .I1(\u_ras/u_ras_mem/r_x [1]),
        .O(m_wb_sel_o[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \u_ras/u_ras_mem/r_adrs_m_reg 
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,w_scr_w[15:2]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\u_ras/B }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\r_x[11]_i_2_n_0 ,\r_x[10]_i_1_n_0 ,\r_x[9]_i_1_n_0 ,\r_x[8]_i_1_n_0 ,\r_x[7]_i_1_n_0 ,\r_x[6]_i_1_n_0 ,\r_x[5]_i_1_n_0 ,\r_x[4]_i_1_n_0 ,\r_x[3]_i_1_n_0 ,\r_x[2]_i_1_n_0 }),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\u_ras/u_ras_line/r_x ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(r_adrs_m_reg_i_1_n_0),
        .CLK(clk_i),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\u_ras/u_ras_mem/r_adrs_m_reg_n_58 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_59 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_60 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_61 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_62 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_63 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_64 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_65 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_66 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_67 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_68 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_69 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_70 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_71 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_72 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_73 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_74 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_75 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_76 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_77 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_78 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_79 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_80 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_81 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_82 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_83 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_84 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_85 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_86 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_87 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_88 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_89 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_90 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_91 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_92 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_93 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_94 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_95 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_96 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_97 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_98 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_99 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_100 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_101 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_102 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_103 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_104 ,\u_ras/u_ras_mem/r_adrs_m_reg_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_mem/r_state_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_state_i_1_n_0),
        .Q(\u_ras/u_ras_mem/r_state ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_mem/r_x_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_ras_mem/r_x ),
        .Q(\u_ras/u_ras_mem/r_x [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_mem/r_x_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\u_ras_mem/r_x[1]_i_1_n_0 ),
        .Q(\u_ras/u_ras_mem/r_x [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_mem/w_y0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_mem/w_y0_carry_n_0 ,\u_ras/u_ras_mem/w_y0_carry_n_1 ,\u_ras/u_ras_mem/w_y0_carry_n_2 ,\u_ras/u_ras_mem/w_y0_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI(w_scr_h_m1[3:0]),
        .O({\u_ras/u_ras_mem/w_y0_carry_n_4 ,\u_ras/u_ras_mem/w_y0_carry_n_5 ,\u_ras/u_ras_mem/w_y0_carry_n_6 ,\u_ras/u_ras_mem/w_y0_carry_n_7 }),
        .S({w_y0_carry_i_1__1_n_0,w_y0_carry_i_2__1_n_0,w_y0_carry_i_3__1_n_0,w_y0_carry_i_4__1_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_mem/w_y0_carry__0 
       (.CI(\u_ras/u_ras_mem/w_y0_carry_n_0 ),
        .CO({\u_ras/u_ras_mem/w_y0_carry__0_n_0 ,\u_ras/u_ras_mem/w_y0_carry__0_n_1 ,\u_ras/u_ras_mem/w_y0_carry__0_n_2 ,\u_ras/u_ras_mem/w_y0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(w_scr_h_m1[7:4]),
        .O({\u_ras/u_ras_mem/w_y0_carry__0_n_4 ,\u_ras/u_ras_mem/w_y0_carry__0_n_5 ,\u_ras/u_ras_mem/w_y0_carry__0_n_6 ,\u_ras/u_ras_mem/w_y0_carry__0_n_7 }),
        .S({w_y0_carry_i_1__0_n_0,w_y0_carry_i_2__0_n_0,w_y0_carry_i_3__0_n_0,w_y0_carry_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras/u_ras_mem/w_y0_carry__1 
       (.CI(\u_ras/u_ras_mem/w_y0_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,w_scr_h_m1[10:8]}),
        .O({\u_ras/u_ras_mem/w_y0_carry__1_n_4 ,\u_ras/u_ras_mem/w_y0_carry__1_n_5 ,\u_ras/u_ras_mem/w_y0_carry__1_n_6 ,\u_ras/u_ras_mem/w_y0_carry__1_n_7 }),
        .S({w_y0_carry_i_1_n_0,w_y0_carry_i_2_n_0,w_y0_carry_i_3_n_0,w_y0_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \u_ras/u_ras_state/ 
       (.I0(\u_ras/u_ras_state/r_state [0]),
        .I1(\u_ras/u_ras_state/r_state [1]),
        .O(w_ack));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFFFFFB8FF0000)) 
    \u_ras/u_ras_state/FSM_sequential_r_state[1]_i_2 
       (.I0(\u_ras/u_ras_state/f_reject1_return ),
        .I1(\u_ras/u_ras_state/r_state [1]),
        .I2(\u_ras/u_ras_state/f_reject_return ),
        .I3(w_sy_flag1_carry_i_10_n_0),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .I5(\u_ras/u_ras_state/FSM_sequential_r_state[1]_i_5_n_0 ),
        .O(\u_ras/u_ras_state/FSM_sequential_r_state ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBFB0)) 
    \u_ras/u_ras_state/FSM_sequential_r_state[1]_i_5 
       (.I0(\u_ras/u_ras_state/f_reject0_return ),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(\u_ras/u_ras_state/r_state [1]),
        .I3(w_en),
        .O(\u_ras/u_ras_state/FSM_sequential_r_state[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/FSM_sequential_r_state_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[0]_i_1__1_n_0 ),
        .Q(\u_ras/u_ras_state/r_state [0]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/FSM_sequential_r_state_reg[0]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/FSM_sequential_r_state_reg[0]_replica 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[0]_i_1__1_n_0 ),
        .Q(\u_ras/u_ras_state/r_state[0]_repN ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/FSM_sequential_r_state_reg[0]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/FSM_sequential_r_state_reg[0]_replica_1 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[0]_i_1__1_n_0 ),
        .Q(\u_ras/u_ras_state/r_state[0]_repN_1 ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/FSM_sequential_r_state_reg[0]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/FSM_sequential_r_state_reg[0]_replica_2 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[0]_i_1__1_n_0 ),
        .Q(\u_ras/u_ras_state/r_state[0]_repN_2 ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/FSM_sequential_r_state_reg[0]_replica" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/FSM_sequential_r_state_reg[0]_replica_3 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[0]_i_1__1_n_0 ),
        .Q(\u_ras/u_ras_state/r_state[0]_repN_3 ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/FSM_sequential_r_state_reg[0]_replica" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/FSM_sequential_r_state_reg[0]_replica_4 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[0]_i_1__1_n_0 ),
        .Q(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/FSM_sequential_r_state_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[1]_i_1__0_n_0 ),
        .Q(\u_ras/u_ras_state/r_state [1]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/FSM_sequential_r_state_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/FSM_sequential_r_state_reg[1]_replica 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[1]_i_1__0_n_0 ),
        .Q(\u_ras/u_ras_state/r_state[1]_repN ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/FSM_sequential_r_state_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/FSM_sequential_r_state_reg[1]_replica_1 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[1]_i_1__0_n_0 ),
        .Q(\u_ras/u_ras_state/r_state[1]_repN_1 ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/FSM_sequential_r_state_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/FSM_sequential_r_state_reg[1]_replica_2 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[1]_i_1__0_n_0 ),
        .Q(\u_ras/u_ras_state/r_state[1]_repN_2 ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/FSM_sequential_r_state_reg[1]_replica" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/FSM_sequential_r_state_reg[1]_replica_3 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\FSM_sequential_r_state[1]_i_1__0_n_0 ),
        .Q(\u_ras/u_ras_state/r_state[1]_repN_3 ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[0] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[0]),
        .Q(\u_ras/u_ras_state/r_v0_x_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[10] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[10]),
        .Q(\u_ras/u_ras_state/r_v0_x_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_v0_x_reg[10]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[10]_replica 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[10]),
        .Q(\u_ras/u_ras_state/r_v0_x_reg_n_0_[10]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[11] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[11]),
        .Q(\u_ras/u_ras_state/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[1] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[1]),
        .Q(\u_ras/u_ras_state/r_v0_x_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[2] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[2]),
        .Q(\u_ras/u_ras_state/r_v0_x_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[3] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[3]),
        .Q(\u_ras/u_ras_state/r_v0_x_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[4] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[4]),
        .Q(\u_ras/u_ras_state/r_v0_x_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[5] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[5]),
        .Q(\u_ras/u_ras_state/r_v0_x_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[6] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[6]),
        .Q(\u_ras/u_ras_state/r_v0_x_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[7] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[7]),
        .Q(\u_ras/u_ras_state/r_v0_x_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[8] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[8]),
        .Q(\u_ras/u_ras_state/r_v0_x_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_x_reg[9] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_x[9]),
        .Q(\u_ras/u_ras_state/r_v0_x_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[0] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[0]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[10] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[10]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_v0_y_reg[10]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[10]_replica 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[10]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_[10]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[11] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[11]),
        .Q(\u_ras/u_ras_state/p_0_in0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[1] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[1]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_v0_y_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[1]_replica 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[1]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_[1]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[2] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[2]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[3] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[3]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[4] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[4]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[5] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[5]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[6] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[6]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[7] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[7]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[8] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[8]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v0_y_reg[9] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v0_y[9]),
        .Q(\u_ras/u_ras_state/r_v0_y_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[0] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[0]),
        .Q(\u_ras/u_ras_state/r_v1_x_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[10] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[10]),
        .Q(\u_ras/u_ras_state/r_v1_x_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_v1_x_reg[10]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[10]_replica 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[10]),
        .Q(\u_ras/u_ras_state/r_v1_x_reg_n_0_[10]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[11] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[11]),
        .Q(\u_ras/u_ras_state/p_1_in8_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[1] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[1]),
        .Q(\u_ras/u_ras_state/r_v1_x_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[2] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[2]),
        .Q(\u_ras/u_ras_state/r_v1_x_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[3] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[3]),
        .Q(\u_ras/u_ras_state/r_v1_x_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[4] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[4]),
        .Q(\u_ras/u_ras_state/r_v1_x_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[5] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[5]),
        .Q(\u_ras/u_ras_state/r_v1_x_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[6] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[6]),
        .Q(\u_ras/u_ras_state/r_v1_x_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[7] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[7]),
        .Q(\u_ras/u_ras_state/r_v1_x_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[8] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[8]),
        .Q(\u_ras/u_ras_state/r_v1_x_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_x_reg[9] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_x[9]),
        .Q(\u_ras/u_ras_state/r_v1_x_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[0] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[0]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_v1_y_reg[0]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[0]_replica 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[0]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[0]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[10] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[10]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[11] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[11]),
        .Q(\u_ras/u_ras_state/p_1_in10_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[1] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[1]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_v1_y_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[1]_replica 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[1]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[1]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[2] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[2]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[3] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[3]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[4] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[4]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[5] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[5]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_v1_y_reg[5]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[5]_replica 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[5]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[5]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[6] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[6]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_v1_y_reg[6]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[6]_replica 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[6]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[6]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[7] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[7]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_v1_y_reg[7]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[7]_replica 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[7]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[7]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[8] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[8]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_v1_y_reg[8]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[8]_replica 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[8]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[8]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v1_y_reg[9] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v1_y[9]),
        .Q(\u_ras/u_ras_state/r_v1_y_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_x_reg[0] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_x[0]),
        .Q(\u_ras/u_ras_state/r_v2_x_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_x_reg[10] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_x[10]),
        .Q(\u_ras/u_ras_state/r_v2_x_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_x_reg[11] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_x[11]),
        .Q(\u_ras/u_ras_state/p_1_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_x_reg[1] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_x[1]),
        .Q(\u_ras/u_ras_state/r_v2_x_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_x_reg[2] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_x[2]),
        .Q(\u_ras/u_ras_state/r_v2_x_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_x_reg[3] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_x[3]),
        .Q(\u_ras/u_ras_state/r_v2_x_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_x_reg[4] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_x[4]),
        .Q(\u_ras/u_ras_state/r_v2_x_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_x_reg[5] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_x[5]),
        .Q(\u_ras/u_ras_state/r_v2_x_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_x_reg[6] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_x[6]),
        .Q(\u_ras/u_ras_state/r_v2_x_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_x_reg[7] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_x[7]),
        .Q(\u_ras/u_ras_state/r_v2_x_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_x_reg[8] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_x[8]),
        .Q(\u_ras/u_ras_state/r_v2_x_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_x_reg[9] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_x[9]),
        .Q(\u_ras/u_ras_state/r_v2_x_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[0] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[0]),
        .Q(\u_ras/u_ras_state/r_v2_y_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[10] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[10]),
        .Q(\u_ras/u_ras_state/r_v2_y_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[11] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[11]),
        .Q(\u_ras/u_ras_state/p_1_in1_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[1] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[1]),
        .Q(\u_ras/u_ras_state/r_v2_y_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[2] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[2]),
        .Q(\u_ras/u_ras_state/r_v2_y_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[3] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[3]),
        .Q(\u_ras/u_ras_state/r_v2_y_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[4] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[4]),
        .Q(\u_ras/u_ras_state/r_v2_y_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[5] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[5]),
        .Q(\u_ras/u_ras_state/r_v2_y_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[6] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[6]),
        .Q(\u_ras/u_ras_state/r_v2_y_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_v2_y_reg[6]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[6]_replica 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[6]),
        .Q(\u_ras/u_ras_state/r_v2_y_reg_n_0_[6]_repN ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[7] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[7]),
        .Q(\u_ras/u_ras_state/r_v2_y_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[8] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[8]),
        .Q(\u_ras/u_ras_state/r_v2_y_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_ras/u_ras_state/r_v2_y_reg[9] 
       (.C(clk_i),
        .CE(\u_ras/u_ras_state/w_set_vtx ),
        .D(w_v2_y[9]),
        .Q(\u_ras/u_ras_state/r_v2_y_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[0]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_ ),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_ ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_1 ),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_ ),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .O(\u_ras/w_v0_x [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[10]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[10] ),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_[10]_repN ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[10] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v0_x [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_x0[10]_i_1" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[10]_i_1_replica 
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[10]_repN ),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_[10]_repN ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[10] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v0_x[10]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[11]_i_1 
       (.I0(\u_ras/u_ras_state/p_0_in ),
        .I1(\u_ras/u_ras_state/p_1_in8_in ),
        .I2(\u_ras/u_ras_state/r_state [1]),
        .I3(\u_ras/u_ras_state/p_1_in ),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .O(\u_ras/w_v0_x [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[1]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[1] ),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_[1] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_1 ),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[1] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_1 ),
        .O(\u_ras/w_v0_x [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[2]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[2] ),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_[2] ),
        .I2(\u_ras/u_ras_state/r_state [1]),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[2] ),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .O(\u_ras/w_v0_x [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[3]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[3] ),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_[3] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_1 ),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[3] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_1 ),
        .O(\u_ras/w_v0_x [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[4]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[4] ),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_[4] ),
        .I2(\u_ras/u_ras_state/r_state [1]),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[4] ),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .O(\u_ras/w_v0_x [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[5]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[5] ),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_[5] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[5] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v0_x [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[6]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[6] ),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_[6] ),
        .I2(\u_ras/u_ras_state/r_state [1]),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[6] ),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .O(\u_ras/w_v0_x [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[7]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[7] ),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_[7] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_1 ),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[7] ),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .O(\u_ras/w_v0_x [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[8]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[8] ),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_[8] ),
        .I2(\u_ras/u_ras_state/r_state [1]),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[8] ),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .O(\u_ras/w_v0_x [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x0[9]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_x_reg_n_0_[9] ),
        .I1(\u_ras/u_ras_state/r_v1_x_reg_n_0_[9] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_2 ),
        .I3(\u_ras/u_ras_state/r_v2_x_reg_n_0_[9] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_1 ),
        .O(\u_ras/w_v0_x [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x1[0]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_ ),
        .I1(\u_ras/u_ras_state/r_v2_x_reg_n_0_ ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_1 ),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_ ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_1 ),
        .O(\u_ras/w_v1_x [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x1[10]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[10] ),
        .I1(\u_ras/u_ras_state/r_v2_x_reg_n_0_[10] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_2 ),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[10] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_1 ),
        .O(\u_ras/w_v1_x [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x1[11]_i_1 
       (.I0(\u_ras/u_ras_state/p_1_in8_in ),
        .I1(\u_ras/u_ras_state/p_1_in ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_1 ),
        .I3(\u_ras/u_ras_state/p_0_in ),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .O(\u_ras/w_v1_x [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x1[1]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[1] ),
        .I1(\u_ras/u_ras_state/r_v2_x_reg_n_0_[1] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_1 ),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[1] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_1 ),
        .O(\u_ras/w_v1_x [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x1[2]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[2] ),
        .I1(\u_ras/u_ras_state/r_v2_x_reg_n_0_[2] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_1 ),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[2] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_1 ),
        .O(\u_ras/w_v1_x [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x1[3]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[3] ),
        .I1(\u_ras/u_ras_state/r_v2_x_reg_n_0_[3] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_1 ),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[3] ),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .O(\u_ras/w_v1_x [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x1[4]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[4] ),
        .I1(\u_ras/u_ras_state/r_v2_x_reg_n_0_[4] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[4] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v1_x [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x1[5]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[5] ),
        .I1(\u_ras/u_ras_state/r_v2_x_reg_n_0_[5] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[5] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN ),
        .O(\u_ras/w_v1_x [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x1[6]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[6] ),
        .I1(\u_ras/u_ras_state/r_v2_x_reg_n_0_[6] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[6] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v1_x [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x1[7]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[7] ),
        .I1(\u_ras/u_ras_state/r_v2_x_reg_n_0_[7] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_1 ),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[7] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_1 ),
        .O(\u_ras/w_v1_x [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x1[8]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[8] ),
        .I1(\u_ras/u_ras_state/r_v2_x_reg_n_0_[8] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_1 ),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[8] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_1 ),
        .O(\u_ras/w_v1_x [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_x1[9]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_x_reg_n_0_[9] ),
        .I1(\u_ras/u_ras_state/r_v2_x_reg_n_0_[9] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_2 ),
        .I3(\u_ras/u_ras_state/r_v0_x_reg_n_0_[9] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_1 ),
        .O(\u_ras/w_v1_x [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[0]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_ ),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[0]_repN ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_3 ),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_ ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_3 ),
        .O(\u_ras/w_v0_y [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[10]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[10]_repN ),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[10] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[10] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN ),
        .O(\u_ras/w_v0_y [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "u_ras/u_ras_state/r_y0[10]_i_1" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[10]_i_1_replica 
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[10]_repN ),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[10] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_3 ),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[10] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_3 ),
        .O(\u_ras/w_v0_y[10]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[11]_i_1 
       (.I0(\u_ras/u_ras_state/p_0_in0_in ),
        .I1(\u_ras/u_ras_state/p_1_in10_in ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/p_1_in1_in ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN ),
        .O(\u_ras/w_v0_y [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[1]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[1]_repN ),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[1]_repN ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[1] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v0_y [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[2]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[2] ),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[2] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[2] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v0_y [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[3]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[3] ),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[3] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[3] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v0_y [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[4]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[4] ),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[4] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[4] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v0_y [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[5]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[5] ),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[5]_repN ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[5] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v0_y [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[6]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[6] ),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[6]_repN ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[6]_repN ),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .O(\u_ras/w_v0_y [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[7]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[7] ),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[7]_repN ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[7] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v0_y [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[8]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[8] ),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[8]_repN ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[8] ),
        .I4(\u_ras/u_ras_state/r_state [0]),
        .O(\u_ras/w_v0_y [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y0[9]_i_1 
       (.I0(\u_ras/u_ras_state/r_v0_y_reg_n_0_[9] ),
        .I1(\u_ras/u_ras_state/r_v1_y_reg_n_0_[9] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v2_y_reg_n_0_[9] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v0_y [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y1[0]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[0]_repN ),
        .I1(\u_ras/u_ras_state/r_v2_y_reg_n_0_ ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_ ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v1_y [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y1[10]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[10] ),
        .I1(\u_ras/u_ras_state/r_v2_y_reg_n_0_[10] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_3 ),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[10]_repN ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_3 ),
        .O(\u_ras/w_v1_y [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y1[11]_i_2 
       (.I0(\u_ras/u_ras_state/p_1_in10_in ),
        .I1(\u_ras/u_ras_state/p_1_in1_in ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN_3 ),
        .I3(\u_ras/u_ras_state/p_0_in0_in ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_2 ),
        .O(\u_ras/w_v1_y [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y1[1]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[1] ),
        .I1(\u_ras/u_ras_state/r_v2_y_reg_n_0_[1] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[1] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v1_y [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y1[2]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[2] ),
        .I1(\u_ras/u_ras_state/r_v2_y_reg_n_0_[2] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[2] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v1_y [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y1[3]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[3] ),
        .I1(\u_ras/u_ras_state/r_v2_y_reg_n_0_[3] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[3] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v1_y [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y1[4]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[4] ),
        .I1(\u_ras/u_ras_state/r_v2_y_reg_n_0_[4] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[4] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v1_y [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y1[5]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[5]_repN ),
        .I1(\u_ras/u_ras_state/r_v2_y_reg_n_0_[5] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[5] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v1_y [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y1[6]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[6]_repN ),
        .I1(\u_ras/u_ras_state/r_v2_y_reg_n_0_[6]_repN ),
        .I2(\u_ras/u_ras_state/r_state [1]),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[6] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v1_y [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y1[7]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[7]_repN ),
        .I1(\u_ras/u_ras_state/r_v2_y_reg_n_0_[7] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[7] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v1_y [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y1[8]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[8]_repN ),
        .I1(\u_ras/u_ras_state/r_v2_y_reg_n_0_[8] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[8] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v1_y [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFA0ACFC0)) 
    \u_ras/u_ras_state/r_y1[9]_i_1 
       (.I0(\u_ras/u_ras_state/r_v1_y_reg_n_0_[9] ),
        .I1(\u_ras/u_ras_state/r_v2_y_reg_n_0_[9] ),
        .I2(\u_ras/u_ras_state/r_state[1]_repN ),
        .I3(\u_ras/u_ras_state/r_v0_y_reg_n_0_[9] ),
        .I4(\u_ras/u_ras_state/r_state[0]_repN_4 ),
        .O(\u_ras/w_v1_y [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_state/result3_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_state/result3_carry_n_0 ,\u_ras/u_ras_state/result3_carry_n_1 ,\u_ras/u_ras_state/result3_carry_n_2 ,\u_ras/u_ras_state/result3_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({result3_carry_i_1_n_0,result3_carry_i_2_n_0,result3_carry_i_3_n_0,result3_carry_i_4_n_0}),
        .S({result3_carry_i_5_n_0,result3_carry_i_6_n_0,result3_carry_i_7_n_0,result3_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_state/result3_carry__0 
       (.CI(\u_ras/u_ras_state/result3_carry_n_0 ),
        .CO({\u_ras/u_ras_state/result324_in ,\u_ras/u_ras_state/result3_carry__0_n_1 ,\u_ras/u_ras_state/result3_carry__0_n_2 ,\u_ras/u_ras_state/result3_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,result3_carry__0_i_1_n_0,result3_carry__0_i_2_n_0}),
        .S({result3_carry__0_i_3_n_0,result3_carry__0_i_4_n_0,result3_carry__0_i_5_n_0,result3_carry__0_i_6_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_state/result3_inferred__0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_state/result3_inferred__0_carry_n_0 ,\u_ras/u_ras_state/result3_inferred__0_carry_n_1 ,\u_ras/u_ras_state/result3_inferred__0_carry_n_2 ,\u_ras/u_ras_state/result3_inferred__0_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({result3_inferred__0_carry_i_1_n_0,result3_inferred__0_carry_i_2_n_0,result3_inferred__0_carry_i_3_n_0,result3_inferred__0_carry_i_4_n_0}),
        .S({result3_inferred__0_carry_i_5_n_0,result3_inferred__0_carry_i_6_n_0,result3_inferred__0_carry_i_7_n_0,result3_inferred__0_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_state/result3_inferred__0_carry__0 
       (.CI(\u_ras/u_ras_state/result3_inferred__0_carry_n_0 ),
        .CO({\u_ras/u_ras_state/result327_in ,\u_ras/u_ras_state/result3_inferred__0_carry__0_n_1 ,\u_ras/u_ras_state/result3_inferred__0_carry__0_n_2 ,\u_ras/u_ras_state/result3_inferred__0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,result3_inferred__0_carry__0_i_1_n_0,result3_inferred__0_carry__0_i_2_n_0}),
        .S({result3_inferred__0_carry__0_i_3_n_0,result3_inferred__0_carry__0_i_4_n_0,result3_inferred__0_carry__0_i_5_n_0,result3_inferred__0_carry__0_i_6_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_state/result3_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_state/result3_inferred__1_carry_n_0 ,\u_ras/u_ras_state/result3_inferred__1_carry_n_1 ,\u_ras/u_ras_state/result3_inferred__1_carry_n_2 ,\u_ras/u_ras_state/result3_inferred__1_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({result3_inferred__1_carry_i_1_n_0,result3_inferred__1_carry_i_2_n_0,result3_inferred__1_carry_i_3_n_0,result3_inferred__1_carry_i_4_n_0}),
        .S({result3_inferred__1_carry_i_5_n_0,result3_inferred__1_carry_i_6_n_0,result3_inferred__1_carry_i_7_n_0,result3_inferred__1_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_state/result3_inferred__1_carry__0 
       (.CI(\u_ras/u_ras_state/result3_inferred__1_carry_n_0 ),
        .CO({\u_ras/u_ras_state/result333_in ,\u_ras/u_ras_state/result3_inferred__1_carry__0_n_1 ,\u_ras/u_ras_state/result3_inferred__1_carry__0_n_2 ,\u_ras/u_ras_state/result3_inferred__1_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,result3_inferred__1_carry__0_i_1_n_0,result3_inferred__1_carry__0_i_2_n_0}),
        .S({result3_inferred__1_carry__0_i_3_n_0,result3_inferred__1_carry__0_i_4_n_0,result3_inferred__1_carry__0_i_5_n_0,result3_inferred__1_carry__0_i_6_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_state/result3_inferred__2_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_state/result3_inferred__2_carry_n_0 ,\u_ras/u_ras_state/result3_inferred__2_carry_n_1 ,\u_ras/u_ras_state/result3_inferred__2_carry_n_2 ,\u_ras/u_ras_state/result3_inferred__2_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({result3_inferred__2_carry_i_1_n_0,result3_inferred__2_carry_i_2_n_0,result3_inferred__2_carry_i_3_n_0,result3_inferred__2_carry_i_4_n_0}),
        .S({result3_inferred__2_carry_i_5_n_0,result3_inferred__2_carry_i_6_n_0,result3_inferred__2_carry_i_7_n_0,result3_inferred__2_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_state/result3_inferred__2_carry__0 
       (.CI(\u_ras/u_ras_state/result3_inferred__2_carry_n_0 ),
        .CO({\u_ras/u_ras_state/result336_in ,\u_ras/u_ras_state/result3_inferred__2_carry__0_n_1 ,\u_ras/u_ras_state/result3_inferred__2_carry__0_n_2 ,\u_ras/u_ras_state/result3_inferred__2_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,result3_inferred__2_carry__0_i_1_n_0,result3_inferred__2_carry__0_i_2_n_0}),
        .S({result3_inferred__2_carry__0_i_3_n_0,result3_inferred__2_carry__0_i_4_n_0,result3_inferred__2_carry__0_i_5_n_0,result3_inferred__2_carry__0_i_6_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_state/result3_inferred__3_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_state/result3_inferred__3_carry_n_0 ,\u_ras/u_ras_state/result3_inferred__3_carry_n_1 ,\u_ras/u_ras_state/result3_inferred__3_carry_n_2 ,\u_ras/u_ras_state/result3_inferred__3_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({result3_inferred__3_carry_i_1_n_0,result3_inferred__3_carry_i_2_n_0,result3_inferred__3_carry_i_3_n_0,result3_inferred__3_carry_i_4_n_0}),
        .S({result3_inferred__3_carry_i_5_n_0,result3_inferred__3_carry_i_6_n_0,result3_inferred__3_carry_i_7_n_0,result3_inferred__3_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_state/result3_inferred__3_carry__0 
       (.CI(\u_ras/u_ras_state/result3_inferred__3_carry_n_0 ),
        .CO({\u_ras/u_ras_state/result3__7 ,\u_ras/u_ras_state/result3_inferred__3_carry__0_n_1 ,\u_ras/u_ras_state/result3_inferred__3_carry__0_n_2 ,\u_ras/u_ras_state/result3_inferred__3_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,result3_inferred__3_carry__0_i_1_n_0,result3_inferred__3_carry__0_i_2_n_0}),
        .S({result3_inferred__3_carry__0_i_3_n_0,result3_inferred__3_carry__0_i_4_n_0,result3_inferred__3_carry__0_i_5_n_0,result3_inferred__3_carry__0_i_6_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_state/result3_inferred__4_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras/u_ras_state/result3_inferred__4_carry_n_0 ,\u_ras/u_ras_state/result3_inferred__4_carry_n_1 ,\u_ras/u_ras_state/result3_inferred__4_carry_n_2 ,\u_ras/u_ras_state/result3_inferred__4_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({result3_inferred__4_carry_i_1_n_0,result3_inferred__4_carry_i_2_n_0,result3_inferred__4_carry_i_3_n_0,result3_inferred__4_carry_i_4_n_0}),
        .S({result3_inferred__4_carry_i_5_n_0,result3_inferred__4_carry_i_6_n_0,result3_inferred__4_carry_i_7_n_0,result3_inferred__4_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \u_ras/u_ras_state/result3_inferred__4_carry__0 
       (.CI(\u_ras/u_ras_state/result3_inferred__4_carry_n_0 ),
        .CO({\u_ras/u_ras_state/result316_in ,\u_ras/u_ras_state/result3_inferred__4_carry__0_n_1 ,\u_ras/u_ras_state/result3_inferred__4_carry__0_n_2 ,\u_ras/u_ras_state/result3_inferred__4_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,result3_inferred__4_carry__0_i_1_n_0,result3_inferred__4_carry__0_i_2_n_0}),
        .S({result3_inferred__4_carry__0_i_3_n_0,result3_inferred__4_carry__0_i_4_n_0,result3_inferred__4_carry__0_i_5_n_0,result3_inferred__4_carry__0_i_6_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u_ras_line/r_state[0]_i_1 
       (.I0(r_state_reg),
        .I1(\u_ras/u_ras_line/r_state_reg_n_0_ ),
        .O(\u_ras_line/r_state ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT5 #(
    .INIT(32'h2AFF2A00)) 
    \u_ras_line/r_state[1]_i_1 
       (.I0(\u_ras/u_ras_line/r_state_reg_n_0_ ),
        .I1(\u_ras/u_ras_line/w_end0__3 ),
        .I2(\u_ras/u_ras_line/w_end00_out ),
        .I3(r_state_reg),
        .I4(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .O(\u_ras_line/r_state[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras_line/r_x0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras_line/r_x0_carry_n_0 ,\u_ras_line/r_x0_carry_n_1 ,\u_ras_line/r_x0_carry_n_2 ,\u_ras_line/r_x0_carry_n_3 }),
        .CYINIT(\u_ras/u_ras_line/r_x_reg_n_0_ ),
        .DI({\u_ras/u_ras_line/r_x_reg_n_0_[3] ,\u_ras/u_ras_line/r_x_reg_n_0_[2] ,\u_ras/u_ras_line/r_x_reg_n_0_[1] ,r_x0_carry_i_1_n_0}),
        .O({\u_ras_line/r_x0_carry_n_4 ,\u_ras_line/r_x0_carry_n_5 ,\u_ras_line/r_x0_carry_n_6 ,\u_ras_line/r_x0_carry_n_7 }),
        .S({r_x0_carry_i_2_n_0,r_x0_carry_i_3_n_0,r_x0_carry_i_4_n_0,r_x0_carry_i_5_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras_line/r_x0_carry__0 
       (.CI(\u_ras_line/r_x0_carry_n_0 ),
        .CO({\u_ras_line/r_x0_carry__0_n_0 ,\u_ras_line/r_x0_carry__0_n_1 ,\u_ras_line/r_x0_carry__0_n_2 ,\u_ras_line/r_x0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\u_ras/u_ras_line/r_x_reg_n_0_[7] ,\u_ras/u_ras_line/r_x_reg_n_0_[6] ,\u_ras/u_ras_line/r_x_reg_n_0_[5] ,\u_ras/u_ras_line/r_x_reg_n_0_[4] }),
        .O({\u_ras_line/r_x0_carry__0_n_4 ,\u_ras_line/r_x0_carry__0_n_5 ,\u_ras_line/r_x0_carry__0_n_6 ,\u_ras_line/r_x0_carry__0_n_7 }),
        .S({r_x0_carry__0_i_1_n_0,r_x0_carry__0_i_2_n_0,r_x0_carry__0_i_3_n_0,r_x0_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras_line/r_x0_carry__1 
       (.CI(\u_ras_line/r_x0_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\u_ras/u_ras_line/r_x_reg_n_0_[9] ,\u_ras/u_ras_line/r_x_reg_n_0_[8] }),
        .O({\u_ras_line/r_x0_carry__1_n_4 ,\u_ras_line/r_x0_carry__1_n_5 ,\u_ras_line/r_x0_carry__1_n_6 ,\u_ras_line/r_x0_carry__1_n_7 }),
        .S({\<const0>__0__0 ,r_x0_carry__1_i_1_n_0,r_x0_carry__1_i_2_n_0,r_x0_carry__1_i_3_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras_line/r_y0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\u_ras_line/r_y0_carry_n_0 ,\u_ras_line/r_y0_carry_n_1 ,\u_ras_line/r_y0_carry_n_2 ,\u_ras_line/r_y0_carry_n_3 }),
        .CYINIT(\u_ras/r_y [0]),
        .DI({\u_ras/r_y [3:1],r_y0_carry_i_1_n_0}),
        .O({\u_ras_line/r_y0_carry_n_4 ,\u_ras_line/r_y0_carry_n_5 ,\u_ras_line/r_y0_carry_n_6 ,\u_ras_line/r_y0_carry_n_7 }),
        .S({r_y0_carry_i_2_n_0,r_y0_carry_i_3_n_0,r_y0_carry_i_4_n_0,r_y0_carry_i_5_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras_line/r_y0_carry__0 
       (.CI(\u_ras_line/r_y0_carry_n_0 ),
        .CO({\u_ras_line/r_y0_carry__0_n_0 ,\u_ras_line/r_y0_carry__0_n_1 ,\u_ras_line/r_y0_carry__0_n_2 ,\u_ras_line/r_y0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\u_ras/r_y [7:4]),
        .O({\u_ras_line/r_y0_carry__0_n_4 ,\u_ras_line/r_y0_carry__0_n_5 ,\u_ras_line/r_y0_carry__0_n_6 ,\u_ras_line/r_y0_carry__0_n_7 }),
        .S({r_y0_carry__0_i_1_n_0,r_y0_carry__0_i_2_n_0,r_y0_carry__0_i_3_n_0,r_y0_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-8 {cell *THIS*}}" *) 
  CARRY4 \u_ras_line/r_y0_carry__1 
       (.CI(\u_ras_line/r_y0_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\u_ras/r_y [9:8]}),
        .O({\u_ras_line/r_y0_carry__1_n_4 ,\u_ras_line/r_y0_carry__1_n_5 ,\u_ras_line/r_y0_carry__1_n_6 ,\u_ras_line/r_y0_carry__1_n_7 }),
        .S({\<const0>__0__0 ,r_y0_carry__1_i_1_n_0,r_y0_carry__1_i_2_n_0,r_y0_carry__1_i_3_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBFFAAAA0800AAAA)) 
    \u_ras_mem/r_x[0]_i_1 
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_ ),
        .I1(\u_ras/w_en_pix ),
        .I2(\u_mem_arb/w_pri__0 ),
        .I3(m_wb_ack_i),
        .I4(\u_ras/u_ras_mem/r_state ),
        .I5(\u_ras/u_ras_mem/r_x [0]),
        .O(\u_ras_mem/r_x ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBFFAAAA0800AAAA)) 
    \u_ras_mem/r_x[1]_i_1 
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[1] ),
        .I1(\u_ras/w_en_pix ),
        .I2(\u_mem_arb/w_pri__0 ),
        .I3(m_wb_ack_i),
        .I4(\u_ras/u_ras_mem/r_state ),
        .I5(\u_ras/u_ras_mem/r_x [1]),
        .O(\u_ras_mem/r_x[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_ccw_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_ccw_i_1_n_0),
        .Q(w_ccw),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[0] 
       (.C(clk_i),
        .CE(\r_dma_size[7]_i_1_n_0 ),
        .D(s_wb_dat_i[0]),
        .Q(w_dma_size[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[10] 
       (.C(clk_i),
        .CE(r_dma_size),
        .D(s_wb_dat_i[10]),
        .Q(w_dma_size[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[11] 
       (.C(clk_i),
        .CE(r_dma_size),
        .D(s_wb_dat_i[11]),
        .Q(w_dma_size[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[12] 
       (.C(clk_i),
        .CE(r_dma_size),
        .D(s_wb_dat_i[12]),
        .Q(w_dma_size[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[13] 
       (.C(clk_i),
        .CE(r_dma_size),
        .D(s_wb_dat_i[13]),
        .Q(w_dma_size[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[14] 
       (.C(clk_i),
        .CE(r_dma_size),
        .D(s_wb_dat_i[14]),
        .Q(w_dma_size[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[15] 
       (.C(clk_i),
        .CE(r_dma_size),
        .D(s_wb_dat_i[15]),
        .Q(w_dma_size[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[1] 
       (.C(clk_i),
        .CE(\r_dma_size[7]_i_1_n_0 ),
        .D(s_wb_dat_i[1]),
        .Q(w_dma_size[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[2] 
       (.C(clk_i),
        .CE(\r_dma_size[7]_i_1_n_0 ),
        .D(s_wb_dat_i[2]),
        .Q(w_dma_size[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[3] 
       (.C(clk_i),
        .CE(\r_dma_size[7]_i_1_n_0 ),
        .D(s_wb_dat_i[3]),
        .Q(w_dma_size[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[4] 
       (.C(clk_i),
        .CE(\r_dma_size[7]_i_1_n_0 ),
        .D(s_wb_dat_i[4]),
        .Q(w_dma_size[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[5] 
       (.C(clk_i),
        .CE(\r_dma_size[7]_i_1_n_0 ),
        .D(s_wb_dat_i[5]),
        .Q(w_dma_size[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[6] 
       (.C(clk_i),
        .CE(\r_dma_size[7]_i_1_n_0 ),
        .D(s_wb_dat_i[6]),
        .Q(w_dma_size[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[7] 
       (.C(clk_i),
        .CE(\r_dma_size[7]_i_1_n_0 ),
        .D(s_wb_dat_i[7]),
        .Q(w_dma_size[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[8] 
       (.C(clk_i),
        .CE(r_dma_size),
        .D(s_wb_dat_i[8]),
        .Q(w_dma_size[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_size_reg[9] 
       (.C(clk_i),
        .CE(r_dma_size),
        .D(s_wb_dat_i[9]),
        .Q(w_dma_size[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_start_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_dma_start_i_1_n_0),
        .Q(w_dma_start),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[0] 
       (.C(clk_i),
        .CE(\r_dma_top_address[5]_i_1_n_0 ),
        .D(s_wb_dat_i[2]),
        .Q(w_dma_top_address[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[10] 
       (.C(clk_i),
        .CE(r_dma_top_address),
        .D(s_wb_dat_i[12]),
        .Q(w_dma_top_address[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[11] 
       (.C(clk_i),
        .CE(r_dma_top_address),
        .D(s_wb_dat_i[13]),
        .Q(w_dma_top_address[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[12] 
       (.C(clk_i),
        .CE(r_dma_top_address),
        .D(s_wb_dat_i[14]),
        .Q(w_dma_top_address[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[13] 
       (.C(clk_i),
        .CE(r_dma_top_address),
        .D(s_wb_dat_i[15]),
        .Q(w_dma_top_address[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[14] 
       (.C(clk_i),
        .CE(\r_dma_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[16]),
        .Q(w_dma_top_address[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[15] 
       (.C(clk_i),
        .CE(\r_dma_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[17]),
        .Q(w_dma_top_address[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[16] 
       (.C(clk_i),
        .CE(\r_dma_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[18]),
        .Q(w_dma_top_address[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[17] 
       (.C(clk_i),
        .CE(\r_dma_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[19]),
        .Q(w_dma_top_address[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[18] 
       (.C(clk_i),
        .CE(\r_dma_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[20]),
        .Q(w_dma_top_address[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[19] 
       (.C(clk_i),
        .CE(\r_dma_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[21]),
        .Q(w_dma_top_address[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[1] 
       (.C(clk_i),
        .CE(\r_dma_top_address[5]_i_1_n_0 ),
        .D(s_wb_dat_i[3]),
        .Q(w_dma_top_address[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[20] 
       (.C(clk_i),
        .CE(\r_dma_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[22]),
        .Q(w_dma_top_address[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[21] 
       (.C(clk_i),
        .CE(\r_dma_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[23]),
        .Q(w_dma_top_address[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[22] 
       (.C(clk_i),
        .CE(\r_dma_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[24]),
        .Q(w_dma_top_address[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[23] 
       (.C(clk_i),
        .CE(\r_dma_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[25]),
        .Q(w_dma_top_address[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[24] 
       (.C(clk_i),
        .CE(\r_dma_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[26]),
        .Q(w_dma_top_address[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[25] 
       (.C(clk_i),
        .CE(\r_dma_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[27]),
        .Q(w_dma_top_address[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[26] 
       (.C(clk_i),
        .CE(\r_dma_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[28]),
        .Q(w_dma_top_address[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[27] 
       (.C(clk_i),
        .CE(\r_dma_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[29]),
        .Q(w_dma_top_address[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[28] 
       (.C(clk_i),
        .CE(\r_dma_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[30]),
        .Q(w_dma_top_address[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[29] 
       (.C(clk_i),
        .CE(\r_dma_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_dma_top_address[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[2] 
       (.C(clk_i),
        .CE(\r_dma_top_address[5]_i_1_n_0 ),
        .D(s_wb_dat_i[4]),
        .Q(w_dma_top_address[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[3] 
       (.C(clk_i),
        .CE(\r_dma_top_address[5]_i_1_n_0 ),
        .D(s_wb_dat_i[5]),
        .Q(w_dma_top_address[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[4] 
       (.C(clk_i),
        .CE(\r_dma_top_address[5]_i_1_n_0 ),
        .D(s_wb_dat_i[6]),
        .Q(w_dma_top_address[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[5] 
       (.C(clk_i),
        .CE(\r_dma_top_address[5]_i_1_n_0 ),
        .D(s_wb_dat_i[7]),
        .Q(w_dma_top_address[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[6] 
       (.C(clk_i),
        .CE(r_dma_top_address),
        .D(s_wb_dat_i[8]),
        .Q(w_dma_top_address[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[7] 
       (.C(clk_i),
        .CE(r_dma_top_address),
        .D(s_wb_dat_i[9]),
        .Q(w_dma_top_address[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[8] 
       (.C(clk_i),
        .CE(r_dma_top_address),
        .D(s_wb_dat_i[10]),
        .Q(w_dma_top_address[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_dma_top_address_reg[9] 
       (.C(clk_i),
        .CE(r_dma_top_address),
        .D(s_wb_dat_i[11]),
        .Q(w_dma_top_address[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_en_cull_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_en_cull_i_1_n_0),
        .Q(w_en_cull),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_int_mask_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_int_mask_i_1_n_0),
        .Q(\u_sys/p_21_in [8]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_int_out_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_int_out_i_1_n_0),
        .Q(int_o),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_int_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_int_i_1_n_0),
        .Q(\u_sys/p_21_in [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[0] 
       (.C(clk_i),
        .CE(\r_m00[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m00[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[10] 
       (.C(clk_i),
        .CE(r_m00),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m00[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[11] 
       (.C(clk_i),
        .CE(r_m00),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m00[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[12] 
       (.C(clk_i),
        .CE(r_m00),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m00[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[13] 
       (.C(clk_i),
        .CE(r_m00),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m00[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[14] 
       (.C(clk_i),
        .CE(r_m00),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m00[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[15] 
       (.C(clk_i),
        .CE(r_m00),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m00[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[16] 
       (.C(clk_i),
        .CE(\r_m00[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m00[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[17] 
       (.C(clk_i),
        .CE(\r_m00[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m00[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[18] 
       (.C(clk_i),
        .CE(\r_m00[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m00[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[19] 
       (.C(clk_i),
        .CE(\r_m00[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m00[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[1] 
       (.C(clk_i),
        .CE(\r_m00[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m00[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[20] 
       (.C(clk_i),
        .CE(\r_m00[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m00[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[21] 
       (.C(clk_i),
        .CE(\r_m00[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m00[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[2] 
       (.C(clk_i),
        .CE(\r_m00[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m00[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[3] 
       (.C(clk_i),
        .CE(\r_m00[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m00[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[4] 
       (.C(clk_i),
        .CE(\r_m00[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m00[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[5] 
       (.C(clk_i),
        .CE(\r_m00[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m00[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[6] 
       (.C(clk_i),
        .CE(\r_m00[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m00[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[7] 
       (.C(clk_i),
        .CE(\r_m00[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m00[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[8] 
       (.C(clk_i),
        .CE(r_m00),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m00[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m00_reg[9] 
       (.C(clk_i),
        .CE(r_m00),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m00[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[0] 
       (.C(clk_i),
        .CE(\r_m01[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m01[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[10] 
       (.C(clk_i),
        .CE(r_m01),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m01[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[11] 
       (.C(clk_i),
        .CE(r_m01),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m01[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[12] 
       (.C(clk_i),
        .CE(r_m01),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m01[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[13] 
       (.C(clk_i),
        .CE(r_m01),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m01[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[14] 
       (.C(clk_i),
        .CE(r_m01),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m01[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[15] 
       (.C(clk_i),
        .CE(r_m01),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m01[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[16] 
       (.C(clk_i),
        .CE(\r_m01[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m01[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[17] 
       (.C(clk_i),
        .CE(\r_m01[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m01[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[18] 
       (.C(clk_i),
        .CE(\r_m01[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m01[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[19] 
       (.C(clk_i),
        .CE(\r_m01[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m01[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[1] 
       (.C(clk_i),
        .CE(\r_m01[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m01[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[20] 
       (.C(clk_i),
        .CE(\r_m01[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m01[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[21] 
       (.C(clk_i),
        .CE(\r_m01[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m01[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[2] 
       (.C(clk_i),
        .CE(\r_m01[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m01[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[3] 
       (.C(clk_i),
        .CE(\r_m01[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m01[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[4] 
       (.C(clk_i),
        .CE(\r_m01[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m01[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[5] 
       (.C(clk_i),
        .CE(\r_m01[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m01[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[6] 
       (.C(clk_i),
        .CE(\r_m01[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m01[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[7] 
       (.C(clk_i),
        .CE(\r_m01[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m01[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[8] 
       (.C(clk_i),
        .CE(r_m01),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m01[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m01_reg[9] 
       (.C(clk_i),
        .CE(r_m01),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m01[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[0] 
       (.C(clk_i),
        .CE(\r_m02[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m02[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[10] 
       (.C(clk_i),
        .CE(r_m02),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m02[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[11] 
       (.C(clk_i),
        .CE(r_m02),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m02[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[12] 
       (.C(clk_i),
        .CE(r_m02),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m02[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[13] 
       (.C(clk_i),
        .CE(r_m02),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m02[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[14] 
       (.C(clk_i),
        .CE(r_m02),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m02[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[15] 
       (.C(clk_i),
        .CE(r_m02),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m02[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[16] 
       (.C(clk_i),
        .CE(\r_m02[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m02[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[17] 
       (.C(clk_i),
        .CE(\r_m02[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m02[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[18] 
       (.C(clk_i),
        .CE(\r_m02[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m02[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[19] 
       (.C(clk_i),
        .CE(\r_m02[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m02[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[1] 
       (.C(clk_i),
        .CE(\r_m02[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m02[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[20] 
       (.C(clk_i),
        .CE(\r_m02[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m02[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[21] 
       (.C(clk_i),
        .CE(\r_m02[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m02[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[2] 
       (.C(clk_i),
        .CE(\r_m02[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m02[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[3] 
       (.C(clk_i),
        .CE(\r_m02[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m02[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[4] 
       (.C(clk_i),
        .CE(\r_m02[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m02[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[5] 
       (.C(clk_i),
        .CE(\r_m02[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m02[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[6] 
       (.C(clk_i),
        .CE(\r_m02[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m02[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[7] 
       (.C(clk_i),
        .CE(\r_m02[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m02[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[8] 
       (.C(clk_i),
        .CE(r_m02),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m02[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m02_reg[9] 
       (.C(clk_i),
        .CE(r_m02),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m02[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[0] 
       (.C(clk_i),
        .CE(\r_m03[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m03[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[10] 
       (.C(clk_i),
        .CE(r_m03),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m03[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[11] 
       (.C(clk_i),
        .CE(r_m03),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m03[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[12] 
       (.C(clk_i),
        .CE(r_m03),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m03[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[13] 
       (.C(clk_i),
        .CE(r_m03),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m03[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[14] 
       (.C(clk_i),
        .CE(r_m03),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m03[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[15] 
       (.C(clk_i),
        .CE(r_m03),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m03[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[16] 
       (.C(clk_i),
        .CE(\r_m03[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m03[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[17] 
       (.C(clk_i),
        .CE(\r_m03[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m03[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[18] 
       (.C(clk_i),
        .CE(\r_m03[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m03[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[19] 
       (.C(clk_i),
        .CE(\r_m03[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m03[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[1] 
       (.C(clk_i),
        .CE(\r_m03[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m03[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[20] 
       (.C(clk_i),
        .CE(\r_m03[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m03[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[21] 
       (.C(clk_i),
        .CE(\r_m03[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m03[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[2] 
       (.C(clk_i),
        .CE(\r_m03[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m03[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[3] 
       (.C(clk_i),
        .CE(\r_m03[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m03[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[4] 
       (.C(clk_i),
        .CE(\r_m03[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m03[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[5] 
       (.C(clk_i),
        .CE(\r_m03[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m03[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[6] 
       (.C(clk_i),
        .CE(\r_m03[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m03[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[7] 
       (.C(clk_i),
        .CE(\r_m03[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m03[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[8] 
       (.C(clk_i),
        .CE(r_m03),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m03[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m03_reg[9] 
       (.C(clk_i),
        .CE(r_m03),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m03[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[0] 
       (.C(clk_i),
        .CE(\r_m10[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m10[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[10] 
       (.C(clk_i),
        .CE(r_m10),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m10[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[11] 
       (.C(clk_i),
        .CE(r_m10),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m10[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[12] 
       (.C(clk_i),
        .CE(r_m10),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m10[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[13] 
       (.C(clk_i),
        .CE(r_m10),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m10[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[14] 
       (.C(clk_i),
        .CE(r_m10),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m10[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[15] 
       (.C(clk_i),
        .CE(r_m10),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m10[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[16] 
       (.C(clk_i),
        .CE(\r_m10[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m10[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[17] 
       (.C(clk_i),
        .CE(\r_m10[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m10[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[18] 
       (.C(clk_i),
        .CE(\r_m10[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m10[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[19] 
       (.C(clk_i),
        .CE(\r_m10[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m10[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[1] 
       (.C(clk_i),
        .CE(\r_m10[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m10[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[20] 
       (.C(clk_i),
        .CE(\r_m10[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m10[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[21] 
       (.C(clk_i),
        .CE(\r_m10[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m10[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[2] 
       (.C(clk_i),
        .CE(\r_m10[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m10[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[3] 
       (.C(clk_i),
        .CE(\r_m10[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m10[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[4] 
       (.C(clk_i),
        .CE(\r_m10[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m10[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[5] 
       (.C(clk_i),
        .CE(\r_m10[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m10[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[6] 
       (.C(clk_i),
        .CE(\r_m10[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m10[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[7] 
       (.C(clk_i),
        .CE(\r_m10[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m10[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[8] 
       (.C(clk_i),
        .CE(r_m10),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m10[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m10_reg[9] 
       (.C(clk_i),
        .CE(r_m10),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m10[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[0] 
       (.C(clk_i),
        .CE(\r_m11[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m11[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[10] 
       (.C(clk_i),
        .CE(r_m11),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m11[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[11] 
       (.C(clk_i),
        .CE(r_m11),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m11[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[12] 
       (.C(clk_i),
        .CE(r_m11),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m11[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[13] 
       (.C(clk_i),
        .CE(r_m11),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m11[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[14] 
       (.C(clk_i),
        .CE(r_m11),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m11[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[15] 
       (.C(clk_i),
        .CE(r_m11),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m11[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[16] 
       (.C(clk_i),
        .CE(\r_m11[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m11[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[17] 
       (.C(clk_i),
        .CE(\r_m11[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m11[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[18] 
       (.C(clk_i),
        .CE(\r_m11[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m11[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[19] 
       (.C(clk_i),
        .CE(\r_m11[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m11[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[1] 
       (.C(clk_i),
        .CE(\r_m11[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m11[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[20] 
       (.C(clk_i),
        .CE(\r_m11[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m11[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[21] 
       (.C(clk_i),
        .CE(\r_m11[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m11[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[2] 
       (.C(clk_i),
        .CE(\r_m11[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m11[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[3] 
       (.C(clk_i),
        .CE(\r_m11[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m11[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[4] 
       (.C(clk_i),
        .CE(\r_m11[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m11[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[5] 
       (.C(clk_i),
        .CE(\r_m11[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m11[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[6] 
       (.C(clk_i),
        .CE(\r_m11[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m11[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[7] 
       (.C(clk_i),
        .CE(\r_m11[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m11[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[8] 
       (.C(clk_i),
        .CE(r_m11),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m11[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m11_reg[9] 
       (.C(clk_i),
        .CE(r_m11),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m11[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[0] 
       (.C(clk_i),
        .CE(\r_m12[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m12[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[10] 
       (.C(clk_i),
        .CE(r_m12),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m12[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[11] 
       (.C(clk_i),
        .CE(r_m12),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m12[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[12] 
       (.C(clk_i),
        .CE(r_m12),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m12[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[13] 
       (.C(clk_i),
        .CE(r_m12),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m12[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[14] 
       (.C(clk_i),
        .CE(r_m12),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m12[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[15] 
       (.C(clk_i),
        .CE(r_m12),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m12[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[16] 
       (.C(clk_i),
        .CE(\r_m12[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m12[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[17] 
       (.C(clk_i),
        .CE(\r_m12[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m12[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[18] 
       (.C(clk_i),
        .CE(\r_m12[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m12[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[19] 
       (.C(clk_i),
        .CE(\r_m12[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m12[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[1] 
       (.C(clk_i),
        .CE(\r_m12[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m12[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[20] 
       (.C(clk_i),
        .CE(\r_m12[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m12[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[21] 
       (.C(clk_i),
        .CE(\r_m12[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m12[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[2] 
       (.C(clk_i),
        .CE(\r_m12[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m12[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[3] 
       (.C(clk_i),
        .CE(\r_m12[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m12[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[4] 
       (.C(clk_i),
        .CE(\r_m12[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m12[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[5] 
       (.C(clk_i),
        .CE(\r_m12[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m12[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[6] 
       (.C(clk_i),
        .CE(\r_m12[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m12[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[7] 
       (.C(clk_i),
        .CE(\r_m12[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m12[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[8] 
       (.C(clk_i),
        .CE(r_m12),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m12[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m12_reg[9] 
       (.C(clk_i),
        .CE(r_m12),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m12[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[0] 
       (.C(clk_i),
        .CE(\r_m13[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m13[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[10] 
       (.C(clk_i),
        .CE(r_m13),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m13[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[11] 
       (.C(clk_i),
        .CE(r_m13),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m13[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[12] 
       (.C(clk_i),
        .CE(r_m13),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m13[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[13] 
       (.C(clk_i),
        .CE(r_m13),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m13[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[14] 
       (.C(clk_i),
        .CE(r_m13),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m13[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[15] 
       (.C(clk_i),
        .CE(r_m13),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m13[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[16] 
       (.C(clk_i),
        .CE(\r_m13[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m13[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[17] 
       (.C(clk_i),
        .CE(\r_m13[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m13[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[18] 
       (.C(clk_i),
        .CE(\r_m13[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m13[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[19] 
       (.C(clk_i),
        .CE(\r_m13[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m13[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[1] 
       (.C(clk_i),
        .CE(\r_m13[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m13[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[20] 
       (.C(clk_i),
        .CE(\r_m13[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m13[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[21] 
       (.C(clk_i),
        .CE(\r_m13[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m13[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[2] 
       (.C(clk_i),
        .CE(\r_m13[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m13[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[3] 
       (.C(clk_i),
        .CE(\r_m13[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m13[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[4] 
       (.C(clk_i),
        .CE(\r_m13[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m13[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[5] 
       (.C(clk_i),
        .CE(\r_m13[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m13[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[6] 
       (.C(clk_i),
        .CE(\r_m13[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m13[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[7] 
       (.C(clk_i),
        .CE(\r_m13[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m13[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[8] 
       (.C(clk_i),
        .CE(r_m13),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m13[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m13_reg[9] 
       (.C(clk_i),
        .CE(r_m13),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m13[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[0] 
       (.C(clk_i),
        .CE(\r_m20[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m20[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[10] 
       (.C(clk_i),
        .CE(r_m20),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m20[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[11] 
       (.C(clk_i),
        .CE(r_m20),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m20[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[12] 
       (.C(clk_i),
        .CE(r_m20),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m20[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[13] 
       (.C(clk_i),
        .CE(r_m20),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m20[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[14] 
       (.C(clk_i),
        .CE(r_m20),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m20[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[15] 
       (.C(clk_i),
        .CE(r_m20),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m20[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[16] 
       (.C(clk_i),
        .CE(\r_m20[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m20[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[17] 
       (.C(clk_i),
        .CE(\r_m20[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m20[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[18] 
       (.C(clk_i),
        .CE(\r_m20[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m20[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[19] 
       (.C(clk_i),
        .CE(\r_m20[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m20[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[1] 
       (.C(clk_i),
        .CE(\r_m20[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m20[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[20] 
       (.C(clk_i),
        .CE(\r_m20[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m20[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[21] 
       (.C(clk_i),
        .CE(\r_m20[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m20[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[2] 
       (.C(clk_i),
        .CE(\r_m20[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m20[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[3] 
       (.C(clk_i),
        .CE(\r_m20[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m20[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[4] 
       (.C(clk_i),
        .CE(\r_m20[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m20[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[5] 
       (.C(clk_i),
        .CE(\r_m20[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m20[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[6] 
       (.C(clk_i),
        .CE(\r_m20[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m20[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[7] 
       (.C(clk_i),
        .CE(\r_m20[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m20[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[8] 
       (.C(clk_i),
        .CE(r_m20),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m20[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m20_reg[9] 
       (.C(clk_i),
        .CE(r_m20),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m20[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[0] 
       (.C(clk_i),
        .CE(\r_m21[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m21[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[10] 
       (.C(clk_i),
        .CE(r_m21),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m21[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[11] 
       (.C(clk_i),
        .CE(r_m21),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m21[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[12] 
       (.C(clk_i),
        .CE(r_m21),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m21[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[13] 
       (.C(clk_i),
        .CE(r_m21),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m21[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[14] 
       (.C(clk_i),
        .CE(r_m21),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m21[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[15] 
       (.C(clk_i),
        .CE(r_m21),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m21[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[16] 
       (.C(clk_i),
        .CE(\r_m21[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m21[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[17] 
       (.C(clk_i),
        .CE(\r_m21[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m21[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[18] 
       (.C(clk_i),
        .CE(\r_m21[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m21[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[19] 
       (.C(clk_i),
        .CE(\r_m21[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m21[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[1] 
       (.C(clk_i),
        .CE(\r_m21[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m21[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[20] 
       (.C(clk_i),
        .CE(\r_m21[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m21[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[21] 
       (.C(clk_i),
        .CE(\r_m21[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m21[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[2] 
       (.C(clk_i),
        .CE(\r_m21[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m21[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[3] 
       (.C(clk_i),
        .CE(\r_m21[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m21[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[4] 
       (.C(clk_i),
        .CE(\r_m21[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m21[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[5] 
       (.C(clk_i),
        .CE(\r_m21[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m21[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[6] 
       (.C(clk_i),
        .CE(\r_m21[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m21[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[7] 
       (.C(clk_i),
        .CE(\r_m21[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m21[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[8] 
       (.C(clk_i),
        .CE(r_m21),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m21[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m21_reg[9] 
       (.C(clk_i),
        .CE(r_m21),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m21[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[0] 
       (.C(clk_i),
        .CE(\r_m22[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m22[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[10] 
       (.C(clk_i),
        .CE(r_m22),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m22[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[11] 
       (.C(clk_i),
        .CE(r_m22),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m22[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[12] 
       (.C(clk_i),
        .CE(r_m22),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m22[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[13] 
       (.C(clk_i),
        .CE(r_m22),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m22[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[14] 
       (.C(clk_i),
        .CE(r_m22),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m22[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[15] 
       (.C(clk_i),
        .CE(r_m22),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m22[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[16] 
       (.C(clk_i),
        .CE(\r_m22[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m22[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[17] 
       (.C(clk_i),
        .CE(\r_m22[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m22[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[18] 
       (.C(clk_i),
        .CE(\r_m22[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m22[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[19] 
       (.C(clk_i),
        .CE(\r_m22[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m22[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[1] 
       (.C(clk_i),
        .CE(\r_m22[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m22[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[20] 
       (.C(clk_i),
        .CE(\r_m22[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m22[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[21] 
       (.C(clk_i),
        .CE(\r_m22[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m22[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[2] 
       (.C(clk_i),
        .CE(\r_m22[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m22[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[3] 
       (.C(clk_i),
        .CE(\r_m22[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m22[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[4] 
       (.C(clk_i),
        .CE(\r_m22[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m22[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[5] 
       (.C(clk_i),
        .CE(\r_m22[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m22[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[6] 
       (.C(clk_i),
        .CE(\r_m22[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m22[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[7] 
       (.C(clk_i),
        .CE(\r_m22[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m22[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[8] 
       (.C(clk_i),
        .CE(r_m22),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m22[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m22_reg[9] 
       (.C(clk_i),
        .CE(r_m22),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m22[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[0] 
       (.C(clk_i),
        .CE(\r_m23[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m23[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[10] 
       (.C(clk_i),
        .CE(r_m23),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m23[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[11] 
       (.C(clk_i),
        .CE(r_m23),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m23[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[12] 
       (.C(clk_i),
        .CE(r_m23),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m23[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[13] 
       (.C(clk_i),
        .CE(r_m23),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m23[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[14] 
       (.C(clk_i),
        .CE(r_m23),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m23[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[15] 
       (.C(clk_i),
        .CE(r_m23),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m23[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[16] 
       (.C(clk_i),
        .CE(\r_m23[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m23[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[17] 
       (.C(clk_i),
        .CE(\r_m23[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m23[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[18] 
       (.C(clk_i),
        .CE(\r_m23[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m23[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[19] 
       (.C(clk_i),
        .CE(\r_m23[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m23[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[1] 
       (.C(clk_i),
        .CE(\r_m23[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m23[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[20] 
       (.C(clk_i),
        .CE(\r_m23[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m23[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[21] 
       (.C(clk_i),
        .CE(\r_m23[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m23[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[2] 
       (.C(clk_i),
        .CE(\r_m23[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m23[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[3] 
       (.C(clk_i),
        .CE(\r_m23[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m23[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[4] 
       (.C(clk_i),
        .CE(\r_m23[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m23[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[5] 
       (.C(clk_i),
        .CE(\r_m23[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m23[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[6] 
       (.C(clk_i),
        .CE(\r_m23[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m23[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[7] 
       (.C(clk_i),
        .CE(\r_m23[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m23[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[8] 
       (.C(clk_i),
        .CE(r_m23),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m23[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m23_reg[9] 
       (.C(clk_i),
        .CE(r_m23),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m23[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[0] 
       (.C(clk_i),
        .CE(\r_m30[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m30[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[10] 
       (.C(clk_i),
        .CE(r_m30),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m30[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[11] 
       (.C(clk_i),
        .CE(r_m30),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m30[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[12] 
       (.C(clk_i),
        .CE(r_m30),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m30[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[13] 
       (.C(clk_i),
        .CE(r_m30),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m30[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[14] 
       (.C(clk_i),
        .CE(r_m30),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m30[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[15] 
       (.C(clk_i),
        .CE(r_m30),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m30[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[16] 
       (.C(clk_i),
        .CE(\r_m30[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m30[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[17] 
       (.C(clk_i),
        .CE(\r_m30[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m30[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[18] 
       (.C(clk_i),
        .CE(\r_m30[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m30[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[19] 
       (.C(clk_i),
        .CE(\r_m30[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m30[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[1] 
       (.C(clk_i),
        .CE(\r_m30[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m30[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[20] 
       (.C(clk_i),
        .CE(\r_m30[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m30[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[21] 
       (.C(clk_i),
        .CE(\r_m30[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m30[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[2] 
       (.C(clk_i),
        .CE(\r_m30[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m30[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[3] 
       (.C(clk_i),
        .CE(\r_m30[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m30[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[4] 
       (.C(clk_i),
        .CE(\r_m30[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m30[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[5] 
       (.C(clk_i),
        .CE(\r_m30[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m30[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[6] 
       (.C(clk_i),
        .CE(\r_m30[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m30[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[7] 
       (.C(clk_i),
        .CE(\r_m30[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m30[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[8] 
       (.C(clk_i),
        .CE(r_m30),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m30[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m30_reg[9] 
       (.C(clk_i),
        .CE(r_m30),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m30[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[0] 
       (.C(clk_i),
        .CE(\r_m31[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m31[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[10] 
       (.C(clk_i),
        .CE(r_m31),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m31[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[11] 
       (.C(clk_i),
        .CE(r_m31),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m31[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[12] 
       (.C(clk_i),
        .CE(r_m31),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m31[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[13] 
       (.C(clk_i),
        .CE(r_m31),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m31[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[14] 
       (.C(clk_i),
        .CE(r_m31),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m31[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[15] 
       (.C(clk_i),
        .CE(r_m31),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m31[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[16] 
       (.C(clk_i),
        .CE(\r_m31[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m31[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[17] 
       (.C(clk_i),
        .CE(\r_m31[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m31[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[18] 
       (.C(clk_i),
        .CE(\r_m31[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m31[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[19] 
       (.C(clk_i),
        .CE(\r_m31[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m31[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[1] 
       (.C(clk_i),
        .CE(\r_m31[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m31[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[20] 
       (.C(clk_i),
        .CE(\r_m31[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m31[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[21] 
       (.C(clk_i),
        .CE(\r_m31[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m31[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[2] 
       (.C(clk_i),
        .CE(\r_m31[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m31[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[3] 
       (.C(clk_i),
        .CE(\r_m31[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m31[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[4] 
       (.C(clk_i),
        .CE(\r_m31[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m31[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[5] 
       (.C(clk_i),
        .CE(\r_m31[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m31[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[6] 
       (.C(clk_i),
        .CE(\r_m31[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m31[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[7] 
       (.C(clk_i),
        .CE(\r_m31[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m31[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[8] 
       (.C(clk_i),
        .CE(r_m31),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m31[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m31_reg[9] 
       (.C(clk_i),
        .CE(r_m31),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m31[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[0] 
       (.C(clk_i),
        .CE(\r_m32[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m32[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[10] 
       (.C(clk_i),
        .CE(r_m32),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m32[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[11] 
       (.C(clk_i),
        .CE(r_m32),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m32[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[12] 
       (.C(clk_i),
        .CE(r_m32),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m32[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[13] 
       (.C(clk_i),
        .CE(r_m32),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m32[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[14] 
       (.C(clk_i),
        .CE(r_m32),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m32[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[15] 
       (.C(clk_i),
        .CE(r_m32),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m32[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[16] 
       (.C(clk_i),
        .CE(\r_m32[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m32[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[17] 
       (.C(clk_i),
        .CE(\r_m32[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m32[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[18] 
       (.C(clk_i),
        .CE(\r_m32[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m32[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[19] 
       (.C(clk_i),
        .CE(\r_m32[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m32[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[1] 
       (.C(clk_i),
        .CE(\r_m32[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m32[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[20] 
       (.C(clk_i),
        .CE(\r_m32[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m32[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[21] 
       (.C(clk_i),
        .CE(\r_m32[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m32[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[2] 
       (.C(clk_i),
        .CE(\r_m32[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m32[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[3] 
       (.C(clk_i),
        .CE(\r_m32[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m32[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[4] 
       (.C(clk_i),
        .CE(\r_m32[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m32[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[5] 
       (.C(clk_i),
        .CE(\r_m32[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m32[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[6] 
       (.C(clk_i),
        .CE(\r_m32[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m32[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[7] 
       (.C(clk_i),
        .CE(\r_m32[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m32[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[8] 
       (.C(clk_i),
        .CE(r_m32),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m32[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m32_reg[9] 
       (.C(clk_i),
        .CE(r_m32),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m32[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[0] 
       (.C(clk_i),
        .CE(\r_m33[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_m33[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[10] 
       (.C(clk_i),
        .CE(r_m33),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_m33[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[11] 
       (.C(clk_i),
        .CE(r_m33),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_m33[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[12] 
       (.C(clk_i),
        .CE(r_m33),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_m33[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[13] 
       (.C(clk_i),
        .CE(r_m33),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_m33[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[14] 
       (.C(clk_i),
        .CE(r_m33),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_m33[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[15] 
       (.C(clk_i),
        .CE(r_m33),
        .D(\u_sys/w_f22 [15]),
        .Q(w_m33[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[16] 
       (.C(clk_i),
        .CE(\r_m33[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_m33[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[17] 
       (.C(clk_i),
        .CE(\r_m33[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_m33[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[18] 
       (.C(clk_i),
        .CE(\r_m33[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_m33[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[19] 
       (.C(clk_i),
        .CE(\r_m33[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_m33[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[1] 
       (.C(clk_i),
        .CE(\r_m33[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_m33[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[20] 
       (.C(clk_i),
        .CE(\r_m33[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_m33[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[21] 
       (.C(clk_i),
        .CE(\r_m33[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_m33[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[2] 
       (.C(clk_i),
        .CE(\r_m33[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_m33[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[3] 
       (.C(clk_i),
        .CE(\r_m33[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_m33[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[4] 
       (.C(clk_i),
        .CE(\r_m33[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_m33[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[5] 
       (.C(clk_i),
        .CE(\r_m33[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_m33[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[6] 
       (.C(clk_i),
        .CE(\r_m33[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_m33[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[7] 
       (.C(clk_i),
        .CE(\r_m33[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_m33[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[8] 
       (.C(clk_i),
        .CE(r_m33),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_m33[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_m33_reg[9] 
       (.C(clk_i),
        .CE(r_m33),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_m33[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_color_reg[0] 
       (.C(clk_i),
        .CE(\u_sys/r_pixel_color ),
        .D(s_wb_dat_i[0]),
        .Q(\^m_wb_dat_o [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_color_reg[1] 
       (.C(clk_i),
        .CE(\u_sys/r_pixel_color ),
        .D(s_wb_dat_i[1]),
        .Q(\^m_wb_dat_o [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_color_reg[2] 
       (.C(clk_i),
        .CE(\u_sys/r_pixel_color ),
        .D(s_wb_dat_i[2]),
        .Q(\^m_wb_dat_o [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_color_reg[3] 
       (.C(clk_i),
        .CE(\u_sys/r_pixel_color ),
        .D(s_wb_dat_i[3]),
        .Q(\^m_wb_dat_o [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_color_reg[4] 
       (.C(clk_i),
        .CE(\u_sys/r_pixel_color ),
        .D(s_wb_dat_i[4]),
        .Q(\^m_wb_dat_o [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_color_reg[5] 
       (.C(clk_i),
        .CE(\u_sys/r_pixel_color ),
        .D(s_wb_dat_i[5]),
        .Q(\^m_wb_dat_o [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_color_reg[6] 
       (.C(clk_i),
        .CE(\u_sys/r_pixel_color ),
        .D(s_wb_dat_i[6]),
        .Q(\^m_wb_dat_o [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_color_reg[7] 
       (.C(clk_i),
        .CE(\u_sys/r_pixel_color ),
        .D(s_wb_dat_i[7]),
        .Q(\^m_wb_dat_o [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[0] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[5]_i_1_n_0 ),
        .D(s_wb_dat_i[2]),
        .Q(w_pixel_top_address[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[10] 
       (.C(clk_i),
        .CE(r_pixel_top_address),
        .D(s_wb_dat_i[12]),
        .Q(w_pixel_top_address[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[11] 
       (.C(clk_i),
        .CE(r_pixel_top_address),
        .D(s_wb_dat_i[13]),
        .Q(w_pixel_top_address[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[12] 
       (.C(clk_i),
        .CE(r_pixel_top_address),
        .D(s_wb_dat_i[14]),
        .Q(w_pixel_top_address[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[13] 
       (.C(clk_i),
        .CE(r_pixel_top_address),
        .D(s_wb_dat_i[15]),
        .Q(w_pixel_top_address[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[14] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[16]),
        .Q(w_pixel_top_address[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[15] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[17]),
        .Q(w_pixel_top_address[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[16] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[18]),
        .Q(w_pixel_top_address[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[17] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[19]),
        .Q(w_pixel_top_address[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[18] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[20]),
        .Q(w_pixel_top_address[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[19] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[21]),
        .Q(w_pixel_top_address[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[1] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[5]_i_1_n_0 ),
        .D(s_wb_dat_i[3]),
        .Q(w_pixel_top_address[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[20] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[22]),
        .Q(w_pixel_top_address[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[21] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[21]_i_1_n_0 ),
        .D(s_wb_dat_i[23]),
        .Q(w_pixel_top_address[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[22] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[24]),
        .Q(w_pixel_top_address[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[23] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[25]),
        .Q(w_pixel_top_address[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[24] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[26]),
        .Q(w_pixel_top_address[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[25] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[27]),
        .Q(w_pixel_top_address[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[26] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[28]),
        .Q(w_pixel_top_address[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[27] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[29]),
        .Q(w_pixel_top_address[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[28] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[30]),
        .Q(w_pixel_top_address[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[29] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[29]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_pixel_top_address[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[2] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[5]_i_1_n_0 ),
        .D(s_wb_dat_i[4]),
        .Q(w_pixel_top_address[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[3] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[5]_i_1_n_0 ),
        .D(s_wb_dat_i[5]),
        .Q(w_pixel_top_address[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[4] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[5]_i_1_n_0 ),
        .D(s_wb_dat_i[6]),
        .Q(w_pixel_top_address[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[5] 
       (.C(clk_i),
        .CE(\r_pixel_top_address[5]_i_1_n_0 ),
        .D(s_wb_dat_i[7]),
        .Q(w_pixel_top_address[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[6] 
       (.C(clk_i),
        .CE(r_pixel_top_address),
        .D(s_wb_dat_i[8]),
        .Q(w_pixel_top_address[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[7] 
       (.C(clk_i),
        .CE(r_pixel_top_address),
        .D(s_wb_dat_i[9]),
        .Q(w_pixel_top_address[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[8] 
       (.C(clk_i),
        .CE(r_pixel_top_address),
        .D(s_wb_dat_i[10]),
        .Q(w_pixel_top_address[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_pixel_top_address_reg[9] 
       (.C(clk_i),
        .CE(r_pixel_top_address),
        .D(s_wb_dat_i[11]),
        .Q(w_pixel_top_address[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[0] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[0]_i_1_n_0 ),
        .Q(s_wb_dat_o[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[10] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[10]_i_1_n_0 ),
        .Q(s_wb_dat_o[10]),
        .R(\u_sys/w_rd [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[11] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[11]_i_1_n_0 ),
        .Q(s_wb_dat_o[11]),
        .R(\u_sys/w_rd [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[12] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[12]_i_1_n_0 ),
        .Q(s_wb_dat_o[12]),
        .R(\u_sys/w_rd [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[13] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[13]_i_1_n_0 ),
        .Q(s_wb_dat_o[13]),
        .R(\u_sys/w_rd [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[14] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[14]_i_1_n_0 ),
        .Q(s_wb_dat_o[14]),
        .R(\u_sys/w_rd [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[15] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[15]_i_2_n_0 ),
        .Q(s_wb_dat_o[15]),
        .R(\u_sys/w_rd [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[16] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[16]_i_1_n_0 ),
        .Q(s_wb_dat_o[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[17] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd_reg[17]_i_1_n_0 ),
        .Q(s_wb_dat_o[17]),
        .R(\u_sys/w_rd [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[18] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd_reg[18]_i_1_n_0 ),
        .Q(s_wb_dat_o[18]),
        .R(\u_sys/w_rd [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[19] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd_reg[19]_i_1_n_0 ),
        .Q(s_wb_dat_o[19]),
        .R(\u_sys/w_rd [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[1] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[1]_i_1_n_0 ),
        .Q(s_wb_dat_o[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[20] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd_reg[20]_i_1_n_0 ),
        .Q(s_wb_dat_o[20]),
        .R(\u_sys/w_rd [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[21] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd_reg[21]_i_2_n_0 ),
        .Q(s_wb_dat_o[21]),
        .R(\u_sys/w_rd [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[22] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[22]_i_1_n_0 ),
        .Q(s_wb_dat_o[22]),
        .R(\u_sys/w_rd [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[23] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[23]_i_1_n_0 ),
        .Q(s_wb_dat_o[23]),
        .R(\u_sys/w_rd [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[24] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[24]_i_1_n_0 ),
        .Q(s_wb_dat_o[24]),
        .R(\u_sys/w_rd [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[25] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[25]_i_1_n_0 ),
        .Q(s_wb_dat_o[25]),
        .R(\u_sys/w_rd [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[26] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[26]_i_1_n_0 ),
        .Q(s_wb_dat_o[26]),
        .R(\u_sys/w_rd [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[27] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[27]_i_1_n_0 ),
        .Q(s_wb_dat_o[27]),
        .R(\u_sys/w_rd [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[28] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[28]_i_1_n_0 ),
        .Q(s_wb_dat_o[28]),
        .R(\u_sys/w_rd [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[29] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[29]_i_1_n_0 ),
        .Q(s_wb_dat_o[29]),
        .R(\u_sys/w_rd [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[2] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[2]_i_1_n_0 ),
        .Q(s_wb_dat_o[2]),
        .R(\u_sys/w_rd [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[30] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[30]_i_1_n_0 ),
        .Q(s_wb_dat_o[30]),
        .R(\u_sys/w_rd [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[31] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[31]_i_2_n_0 ),
        .Q(s_wb_dat_o[31]),
        .R(\u_sys/w_rd [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[3] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[3]_i_1_n_0 ),
        .Q(s_wb_dat_o[3]),
        .R(\u_sys/w_rd [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[4] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[4]_i_1_n_0 ),
        .Q(s_wb_dat_o[4]),
        .R(\u_sys/w_rd [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[5] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[5]_i_1_n_0 ),
        .Q(s_wb_dat_o[5]),
        .R(\u_sys/w_rd [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[6] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[6]_i_1_n_0 ),
        .Q(s_wb_dat_o[6]),
        .R(\u_sys/w_rd [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[7] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[7]_i_2_n_0 ),
        .Q(s_wb_dat_o[7]),
        .R(\u_sys/w_rd [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[8] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[8]_i_1_n_0 ),
        .Q(s_wb_dat_o[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rd_reg[9] 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(\r_rd[9]_i_1_n_0 ),
        .Q(s_wb_dat_o[9]),
        .R(\u_sys/w_rd [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_rstr_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_rstr_i_1_n_0),
        .Q(\u_sys/r_rstr ),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[0] 
       (.C(clk_i),
        .CE(\r_scr_h_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[0]),
        .Q(w_scr_h_m1[0]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[10] 
       (.C(clk_i),
        .CE(r_scr_h_m1),
        .D(s_wb_dat_i[10]),
        .Q(w_scr_h_m1[10]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[11] 
       (.C(clk_i),
        .CE(r_scr_h_m1),
        .D(s_wb_dat_i[11]),
        .Q(w_scr_h_m1[11]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[12] 
       (.C(clk_i),
        .CE(r_scr_h_m1),
        .D(s_wb_dat_i[12]),
        .Q(w_scr_h_m1[12]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[13] 
       (.C(clk_i),
        .CE(r_scr_h_m1),
        .D(s_wb_dat_i[13]),
        .Q(w_scr_h_m1[13]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[14] 
       (.C(clk_i),
        .CE(r_scr_h_m1),
        .D(s_wb_dat_i[14]),
        .Q(w_scr_h_m1[14]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[15] 
       (.C(clk_i),
        .CE(r_scr_h_m1),
        .D(s_wb_dat_i[15]),
        .Q(w_scr_h_m1[15]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[1] 
       (.C(clk_i),
        .CE(\r_scr_h_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[1]),
        .Q(w_scr_h_m1[1]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[2] 
       (.C(clk_i),
        .CE(\r_scr_h_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[2]),
        .Q(w_scr_h_m1[2]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[3] 
       (.C(clk_i),
        .CE(\r_scr_h_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[3]),
        .Q(w_scr_h_m1[3]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[4] 
       (.C(clk_i),
        .CE(\r_scr_h_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[4]),
        .Q(w_scr_h_m1[4]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[5] 
       (.C(clk_i),
        .CE(\r_scr_h_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[5]),
        .Q(w_scr_h_m1[5]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[6] 
       (.C(clk_i),
        .CE(\r_scr_h_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[6]),
        .Q(w_scr_h_m1[6]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[7] 
       (.C(clk_i),
        .CE(\r_scr_h_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[7]),
        .Q(w_scr_h_m1[7]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[8] 
       (.C(clk_i),
        .CE(r_scr_h_m1),
        .D(s_wb_dat_i[8]),
        .Q(w_scr_h_m1[8]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_h_m1_reg[9] 
       (.C(clk_i),
        .CE(r_scr_h_m1),
        .D(s_wb_dat_i[9]),
        .Q(w_scr_h_m1[9]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[0] 
       (.C(clk_i),
        .CE(\r_scr_w_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[0]),
        .Q(w_scr_w_m1[0]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[10] 
       (.C(clk_i),
        .CE(r_scr_w_m1),
        .D(s_wb_dat_i[10]),
        .Q(w_scr_w_m1[10]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[11] 
       (.C(clk_i),
        .CE(r_scr_w_m1),
        .D(s_wb_dat_i[11]),
        .Q(w_scr_w_m1[11]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[12] 
       (.C(clk_i),
        .CE(r_scr_w_m1),
        .D(s_wb_dat_i[12]),
        .Q(w_scr_w_m1[12]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[13] 
       (.C(clk_i),
        .CE(r_scr_w_m1),
        .D(s_wb_dat_i[13]),
        .Q(w_scr_w_m1[13]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[14] 
       (.C(clk_i),
        .CE(r_scr_w_m1),
        .D(s_wb_dat_i[14]),
        .Q(w_scr_w_m1[14]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[15] 
       (.C(clk_i),
        .CE(r_scr_w_m1),
        .D(s_wb_dat_i[15]),
        .Q(w_scr_w_m1[15]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[1] 
       (.C(clk_i),
        .CE(\r_scr_w_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[1]),
        .Q(w_scr_w_m1[1]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[2] 
       (.C(clk_i),
        .CE(\r_scr_w_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[2]),
        .Q(w_scr_w_m1[2]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[3] 
       (.C(clk_i),
        .CE(\r_scr_w_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[3]),
        .Q(w_scr_w_m1[3]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[4] 
       (.C(clk_i),
        .CE(\r_scr_w_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[4]),
        .Q(w_scr_w_m1[4]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[5] 
       (.C(clk_i),
        .CE(\r_scr_w_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[5]),
        .Q(w_scr_w_m1[5]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[6] 
       (.C(clk_i),
        .CE(\r_scr_w_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[6]),
        .Q(w_scr_w_m1[6]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[7] 
       (.C(clk_i),
        .CE(\r_scr_w_m1[7]_i_1_n_0 ),
        .D(s_wb_dat_i[7]),
        .Q(w_scr_w_m1[7]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[8] 
       (.C(clk_i),
        .CE(r_scr_w_m1),
        .D(s_wb_dat_i[8]),
        .Q(w_scr_w_m1[8]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_w_m1_reg[9] 
       (.C(clk_i),
        .CE(r_scr_w_m1),
        .D(s_wb_dat_i[9]),
        .Q(w_scr_w_m1[9]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[0] 
       (.C(clk_i),
        .CE(\r_scr_w[7]_i_1_n_0 ),
        .D(s_wb_dat_i[0]),
        .Q(w_scr_w[0]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[10] 
       (.C(clk_i),
        .CE(r_scr_w),
        .D(s_wb_dat_i[10]),
        .Q(w_scr_w[10]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[11] 
       (.C(clk_i),
        .CE(r_scr_w),
        .D(s_wb_dat_i[11]),
        .Q(w_scr_w[11]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[12] 
       (.C(clk_i),
        .CE(r_scr_w),
        .D(s_wb_dat_i[12]),
        .Q(w_scr_w[12]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[13] 
       (.C(clk_i),
        .CE(r_scr_w),
        .D(s_wb_dat_i[13]),
        .Q(w_scr_w[13]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[14] 
       (.C(clk_i),
        .CE(r_scr_w),
        .D(s_wb_dat_i[14]),
        .Q(w_scr_w[14]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[15] 
       (.C(clk_i),
        .CE(r_scr_w),
        .D(s_wb_dat_i[15]),
        .Q(w_scr_w[15]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[1] 
       (.C(clk_i),
        .CE(\r_scr_w[7]_i_1_n_0 ),
        .D(s_wb_dat_i[1]),
        .Q(w_scr_w[1]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[2] 
       (.C(clk_i),
        .CE(\r_scr_w[7]_i_1_n_0 ),
        .D(s_wb_dat_i[2]),
        .Q(w_scr_w[2]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[3] 
       (.C(clk_i),
        .CE(\r_scr_w[7]_i_1_n_0 ),
        .D(s_wb_dat_i[3]),
        .Q(w_scr_w[3]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[4] 
       (.C(clk_i),
        .CE(\r_scr_w[7]_i_1_n_0 ),
        .D(s_wb_dat_i[4]),
        .Q(w_scr_w[4]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[5] 
       (.C(clk_i),
        .CE(\r_scr_w[7]_i_1_n_0 ),
        .D(s_wb_dat_i[5]),
        .Q(w_scr_w[5]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[6] 
       (.C(clk_i),
        .CE(\r_scr_w[7]_i_1_n_0 ),
        .D(s_wb_dat_i[6]),
        .Q(w_scr_w[6]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[7] 
       (.C(clk_i),
        .CE(\r_scr_w[7]_i_1_n_0 ),
        .D(s_wb_dat_i[7]),
        .Q(w_scr_w[7]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[8] 
       (.C(clk_i),
        .CE(r_scr_w),
        .D(s_wb_dat_i[8]),
        .Q(w_scr_w[8]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_scr_w_reg[9] 
       (.C(clk_i),
        .CE(r_scr_w),
        .D(s_wb_dat_i[9]),
        .Q(w_scr_w[9]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[0] 
       (.C(clk_i),
        .CE(\r_vh[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_vh[0]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[10] 
       (.C(clk_i),
        .CE(r_vh),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_vh[10]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[11] 
       (.C(clk_i),
        .CE(r_vh),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_vh[11]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[12] 
       (.C(clk_i),
        .CE(r_vh),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_vh[12]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[13] 
       (.C(clk_i),
        .CE(r_vh),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_vh[13]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[14] 
       (.C(clk_i),
        .CE(r_vh),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_vh[14]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[15] 
       (.C(clk_i),
        .CE(r_vh),
        .D(\u_sys/w_f22 [15]),
        .Q(w_vh[15]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[16] 
       (.C(clk_i),
        .CE(\r_vh[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_vh[16]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[17] 
       (.C(clk_i),
        .CE(\r_vh[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_vh[17]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[18] 
       (.C(clk_i),
        .CE(\r_vh[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_vh[18]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[19] 
       (.C(clk_i),
        .CE(\r_vh[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_vh[19]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[1] 
       (.C(clk_i),
        .CE(\r_vh[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_vh[1]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[20] 
       (.C(clk_i),
        .CE(\r_vh[21]_i_1_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_vh[20]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[21] 
       (.C(clk_i),
        .CE(\r_vh[21]_i_1_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_vh[21]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[2] 
       (.C(clk_i),
        .CE(\r_vh[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_vh[2]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[3] 
       (.C(clk_i),
        .CE(\r_vh[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_vh[3]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[4] 
       (.C(clk_i),
        .CE(\r_vh[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_vh[4]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[5] 
       (.C(clk_i),
        .CE(\r_vh[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_vh[5]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[6] 
       (.C(clk_i),
        .CE(\r_vh[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_vh[6]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[7] 
       (.C(clk_i),
        .CE(\r_vh[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_vh[7]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[8] 
       (.C(clk_i),
        .CE(r_vh),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_vh[8]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vh_reg[9] 
       (.C(clk_i),
        .CE(r_vh),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_vh[9]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[0] 
       (.C(clk_i),
        .CE(\r_vw[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_7 ),
        .Q(w_vw[0]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[10] 
       (.C(clk_i),
        .CE(r_vw),
        .D(\r_m00_reg[11]_i_1_n_5 ),
        .Q(w_vw[10]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[11] 
       (.C(clk_i),
        .CE(r_vw),
        .D(\r_m00_reg[11]_i_1_n_4 ),
        .Q(w_vw[11]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[12] 
       (.C(clk_i),
        .CE(r_vw),
        .D(\r_m00_reg[14]_i_1_n_7 ),
        .Q(w_vw[12]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[13] 
       (.C(clk_i),
        .CE(r_vw),
        .D(\r_m00_reg[14]_i_1_n_6 ),
        .Q(w_vw[13]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[14] 
       (.C(clk_i),
        .CE(r_vw),
        .D(\r_m00_reg[14]_i_1_n_5 ),
        .Q(w_vw[14]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[15] 
       (.C(clk_i),
        .CE(r_vw),
        .D(\u_sys/w_f22 [15]),
        .Q(w_vw[15]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[16] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1__0_n_0 ),
        .D(\u_sys/w_f22 [16]),
        .Q(w_vw[16]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[17] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1__0_n_0 ),
        .D(\u_sys/w_f22 [17]),
        .Q(w_vw[17]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[18] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1__0_n_0 ),
        .D(\u_sys/w_f22 [18]),
        .Q(w_vw[18]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[19] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1__0_n_0 ),
        .D(\u_sys/w_f22 [19]),
        .Q(w_vw[19]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[1] 
       (.C(clk_i),
        .CE(\r_vw[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_6 ),
        .Q(w_vw[1]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[20] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1__0_n_0 ),
        .D(\u_sys/w_f22 [20]),
        .Q(w_vw[20]),
        .S(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[21] 
       (.C(clk_i),
        .CE(\r_vw[21]_i_1__0_n_0 ),
        .D(s_wb_dat_i[31]),
        .Q(w_vw[21]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[2] 
       (.C(clk_i),
        .CE(\r_vw[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_5 ),
        .Q(w_vw[2]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[3] 
       (.C(clk_i),
        .CE(\r_vw[7]_i_1_n_0 ),
        .D(\r_m00_reg[3]_i_1_n_4 ),
        .Q(w_vw[3]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[4] 
       (.C(clk_i),
        .CE(\r_vw[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_7 ),
        .Q(w_vw[4]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[5] 
       (.C(clk_i),
        .CE(\r_vw[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_6 ),
        .Q(w_vw[5]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[6] 
       (.C(clk_i),
        .CE(\r_vw[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_5 ),
        .Q(w_vw[6]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[7] 
       (.C(clk_i),
        .CE(\r_vw[7]_i_1_n_0 ),
        .D(\r_m00_reg[7]_i_2_n_4 ),
        .Q(w_vw[7]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[8] 
       (.C(clk_i),
        .CE(r_vw),
        .D(\r_m00_reg[11]_i_1_n_7 ),
        .Q(w_vw[8]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_vw_reg[9] 
       (.C(clk_i),
        .CE(r_vw),
        .D(\r_m00_reg[11]_i_1_n_6 ),
        .Q(w_vw[9]),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u_sys/r_y_flip_reg 
       (.C(clk_i),
        .CE(\<const1>__0__0 ),
        .D(r_y_flip_i_1_n_0),
        .Q(w_y_flip),
        .R(rst_i));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_1
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [14]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_82 ),
        .O(w_cf_tmp_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_1__0
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [11]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_85 ),
        .O(w_cf_tmp_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_1__1
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [7]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_89 ),
        .O(w_cf_tmp_carry_i_1__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_1__2
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [3]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_93 ),
        .O(w_cf_tmp_carry_i_1__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_2
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [13]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_83 ),
        .O(w_cf_tmp_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_2__0
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [10]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_86 ),
        .O(w_cf_tmp_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_2__1
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [6]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_90 ),
        .O(w_cf_tmp_carry_i_2__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_2__2
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [2]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_94 ),
        .O(w_cf_tmp_carry_i_2__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_3
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [12]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_84 ),
        .O(w_cf_tmp_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_3__0
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [9]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_87 ),
        .O(w_cf_tmp_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_3__1
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [5]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_91 ),
        .O(w_cf_tmp_carry_i_3__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_3__2
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [1]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_95 ),
        .O(w_cf_tmp_carry_i_3__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_4
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [8]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_88 ),
        .O(w_cf_tmp_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_4__0
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [4]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_92 ),
        .O(w_cf_tmp_carry_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_cf_tmp_carry_i_4__1
       (.I0(\u_geo/u_geo_persdiv/w_rom_base [0]),
        .I1(\u_geo/u_geo_persdiv/u_frcp/w_rom_correct_n_96 ),
        .O(w_cf_tmp_carry_i_4__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_1
       (.I0(w_m10[15]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_33_n_0),
        .O(w_cf_tmp_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_10
       (.I0(w_m10[6]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_42_n_0),
        .O(w_cf_tmp_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_10__0
       (.I0(w_m11[6]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_42__0_n_0),
        .O(w_cf_tmp_i_10__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_10__1
       (.I0(w_m12[6]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_42__1_n_0),
        .O(w_cf_tmp_i_10__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_10__2
       (.I0(w_m13[6]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_26_n_0),
        .O(w_cf_tmp_i_10__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_10__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[6] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [6]),
        .O(w_cf_tmp_i_10__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_10__4
       (.I0(w_vw[6]),
        .I1(w_vh[6]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_11
       (.I0(w_m10[5]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_43_n_0),
        .O(w_cf_tmp_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_11__0
       (.I0(w_m11[5]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_43__0_n_0),
        .O(w_cf_tmp_i_11__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_11__1
       (.I0(w_m12[5]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_43__1_n_0),
        .O(w_cf_tmp_i_11__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_11__2
       (.I0(w_m13[5]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_27_n_0),
        .O(w_cf_tmp_i_11__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_11__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[5] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [5]),
        .O(w_cf_tmp_i_11__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_11__4
       (.I0(w_vw[5]),
        .I1(w_vh[5]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_12
       (.I0(w_m10[4]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_44_n_0),
        .O(w_cf_tmp_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_12__0
       (.I0(w_m11[4]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_44__0_n_0),
        .O(w_cf_tmp_i_12__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_12__1
       (.I0(w_m12[4]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_44__1_n_0),
        .O(w_cf_tmp_i_12__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_12__2
       (.I0(w_m13[4]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_28_n_0),
        .O(w_cf_tmp_i_12__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_12__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[4] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [4]),
        .O(w_cf_tmp_i_12__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_12__4
       (.I0(w_vw[4]),
        .I1(w_vh[4]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_13
       (.I0(w_m10[3]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_45_n_0),
        .O(w_cf_tmp_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_13__0
       (.I0(w_m11[3]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_45__0_n_0),
        .O(w_cf_tmp_i_13__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_13__1
       (.I0(w_m12[3]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_45__1_n_0),
        .O(w_cf_tmp_i_13__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_13__2
       (.I0(w_m13[3]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_29_n_0),
        .O(w_cf_tmp_i_13__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_13__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[3] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [3]),
        .O(w_cf_tmp_i_13__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_13__4
       (.I0(w_vw[3]),
        .I1(w_vh[3]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_14
       (.I0(w_m10[2]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_46_n_0),
        .O(w_cf_tmp_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_14__0
       (.I0(w_m11[2]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_46__0_n_0),
        .O(w_cf_tmp_i_14__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_14__1
       (.I0(w_m12[2]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_46__1_n_0),
        .O(w_cf_tmp_i_14__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_14__2
       (.I0(w_m13[2]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_30_n_0),
        .O(w_cf_tmp_i_14__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_14__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[2] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [2]),
        .O(w_cf_tmp_i_14__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_14__4
       (.I0(w_vw[2]),
        .I1(w_vh[2]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_15
       (.I0(w_m10[1]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_47_n_0),
        .O(w_cf_tmp_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_15__0
       (.I0(w_m11[1]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_47__0_n_0),
        .O(w_cf_tmp_i_15__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_15__1
       (.I0(w_m12[1]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_47__1_n_0),
        .O(w_cf_tmp_i_15__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_15__2
       (.I0(w_m13[1]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_31_n_0),
        .O(w_cf_tmp_i_15__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_15__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[1] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [1]),
        .O(w_cf_tmp_i_15__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_15__4
       (.I0(w_vw[1]),
        .I1(w_vh[1]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_16
       (.I0(w_m10[0]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_48_n_0),
        .O(w_cf_tmp_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_16__0
       (.I0(w_m11[0]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_48__0_n_0),
        .O(w_cf_tmp_i_16__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_16__1
       (.I0(w_m12[0]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_48__1_n_0),
        .O(w_cf_tmp_i_16__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_16__2
       (.I0(w_m13[0]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_32_n_0),
        .O(w_cf_tmp_i_16__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_16__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_ ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [0]),
        .O(w_cf_tmp_i_16__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_16__4
       (.I0(w_vw[0]),
        .I1(w_vh[0]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_17
       (.I0(w_m23[15]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[15]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[15]),
        .O(w_cf_tmp_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_17__0
       (.I0(\u_geo/w_vz_dma [15]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [15]),
        .O(\u_geo/u_geo_matrix/w_vz_in [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_17__1
       (.I0(\u_geo/w_vy_dma [15]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [15]),
        .O(\u_geo/u_geo_matrix/w_vy_in [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_17__2
       (.I0(\u_geo/w_vx_dma [15]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [15]),
        .O(\u_geo/u_geo_matrix/w_vx_in [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_17__3
       (.I0(\u_geo/w_vy_pdiv [15]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [15]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF00FF00FF00FE)) 
    w_cf_tmp_i_17__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [0]),
        .I1(\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [2]),
        .I2(\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [1]),
        .I3(\r_c[20]_i_2__8_n_0 ),
        .I4(\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [4]),
        .I5(\u_geo/u_geo_viewport/u_fadd/norm/f_incdec_return [3]),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_18
       (.I0(w_m23[14]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[14]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[14]),
        .O(w_cf_tmp_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_18__0
       (.I0(\u_geo/w_vz_dma [14]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [14]),
        .O(\u_geo/u_geo_matrix/w_vz_in [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_18__1
       (.I0(\u_geo/w_vy_dma [14]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [14]),
        .O(\u_geo/u_geo_matrix/w_vy_in [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_18__2
       (.I0(\u_geo/w_vx_dma [14]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [14]),
        .O(\u_geo/u_geo_matrix/w_vx_in [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_18__3
       (.I0(\u_geo/w_vy_pdiv [14]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [14]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC000E020F0F0F0F0)) 
    w_cf_tmp_i_18__4
       (.I0(w_cf_tmp_i_33__2_n_0),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I2(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [15]),
        .I4(w_cf_tmp_i_34__2_n_0),
        .I5(w_cf_tmp_i_35__2_n_0),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_19
       (.I0(w_m23[13]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[13]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[13]),
        .O(w_cf_tmp_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_19__0
       (.I0(\u_geo/w_vz_dma [13]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [13]),
        .O(\u_geo/u_geo_matrix/w_vz_in [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_19__1
       (.I0(\u_geo/w_vy_dma [13]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [13]),
        .O(\u_geo/u_geo_matrix/w_vy_in [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_19__2
       (.I0(\u_geo/w_vx_dma [13]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [13]),
        .O(\u_geo/u_geo_matrix/w_vx_in [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_19__3
       (.I0(\u_geo/w_vy_pdiv [13]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [13]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88880A0088880AAA)) 
    w_cf_tmp_i_19__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [14]),
        .I2(w_cf_tmp_i_36__2_n_0),
        .I3(w_cf_tmp_i_33__2_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I5(w_cf_tmp_i_34__2_n_0),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_1__0
       (.I0(w_m11[15]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_33__0_n_0),
        .O(w_cf_tmp_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_1__1
       (.I0(w_m12[15]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_33__1_n_0),
        .O(w_cf_tmp_i_1__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_1__2
       (.I0(w_m13[15]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_17_n_0),
        .O(w_cf_tmp_i_1__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_1__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[15] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [15]),
        .O(w_cf_tmp_i_1__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_1__4
       (.I0(w_vw[15]),
        .I1(w_vh[15]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_2
       (.I0(w_m10[14]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_34_n_0),
        .O(w_cf_tmp_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_20
       (.I0(w_m23[12]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[12]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[12]),
        .O(w_cf_tmp_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_20__0
       (.I0(\u_geo/w_vz_dma [12]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [12]),
        .O(\u_geo/u_geo_matrix/w_vz_in [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_20__1
       (.I0(\u_geo/w_vy_dma [12]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [12]),
        .O(\u_geo/u_geo_matrix/w_vy_in [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_20__2
       (.I0(\u_geo/w_vx_dma [12]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [12]),
        .O(\u_geo/u_geo_matrix/w_vx_in [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_20__3
       (.I0(\u_geo/w_vy_pdiv [12]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [12]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88880A0088880AAA)) 
    w_cf_tmp_i_20__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [13]),
        .I2(w_cf_tmp_i_37__2_n_0),
        .I3(w_cf_tmp_i_33__2_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I5(w_cf_tmp_i_36__2_n_0),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_21
       (.I0(w_m23[11]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[11]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[11]),
        .O(w_cf_tmp_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_21__0
       (.I0(\u_geo/w_vz_dma [11]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [11]),
        .O(\u_geo/u_geo_matrix/w_vz_in [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_21__1
       (.I0(\u_geo/w_vy_dma [11]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [11]),
        .O(\u_geo/u_geo_matrix/w_vy_in [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_21__2
       (.I0(\u_geo/w_vx_dma [11]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [11]),
        .O(\u_geo/u_geo_matrix/w_vx_in [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_21__3
       (.I0(\u_geo/w_vy_pdiv [11]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [11]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8800880A88AA880A)) 
    w_cf_tmp_i_21__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [12]),
        .I2(w_cf_tmp_i_37__2_n_0),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I4(w_cf_tmp_i_33__2_n_0),
        .I5(w_cf_tmp_i_38__2_n_0),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_22
       (.I0(w_m23[10]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[10]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[10]),
        .O(w_cf_tmp_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_22__0
       (.I0(\u_geo/w_vz_dma [10]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [10]),
        .O(\u_geo/u_geo_matrix/w_vz_in [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_22__1
       (.I0(\u_geo/w_vy_dma [10]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [10]),
        .O(\u_geo/u_geo_matrix/w_vy_in [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_22__2
       (.I0(\u_geo/w_vx_dma [10]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [10]),
        .O(\u_geo/u_geo_matrix/w_vx_in [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_22__3
       (.I0(\u_geo/w_vy_pdiv [10]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [10]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA02A2000002A2)) 
    w_cf_tmp_i_22__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(w_cf_tmp_i_38__2_n_0),
        .I2(w_cf_tmp_i_33__2_n_0),
        .I3(w_cf_tmp_i_39__2_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I5(\u_geo/u_geo_viewport/u_fadd/r_mats [11]),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_23
       (.I0(w_m23[9]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[9]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[9]),
        .O(w_cf_tmp_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_23__0
       (.I0(\u_geo/w_vz_dma [9]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [9]),
        .O(\u_geo/u_geo_matrix/w_vz_in [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_23__1
       (.I0(\u_geo/w_vy_dma [9]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [9]),
        .O(\u_geo/u_geo_matrix/w_vy_in [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_23__2
       (.I0(\u_geo/w_vx_dma [9]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [9]),
        .O(\u_geo/u_geo_matrix/w_vx_in [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_23__3
       (.I0(\u_geo/w_vy_pdiv [9]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [9]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88880A0088880AAA)) 
    w_cf_tmp_i_23__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [10]),
        .I2(w_cf_tmp_i_40__2_n_0),
        .I3(w_cf_tmp_i_33__2_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I5(w_cf_tmp_i_39__2_n_0),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_24
       (.I0(w_m23[8]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[8]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[8]),
        .O(w_cf_tmp_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_24__0
       (.I0(\u_geo/w_vz_dma [8]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [8]),
        .O(\u_geo/u_geo_matrix/w_vz_in [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_24__1
       (.I0(\u_geo/w_vy_dma [8]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [8]),
        .O(\u_geo/u_geo_matrix/w_vy_in [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_24__2
       (.I0(\u_geo/w_vx_dma [8]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [8]),
        .O(\u_geo/u_geo_matrix/w_vx_in [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_24__3
       (.I0(\u_geo/w_vy_pdiv [8]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [8]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA02A2000002A2)) 
    w_cf_tmp_i_24__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(w_cf_tmp_i_40__2_n_0),
        .I2(w_cf_tmp_i_33__2_n_0),
        .I3(w_cf_tmp_i_41__2_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I5(\u_geo/u_geo_viewport/u_fadd/r_mats [9]),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_25
       (.I0(w_m23[7]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[7]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[7]),
        .O(w_cf_tmp_i_25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_25__0
       (.I0(\u_geo/w_vz_dma [7]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [7]),
        .O(\u_geo/u_geo_matrix/w_vz_in [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_25__1
       (.I0(\u_geo/w_vy_dma [7]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [7]),
        .O(\u_geo/u_geo_matrix/w_vy_in [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_25__2
       (.I0(\u_geo/w_vx_dma [7]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [7]),
        .O(\u_geo/u_geo_matrix/w_vx_in [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_25__3
       (.I0(\u_geo/w_vy_pdiv [7]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [7]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8800880A88AA880A)) 
    w_cf_tmp_i_25__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [8]),
        .I2(w_cf_tmp_i_41__2_n_0),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I4(w_cf_tmp_i_33__2_n_0),
        .I5(w_cf_tmp_i_42__2_n_0),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_26
       (.I0(w_m23[6]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[6]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[6]),
        .O(w_cf_tmp_i_26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_26__0
       (.I0(\u_geo/w_vz_dma [6]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [6]),
        .O(\u_geo/u_geo_matrix/w_vz_in [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_26__1
       (.I0(\u_geo/w_vy_dma [6]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [6]),
        .O(\u_geo/u_geo_matrix/w_vy_in [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_26__2
       (.I0(\u_geo/w_vx_dma [6]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [6]),
        .O(\u_geo/u_geo_matrix/w_vx_in [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_26__3
       (.I0(\u_geo/w_vy_pdiv [6]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [6]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8800880A88AA880A)) 
    w_cf_tmp_i_26__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [7]),
        .I2(w_cf_tmp_i_42__2_n_0),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I4(w_cf_tmp_i_33__2_n_0),
        .I5(w_cf_tmp_i_43__2_n_0),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_27
       (.I0(w_m23[5]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[5]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[5]),
        .O(w_cf_tmp_i_27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_27__0
       (.I0(\u_geo/w_vz_dma [5]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [5]),
        .O(\u_geo/u_geo_matrix/w_vz_in [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_27__1
       (.I0(\u_geo/w_vy_dma [5]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [5]),
        .O(\u_geo/u_geo_matrix/w_vy_in [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_27__2
       (.I0(\u_geo/w_vx_dma [5]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [5]),
        .O(\u_geo/u_geo_matrix/w_vx_in [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_27__3
       (.I0(\u_geo/w_vy_pdiv [5]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [5]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA02A2000002A2)) 
    w_cf_tmp_i_27__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(w_cf_tmp_i_43__2_n_0),
        .I2(w_cf_tmp_i_33__2_n_0),
        .I3(w_cf_tmp_i_44__2_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I5(\u_geo/u_geo_viewport/u_fadd/r_mats [6]),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_28
       (.I0(w_m23[4]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[4]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[4]),
        .O(w_cf_tmp_i_28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_28__0
       (.I0(\u_geo/w_vz_dma [4]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [4]),
        .O(\u_geo/u_geo_matrix/w_vz_in [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_28__1
       (.I0(\u_geo/w_vy_dma [4]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [4]),
        .O(\u_geo/u_geo_matrix/w_vy_in [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_28__2
       (.I0(\u_geo/w_vx_dma [4]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [4]),
        .O(\u_geo/u_geo_matrix/w_vx_in [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_28__3
       (.I0(\u_geo/w_vy_pdiv [4]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [4]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA02A2000002A2)) 
    w_cf_tmp_i_28__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(w_cf_tmp_i_44__2_n_0),
        .I2(w_cf_tmp_i_33__2_n_0),
        .I3(w_cf_tmp_i_45__2_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I5(\u_geo/u_geo_viewport/u_fadd/r_mats [5]),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_29
       (.I0(w_m23[3]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[3]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[3]),
        .O(w_cf_tmp_i_29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_29__0
       (.I0(\u_geo/w_vz_dma [3]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [3]),
        .O(\u_geo/u_geo_matrix/w_vz_in [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_29__1
       (.I0(\u_geo/w_vy_dma [3]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [3]),
        .O(\u_geo/u_geo_matrix/w_vy_in [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_29__2
       (.I0(\u_geo/w_vx_dma [3]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [3]),
        .O(\u_geo/u_geo_matrix/w_vx_in [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_29__3
       (.I0(\u_geo/w_vy_pdiv [3]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [3]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA02A2000002A2)) 
    w_cf_tmp_i_29__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(w_cf_tmp_i_45__2_n_0),
        .I2(w_cf_tmp_i_33__2_n_0),
        .I3(w_cf_tmp_i_46__2_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I5(\u_geo/u_geo_viewport/u_fadd/r_mats [4]),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_2__0
       (.I0(w_m11[14]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_34__0_n_0),
        .O(w_cf_tmp_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_2__1
       (.I0(w_m12[14]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_34__1_n_0),
        .O(w_cf_tmp_i_2__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_2__2
       (.I0(w_m13[14]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_18_n_0),
        .O(w_cf_tmp_i_2__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_2__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[14] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [14]),
        .O(w_cf_tmp_i_2__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_2__4
       (.I0(w_vw[14]),
        .I1(w_vh[14]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_3
       (.I0(w_m10[13]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_35_n_0),
        .O(w_cf_tmp_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_30
       (.I0(w_m23[2]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[2]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[2]),
        .O(w_cf_tmp_i_30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_30__0
       (.I0(\u_geo/w_vz_dma [2]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [2]),
        .O(\u_geo/u_geo_matrix/w_vz_in [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_30__1
       (.I0(\u_geo/w_vy_dma [2]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [2]),
        .O(\u_geo/u_geo_matrix/w_vy_in [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_30__2
       (.I0(\u_geo/w_vx_dma [2]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [2]),
        .O(\u_geo/u_geo_matrix/w_vx_in [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_30__3
       (.I0(\u_geo/w_vy_pdiv [2]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [2]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA008080AA00A2A2)) 
    w_cf_tmp_i_30__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(w_cf_tmp_i_33__2_n_0),
        .I2(w_cf_tmp_i_47__2_n_0),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [3]),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I5(w_cf_tmp_i_46__2_n_0),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_31
       (.I0(w_m23[1]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[1]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[1]),
        .O(w_cf_tmp_i_31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_31__0
       (.I0(\u_geo/w_vz_dma [1]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [1]),
        .O(\u_geo/u_geo_matrix/w_vz_in [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_31__1
       (.I0(\u_geo/w_vy_dma [1]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [1]),
        .O(\u_geo/u_geo_matrix/w_vy_in [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_31__2
       (.I0(\u_geo/w_vx_dma [1]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [1]),
        .O(\u_geo/u_geo_matrix/w_vx_in [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_31__3
       (.I0(\u_geo/w_vy_pdiv [1]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [1]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    w_cf_tmp_i_31__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I1(w_cf_tmp_i_48__2_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [2]),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_32
       (.I0(w_m23[0]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m33[0]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m03[0]),
        .O(w_cf_tmp_i_32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_32__0
       (.I0(\u_geo/w_vz_dma [0]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vz_in [0]),
        .O(\u_geo/u_geo_matrix/w_vz_in [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_32__1
       (.I0(\u_geo/w_vy_dma [0]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vy_in [0]),
        .O(\u_geo/u_geo_matrix/w_vy_in [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_32__2
       (.I0(\u_geo/w_vx_dma [0]),
        .I1(\u_geo/w_state_mat ),
        .I2(\u_geo/u_geo_matrix/r_vx_in [0]),
        .O(\u_geo/u_geo_matrix/w_vx_in [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAABAAA8A)) 
    w_cf_tmp_i_32__3
       (.I0(\u_geo/w_vy_pdiv [0]),
        .I1(\u_geo/u_geo_persdiv/r_state [0]),
        .I2(\u_geo/u_geo_persdiv/r_state [1]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/w_vx_pdiv [0]),
        .O(\u_geo/u_geo_persdiv/w_fmul_a [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB010A000)) 
    w_cf_tmp_i_32__4
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I1(w_cf_tmp_i_33__2_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/w_c [15]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [1]),
        .I4(w_cf_tmp_i_49_n_0),
        .O(\u_geo/u_geo_viewport/u_fadd/w_c [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_33
       (.I0(w_m20[15]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[15]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[15]),
        .O(w_cf_tmp_i_33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_33__0
       (.I0(w_m21[15]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[15]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[15]),
        .O(w_cf_tmp_i_33__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_33__1
       (.I0(w_m22[15]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[15]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[15]),
        .O(w_cf_tmp_i_33__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000F000F0000000E)) 
    w_cf_tmp_i_33__2
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [6]),
        .I1(w_cf_tmp_i_50_n_0),
        .I2(w_cf_tmp_i_51_n_0),
        .I3(w_cf_tmp_i_52_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [7]),
        .I5(w_cf_tmp_i_53_n_0),
        .O(w_cf_tmp_i_33__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_34
       (.I0(w_m20[14]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[14]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[14]),
        .O(w_cf_tmp_i_34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_34__0
       (.I0(w_m21[14]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[14]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[14]),
        .O(w_cf_tmp_i_34__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_34__1
       (.I0(w_m22[14]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[14]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[14]),
        .O(w_cf_tmp_i_34__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_34__2
       (.I0(w_cf_tmp_i_54_n_0),
        .I1(_inferred__1_carry_i_8__8_n_0),
        .I2(w_cf_tmp_i_55_n_0),
        .O(w_cf_tmp_i_34__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_35
       (.I0(w_m20[13]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[13]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[13]),
        .O(w_cf_tmp_i_35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_35__0
       (.I0(w_m21[13]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[13]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[13]),
        .O(w_cf_tmp_i_35__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_35__1
       (.I0(w_m22[13]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[13]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[13]),
        .O(w_cf_tmp_i_35__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEFEEEE)) 
    w_cf_tmp_i_35__2
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [16]),
        .I1(w_cf_tmp_i_33__2_n_0),
        .I2(_inferred__1_carry_i_8__8_n_0),
        .I3(w_cf_tmp_i_56_n_0),
        .I4(w_cf_tmp_i_57_n_0),
        .O(w_cf_tmp_i_35__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_36
       (.I0(w_m20[12]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[12]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[12]),
        .O(w_cf_tmp_i_36_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_36__0
       (.I0(w_m21[12]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[12]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[12]),
        .O(w_cf_tmp_i_36__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_36__1
       (.I0(w_m22[12]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[12]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[12]),
        .O(w_cf_tmp_i_36__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_36__2
       (.I0(w_cf_tmp_i_58_n_0),
        .I1(_inferred__1_carry_i_8__8_n_0),
        .I2(w_cf_tmp_i_56_n_0),
        .O(w_cf_tmp_i_36__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_37
       (.I0(w_m20[11]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[11]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[11]),
        .O(w_cf_tmp_i_37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_37__0
       (.I0(w_m21[11]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[11]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[11]),
        .O(w_cf_tmp_i_37__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_37__1
       (.I0(w_m22[11]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[11]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[11]),
        .O(w_cf_tmp_i_37__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_37__2
       (.I0(w_cf_tmp_i_59_n_0),
        .I1(_inferred__1_carry_i_8__8_n_0),
        .I2(w_cf_tmp_i_54_n_0),
        .O(w_cf_tmp_i_37__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_38
       (.I0(w_m20[10]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[10]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[10]),
        .O(w_cf_tmp_i_38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_38__0
       (.I0(w_m21[10]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[10]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[10]),
        .O(w_cf_tmp_i_38__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_38__1
       (.I0(w_m22[10]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[10]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[10]),
        .O(w_cf_tmp_i_38__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_38__2
       (.I0(w_cf_tmp_i_60_n_0),
        .I1(_inferred__1_carry_i_8__8_n_0),
        .I2(w_cf_tmp_i_58_n_0),
        .O(w_cf_tmp_i_38__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_39
       (.I0(w_m20[9]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[9]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[9]),
        .O(w_cf_tmp_i_39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_39__0
       (.I0(w_m21[9]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[9]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[9]),
        .O(w_cf_tmp_i_39__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_39__1
       (.I0(w_m22[9]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[9]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[9]),
        .O(w_cf_tmp_i_39__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    w_cf_tmp_i_39__2
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [3]),
        .I1(_inferred__1_carry_i_7__8_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [7]),
        .I3(_inferred__1_carry_i_6__8_n_0),
        .I4(_inferred__1_carry_i_8__8_n_0),
        .I5(w_cf_tmp_i_59_n_0),
        .O(w_cf_tmp_i_39__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_3__0
       (.I0(w_m11[13]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_35__0_n_0),
        .O(w_cf_tmp_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_3__1
       (.I0(w_m12[13]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_35__1_n_0),
        .O(w_cf_tmp_i_3__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_3__2
       (.I0(w_m13[13]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_19_n_0),
        .O(w_cf_tmp_i_3__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_3__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[13] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [13]),
        .O(w_cf_tmp_i_3__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_3__4
       (.I0(w_vw[13]),
        .I1(w_vh[13]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_4
       (.I0(w_m10[12]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_36_n_0),
        .O(w_cf_tmp_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_40
       (.I0(w_m20[8]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[8]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[8]),
        .O(w_cf_tmp_i_40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_40__0
       (.I0(w_m21[8]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[8]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[8]),
        .O(w_cf_tmp_i_40__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_40__1
       (.I0(w_m22[8]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[8]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[8]),
        .O(w_cf_tmp_i_40__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    w_cf_tmp_i_40__2
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [2]),
        .I1(_inferred__1_carry_i_7__8_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [6]),
        .I3(_inferred__1_carry_i_6__8_n_0),
        .I4(_inferred__1_carry_i_8__8_n_0),
        .I5(w_cf_tmp_i_60_n_0),
        .O(w_cf_tmp_i_40__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_41
       (.I0(w_m20[7]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[7]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[7]),
        .O(w_cf_tmp_i_41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_41__0
       (.I0(w_m21[7]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[7]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[7]),
        .O(w_cf_tmp_i_41__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_41__1
       (.I0(w_m22[7]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[7]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[7]),
        .O(w_cf_tmp_i_41__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    w_cf_tmp_i_41__2
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [1]),
        .I1(_inferred__1_carry_i_7__8_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [5]),
        .I3(_inferred__1_carry_i_6__8_n_0),
        .I4(_inferred__1_carry_i_8__8_n_0),
        .I5(w_cf_tmp_i_61_n_0),
        .O(w_cf_tmp_i_41__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_42
       (.I0(w_m20[6]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[6]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[6]),
        .O(w_cf_tmp_i_42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_42__0
       (.I0(w_m21[6]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[6]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[6]),
        .O(w_cf_tmp_i_42__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_42__1
       (.I0(w_m22[6]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[6]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[6]),
        .O(w_cf_tmp_i_42__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47FFFFFF47FF0000)) 
    w_cf_tmp_i_42__2
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [0]),
        .I1(_inferred__1_carry_i_7__8_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [4]),
        .I3(_inferred__1_carry_i_6__8_n_0),
        .I4(_inferred__1_carry_i_8__8_n_0),
        .I5(w_cf_tmp_i_62_n_0),
        .O(w_cf_tmp_i_42__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_43
       (.I0(w_m20[5]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[5]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[5]),
        .O(w_cf_tmp_i_43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_43__0
       (.I0(w_m21[5]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[5]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[5]),
        .O(w_cf_tmp_i_43__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_43__1
       (.I0(w_m22[5]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[5]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[5]),
        .O(w_cf_tmp_i_43__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    w_cf_tmp_i_43__2
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [3]),
        .I1(_inferred__1_carry_i_8__8_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [1]),
        .I3(_inferred__1_carry_i_7__8_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [5]),
        .I5(_inferred__1_carry_i_6__8_n_0),
        .O(w_cf_tmp_i_43__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_44
       (.I0(w_m20[4]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[4]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[4]),
        .O(w_cf_tmp_i_44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_44__0
       (.I0(w_m21[4]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[4]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[4]),
        .O(w_cf_tmp_i_44__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_44__1
       (.I0(w_m22[4]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[4]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[4]),
        .O(w_cf_tmp_i_44__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    w_cf_tmp_i_44__2
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [2]),
        .I1(_inferred__1_carry_i_8__8_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [0]),
        .I3(_inferred__1_carry_i_7__8_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [4]),
        .I5(_inferred__1_carry_i_6__8_n_0),
        .O(w_cf_tmp_i_44__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_45
       (.I0(w_m20[3]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[3]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[3]),
        .O(w_cf_tmp_i_45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_45__0
       (.I0(w_m21[3]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[3]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[3]),
        .O(w_cf_tmp_i_45__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_45__1
       (.I0(w_m22[3]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[3]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[3]),
        .O(w_cf_tmp_i_45__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    w_cf_tmp_i_45__2
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [1]),
        .I1(_inferred__1_carry_i_8__8_n_0),
        .I2(_inferred__1_carry_i_7__8_n_0),
        .I3(_inferred__1_carry_i_6__8_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [3]),
        .O(w_cf_tmp_i_45__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_46
       (.I0(w_m20[2]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[2]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[2]),
        .O(w_cf_tmp_i_46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_46__0
       (.I0(w_m21[2]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[2]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[2]),
        .O(w_cf_tmp_i_46__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_46__1
       (.I0(w_m22[2]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[2]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[2]),
        .O(w_cf_tmp_i_46__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF4FFF7FF)) 
    w_cf_tmp_i_46__2
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [0]),
        .I1(_inferred__1_carry_i_8__8_n_0),
        .I2(_inferred__1_carry_i_7__8_n_0),
        .I3(_inferred__1_carry_i_6__8_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [2]),
        .O(w_cf_tmp_i_46__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_47
       (.I0(w_m20[1]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[1]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[1]),
        .O(w_cf_tmp_i_47_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_47__0
       (.I0(w_m21[1]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[1]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[1]),
        .O(w_cf_tmp_i_47__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_47__1
       (.I0(w_m22[1]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[1]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[1]),
        .O(w_cf_tmp_i_47__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    w_cf_tmp_i_47__2
       (.I0(_inferred__1_carry_i_8__8_n_0),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [1]),
        .I2(_inferred__1_carry_i_6__8_n_0),
        .I3(_inferred__1_carry_i_7__8_n_0),
        .O(w_cf_tmp_i_47__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_48
       (.I0(w_m20[0]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m30[0]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m00[0]),
        .O(w_cf_tmp_i_48_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_48__0
       (.I0(w_m21[0]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m31[0]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m01[0]),
        .O(w_cf_tmp_i_48__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    w_cf_tmp_i_48__1
       (.I0(w_m22[0]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[2] ),
        .I2(w_m32[0]),
        .I3(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_[3] ),
        .I4(w_m02[0]),
        .O(w_cf_tmp_i_48__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000B080000)) 
    w_cf_tmp_i_48__2
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [0]),
        .I1(w_cf_tmp_i_33__2_n_0),
        .I2(_inferred__1_carry_i_8__8_n_0),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [1]),
        .I4(_inferred__1_carry_i_6__8_n_0),
        .I5(_inferred__1_carry_i_7__8_n_0),
        .O(w_cf_tmp_i_48__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    w_cf_tmp_i_49
       (.I0(_inferred__1_carry_i_8__8_n_0),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [0]),
        .I2(_inferred__1_carry_i_6__8_n_0),
        .I3(_inferred__1_carry_i_7__8_n_0),
        .O(w_cf_tmp_i_49_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_4__0
       (.I0(w_m11[12]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_36__0_n_0),
        .O(w_cf_tmp_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_4__1
       (.I0(w_m12[12]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_36__1_n_0),
        .O(w_cf_tmp_i_4__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_4__2
       (.I0(w_m13[12]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_20_n_0),
        .O(w_cf_tmp_i_4__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_4__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[12] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [12]),
        .O(w_cf_tmp_i_4__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_4__4
       (.I0(w_vw[12]),
        .I1(w_vh[12]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_5
       (.I0(w_m10[11]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_37_n_0),
        .O(w_cf_tmp_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551011)) 
    w_cf_tmp_i_50
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [5]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [3]),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [2]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [1]),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [4]),
        .O(w_cf_tmp_i_50_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    w_cf_tmp_i_51
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [9]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [12]),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [14]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [10]),
        .O(w_cf_tmp_i_51_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00F4)) 
    w_cf_tmp_i_52
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [12]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [11]),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [13]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [14]),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [15]),
        .O(w_cf_tmp_i_52_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    w_cf_tmp_i_53
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [8]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [12]),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [14]),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [10]),
        .O(w_cf_tmp_i_53_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    w_cf_tmp_i_54
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [7]),
        .I1(_inferred__1_carry_i_7__8_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [11]),
        .I3(_inferred__1_carry_i_6__8_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [3]),
        .O(w_cf_tmp_i_54_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505010105F5F101F)) 
    w_cf_tmp_i_55
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [9]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [1]),
        .I2(_inferred__1_carry_i_7__8_n_0),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [5]),
        .I4(_inferred__1_carry_i_6__8_n_0),
        .I5(\u_geo/u_geo_viewport/u_fadd/r_mats [13]),
        .O(w_cf_tmp_i_55_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h303010103F3F101F)) 
    w_cf_tmp_i_56
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [0]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [8]),
        .I2(_inferred__1_carry_i_7__8_n_0),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [4]),
        .I4(_inferred__1_carry_i_6__8_n_0),
        .I5(\u_geo/u_geo_viewport/u_fadd/r_mats [12]),
        .O(w_cf_tmp_i_56_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h303010103F3F101F)) 
    w_cf_tmp_i_57
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [2]),
        .I1(\u_geo/u_geo_viewport/u_fadd/r_mats [10]),
        .I2(_inferred__1_carry_i_7__8_n_0),
        .I3(\u_geo/u_geo_viewport/u_fadd/r_mats [6]),
        .I4(_inferred__1_carry_i_6__8_n_0),
        .I5(\u_geo/u_geo_viewport/u_fadd/r_mats [14]),
        .O(w_cf_tmp_i_57_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44CC77CF)) 
    w_cf_tmp_i_58
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [6]),
        .I1(_inferred__1_carry_i_7__8_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [2]),
        .I3(_inferred__1_carry_i_6__8_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [10]),
        .O(w_cf_tmp_i_58_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h47CC47CF)) 
    w_cf_tmp_i_59
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [5]),
        .I1(_inferred__1_carry_i_7__8_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [9]),
        .I3(_inferred__1_carry_i_6__8_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [1]),
        .O(w_cf_tmp_i_59_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_5__0
       (.I0(w_m11[11]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_37__0_n_0),
        .O(w_cf_tmp_i_5__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_5__1
       (.I0(w_m12[11]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_37__1_n_0),
        .O(w_cf_tmp_i_5__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_5__2
       (.I0(w_m13[11]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_21_n_0),
        .O(w_cf_tmp_i_5__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_5__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[11] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [11]),
        .O(w_cf_tmp_i_5__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_5__4
       (.I0(w_vw[11]),
        .I1(w_vh[11]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_6
       (.I0(w_m10[10]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_38_n_0),
        .O(w_cf_tmp_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44CC77CF)) 
    w_cf_tmp_i_60
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [4]),
        .I1(_inferred__1_carry_i_7__8_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [0]),
        .I3(_inferred__1_carry_i_6__8_n_0),
        .I4(\u_geo/u_geo_viewport/u_fadd/r_mats [8]),
        .O(w_cf_tmp_i_60_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    w_cf_tmp_i_61
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [3]),
        .I1(_inferred__1_carry_i_7__8_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [7]),
        .I3(_inferred__1_carry_i_6__8_n_0),
        .O(w_cf_tmp_i_61_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h47FF)) 
    w_cf_tmp_i_62
       (.I0(\u_geo/u_geo_viewport/u_fadd/r_mats [2]),
        .I1(_inferred__1_carry_i_7__8_n_0),
        .I2(\u_geo/u_geo_viewport/u_fadd/r_mats [6]),
        .I3(_inferred__1_carry_i_6__8_n_0),
        .O(w_cf_tmp_i_62_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_6__0
       (.I0(w_m11[10]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_38__0_n_0),
        .O(w_cf_tmp_i_6__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_6__1
       (.I0(w_m12[10]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_38__1_n_0),
        .O(w_cf_tmp_i_6__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_6__2
       (.I0(w_m13[10]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_22_n_0),
        .O(w_cf_tmp_i_6__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_6__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[10] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [10]),
        .O(w_cf_tmp_i_6__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_6__4
       (.I0(w_vw[10]),
        .I1(w_vh[10]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_7
       (.I0(w_m10[9]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_39_n_0),
        .O(w_cf_tmp_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_7__0
       (.I0(w_m11[9]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_39__0_n_0),
        .O(w_cf_tmp_i_7__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_7__1
       (.I0(w_m12[9]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_39__1_n_0),
        .O(w_cf_tmp_i_7__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_7__2
       (.I0(w_m13[9]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_23_n_0),
        .O(w_cf_tmp_i_7__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_7__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[9] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [9]),
        .O(w_cf_tmp_i_7__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_7__4
       (.I0(w_vw[9]),
        .I1(w_vh[9]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_8
       (.I0(w_m10[8]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_40_n_0),
        .O(w_cf_tmp_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_8__0
       (.I0(w_m11[8]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_40__0_n_0),
        .O(w_cf_tmp_i_8__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_8__1
       (.I0(w_m12[8]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_40__1_n_0),
        .O(w_cf_tmp_i_8__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_8__2
       (.I0(w_m13[8]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_24_n_0),
        .O(w_cf_tmp_i_8__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_8__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[8] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [8]),
        .O(w_cf_tmp_i_8__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_8__4
       (.I0(w_vw[8]),
        .I1(w_vh[8]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_9
       (.I0(w_m10[7]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_41_n_0),
        .O(w_cf_tmp_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_9__0
       (.I0(w_m11[7]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_41__0_n_0),
        .O(w_cf_tmp_i_9__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_9__1
       (.I0(w_m12[7]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_41__1_n_0),
        .O(w_cf_tmp_i_9__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_cf_tmp_i_9__2
       (.I0(w_m13[7]),
        .I1(\u_geo/u_geo_matrix/FSM_onehot_r_state_reg_n_0_ ),
        .I2(w_cf_tmp_i_25_n_0),
        .O(w_cf_tmp_i_9__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFB0008)) 
    w_cf_tmp_i_9__3
       (.I0(\u_geo/u_geo_persdiv/u_frcp/r_c_reg_n_0_[7] ),
        .I1(\u_geo/u_geo_persdiv/r_state [1]),
        .I2(\u_geo/u_geo_persdiv/r_state [0]),
        .I3(\u_geo/u_geo_persdiv/r_state [2]),
        .I4(\u_geo/u_geo_persdiv/r_ivw [7]),
        .O(w_cf_tmp_i_9__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCACCCCCCCCCCCC)) 
    w_cf_tmp_i_9__4
       (.I0(w_vw[7]),
        .I1(w_vh[7]),
        .I2(\u_geo/u_geo_viewport/r_state [2]),
        .I3(\u_geo/u_geo_viewport/r_state [3]),
        .I4(\u_geo/u_geo_viewport/r_state [1]),
        .I5(\u_geo/u_geo_viewport/r_state [0]),
        .O(\u_geo/u_geo_viewport/w_fmul_b [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    w_dym_carry__0_i_1
       (.I0(\u_ras/w_dy [7]),
        .O(w_dym_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    w_dym_carry__0_i_2
       (.I0(\u_ras/w_dy [6]),
        .O(w_dym_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    w_dym_carry__0_i_3
       (.I0(\u_ras/w_dy [5]),
        .O(w_dym_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    w_dym_carry__0_i_4
       (.I0(\u_ras/w_dy [4]),
        .O(w_dym_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    w_dym_carry__1_i_1
       (.I0(\u_ras/w_dy [11]),
        .O(w_dym_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    w_dym_carry__1_i_2
       (.I0(\u_ras/w_dy [10]),
        .O(w_dym_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    w_dym_carry__1_i_3
       (.I0(\u_ras/w_dy [9]),
        .O(w_dym_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    w_dym_carry__1_i_4
       (.I0(\u_ras/w_dy [8]),
        .O(w_dym_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    w_dym_carry_i_1
       (.I0(\u_ras/w_dy [3]),
        .O(w_dym_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    w_dym_carry_i_2
       (.I0(\u_ras/w_dy [2]),
        .O(w_dym_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    w_dym_carry_i_3
       (.I0(\u_ras/w_dy [1]),
        .O(w_dym_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    w_end0_carry_i_1
       (.I0(\u_ras/r_y [9]),
        .I1(\u_ras/w_y1 [9]),
        .I2(\u_ras/w_y1 [11]),
        .I3(\u_ras/w_y ),
        .I4(\u_ras/w_y1 [10]),
        .I5(\u_ras/r_y [10]),
        .O(w_end0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    w_end0_carry_i_2
       (.I0(\u_ras/r_y [6]),
        .I1(\u_ras/w_y1 [6]),
        .I2(\u_ras/w_y1 [8]),
        .I3(\u_ras/r_y [8]),
        .I4(\u_ras/w_y1 [7]),
        .I5(\u_ras/r_y [7]),
        .O(w_end0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    w_end0_carry_i_3
       (.I0(\u_ras/r_y [3]),
        .I1(\u_ras/w_y1 [3]),
        .I2(\u_ras/w_y1 [5]),
        .I3(\u_ras/r_y [5]),
        .I4(\u_ras/w_y1 [4]),
        .I5(\u_ras/r_y [4]),
        .O(w_end0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    w_end0_carry_i_4
       (.I0(\u_ras/r_y [0]),
        .I1(\u_ras/w_y1 [0]),
        .I2(\u_ras/w_y1 [2]),
        .I3(\u_ras/r_y [2]),
        .I4(\u_ras/w_y1 [1]),
        .I5(\u_ras/r_y [1]),
        .O(w_end0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    w_end0_inferred__0_carry_i_1
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[9] ),
        .I1(\u_ras/w_x1 [9]),
        .I2(\u_ras/w_x1 [11]),
        .I3(\u_ras/w_x ),
        .I4(\u_ras/w_x1 [10]),
        .I5(\u_ras/u_ras_line/r_x_reg_n_0_[10] ),
        .O(w_end0_inferred__0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    w_end0_inferred__0_carry_i_2
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[6] ),
        .I1(\u_ras/w_x1 [6]),
        .I2(\u_ras/w_x1 [8]),
        .I3(\u_ras/u_ras_line/r_x_reg_n_0_[8] ),
        .I4(\u_ras/w_x1 [7]),
        .I5(\u_ras/u_ras_line/r_x_reg_n_0_[7] ),
        .O(w_end0_inferred__0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    w_end0_inferred__0_carry_i_3
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[3] ),
        .I1(\u_ras/w_x1 [3]),
        .I2(\u_ras/w_x1 [5]),
        .I3(\u_ras/u_ras_line/r_x_reg_n_0_[5] ),
        .I4(\u_ras/w_x1 [4]),
        .I5(\u_ras/u_ras_line/r_x_reg_n_0_[4] ),
        .O(w_end0_inferred__0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    w_end0_inferred__0_carry_i_4
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_ ),
        .I1(\u_ras/w_x1 [0]),
        .I2(\u_ras/w_x1 [2]),
        .I3(\u_ras/u_ras_line/r_x_reg_n_0_[2] ),
        .I4(\u_ras/w_x1 [1]),
        .I5(\u_ras/u_ras_line/r_x_reg_n_0_[1] ),
        .O(w_end0_inferred__0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair5" *) 
  LUT3 #(
    .INIT(8'hD4)) 
    w_err__0_carry__0_i_1
       (.I0(\u_ras/w_dy [6]),
        .I1(w_err__0_carry__0_i_9_n_0),
        .I2(\u_ras/p_2_in [6]),
        .O(w_err__0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    w_err__0_carry__0_i_10
       (.I0(\u_ras/u_ras_line/r_x1 [5]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x0 [5]),
        .I3(w_err__0_carry__0_i_14_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(w_err__0_carry__0_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    w_err__0_carry__0_i_11
       (.I0(\u_ras/u_ras_line/r_x1 [4]),
        .I1(_inferred__5_carry_i_9_n_0_repN),
        .I2(\u_ras/u_ras_line/r_x0 [4]),
        .I3(w_err__0_carry__0_i_15_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(w_err__0_carry__0_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    w_err__0_carry__0_i_12
       (.I0(\u_ras/u_ras_line/r_x1 [7]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x0 [7]),
        .I3(w_err__0_carry__0_i_16_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(w_err__0_carry__0_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    w_err__0_carry__0_i_13
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_v0_x_reg_n_0_[6] ),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[6] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[6] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(w_err__0_carry__0_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    w_err__0_carry__0_i_14
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_v0_x_reg_n_0_[5] ),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[5] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[5] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(w_err__0_carry__0_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    w_err__0_carry__0_i_15
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_v0_x_reg_n_0_[4] ),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[4] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[4] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(w_err__0_carry__0_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    w_err__0_carry__0_i_16
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_v0_x_reg_n_0_[7] ),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[7] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[7] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(w_err__0_carry__0_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair4" *) 
  LUT3 #(
    .INIT(8'hD4)) 
    w_err__0_carry__0_i_2
       (.I0(\u_ras/w_dy [5]),
        .I1(w_err__0_carry__0_i_10_n_0),
        .I2(\u_ras/p_2_in [5]),
        .O(w_err__0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair3" *) 
  LUT3 #(
    .INIT(8'hD4)) 
    w_err__0_carry__0_i_3
       (.I0(\u_ras/w_dy [4]),
        .I1(w_err__0_carry__0_i_11_n_0),
        .I2(\u_ras/p_2_in [4]),
        .O(w_err__0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair2" *) 
  LUT3 #(
    .INIT(8'hD4)) 
    w_err__0_carry__0_i_4
       (.I0(\u_ras/w_dy [3]),
        .I1(w_err__0_carry_i_11_n_0),
        .I2(\u_ras/p_2_in [3]),
        .O(w_err__0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair6" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    w_err__0_carry__0_i_5
       (.I0(\u_ras/w_dy [7]),
        .I1(w_err__0_carry__0_i_12_n_0),
        .I2(\u_ras/p_2_in [7]),
        .I3(w_err__0_carry__0_i_1_n_0),
        .O(w_err__0_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair5" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    w_err__0_carry__0_i_6
       (.I0(\u_ras/w_dy [6]),
        .I1(w_err__0_carry__0_i_9_n_0),
        .I2(\u_ras/p_2_in [6]),
        .I3(w_err__0_carry__0_i_2_n_0),
        .O(w_err__0_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair4" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    w_err__0_carry__0_i_7
       (.I0(\u_ras/w_dy [5]),
        .I1(w_err__0_carry__0_i_10_n_0),
        .I2(\u_ras/p_2_in [5]),
        .I3(w_err__0_carry__0_i_3_n_0),
        .O(w_err__0_carry__0_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair3" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    w_err__0_carry__0_i_8
       (.I0(\u_ras/w_dy [4]),
        .I1(w_err__0_carry__0_i_11_n_0),
        .I2(\u_ras/p_2_in [4]),
        .I3(w_err__0_carry__0_i_4_n_0),
        .O(w_err__0_carry__0_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    w_err__0_carry__0_i_9
       (.I0(\u_ras/u_ras_line/r_x1 [6]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x0 [6]),
        .I3(w_err__0_carry__0_i_13_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(w_err__0_carry__0_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair7" *) 
  LUT3 #(
    .INIT(8'hD4)) 
    w_err__0_carry__1_i_1
       (.I0(\u_ras/w_dy [8]),
        .I1(w_err__0_carry__1_i_6_n_0),
        .I2(\u_ras/p_2_in [8]),
        .O(w_err__0_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    w_err__0_carry__1_i_10
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_v0_x_reg_n_0_[9] ),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[9] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[9] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(w_err__0_carry__1_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    w_err__0_carry__1_i_11
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_v0_x_reg_n_0_[10] ),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[10] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[10] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(w_err__0_carry__1_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair6" *) 
  LUT3 #(
    .INIT(8'hD4)) 
    w_err__0_carry__1_i_2
       (.I0(\u_ras/w_dy [7]),
        .I1(w_err__0_carry__0_i_12_n_0),
        .I2(\u_ras/p_2_in [7]),
        .O(w_err__0_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8E71718E718E8E71)) 
    w_err__0_carry__1_i_3
       (.I0(\u_ras/p_2_in [9]),
        .I1(w_err__0_carry__1_i_7_n_0),
        .I2(\u_ras/w_dy [9]),
        .I3(\u_ras/w_dy [10]),
        .I4(w_err__0_carry__1_i_8_n_0),
        .I5(\u_ras/p_2_in [10]),
        .O(w_err__0_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    w_err__0_carry__1_i_4
       (.I0(w_err__0_carry__1_i_1_n_0),
        .I1(\u_ras/w_dy [9]),
        .I2(w_err__0_carry__1_i_7_n_0),
        .I3(\u_ras/p_2_in [9]),
        .O(w_err__0_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair7" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    w_err__0_carry__1_i_5
       (.I0(\u_ras/w_dy [8]),
        .I1(w_err__0_carry__1_i_6_n_0),
        .I2(\u_ras/p_2_in [8]),
        .I3(w_err__0_carry__1_i_2_n_0),
        .O(w_err__0_carry__1_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    w_err__0_carry__1_i_6
       (.I0(\u_ras/u_ras_line/r_x1 [8]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x0 [8]),
        .I3(w_err__0_carry__1_i_9_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(w_err__0_carry__1_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    w_err__0_carry__1_i_7
       (.I0(\u_ras/u_ras_line/r_x1 [9]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x0 [9]),
        .I3(w_err__0_carry__1_i_10_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(w_err__0_carry__1_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    w_err__0_carry__1_i_8
       (.I0(\u_ras/u_ras_line/r_x1 [10]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x0 [10]),
        .I3(w_err__0_carry__1_i_11_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(w_err__0_carry__1_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    w_err__0_carry__1_i_9
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_v0_x_reg_n_0_[8] ),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[8] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[8] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(w_err__0_carry__1_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair1" *) 
  LUT3 #(
    .INIT(8'hD4)) 
    w_err__0_carry_i_1
       (.I0(\u_ras/w_dy [2]),
        .I1(w_err__0_carry_i_8_n_0),
        .I2(\u_ras/p_2_in [2]),
        .O(w_err__0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    w_err__0_carry_i_10
       (.I0(\u_ras/u_ras_line/r_x1 [0]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x0 [0]),
        .I3(w_err__0_carry_i_14_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(w_err__0_carry_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    w_err__0_carry_i_11
       (.I0(\u_ras/u_ras_line/r_x1 [3]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x0 [3]),
        .I3(w_err__0_carry_i_15_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(w_err__0_carry_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    w_err__0_carry_i_12
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_v0_x_reg_n_0_[2] ),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[2] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[2] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(w_err__0_carry_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    w_err__0_carry_i_13
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_v0_x_reg_n_0_[1] ),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[1] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[1] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(w_err__0_carry_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    w_err__0_carry_i_14
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_v0_x_reg_n_0_ ),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_ ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_ ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(w_err__0_carry_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDE488E4FADD5088)) 
    w_err__0_carry_i_15
       (.I0(_inferred__5_carry_i_14_n_0),
        .I1(\u_ras/u_ras_state/r_v0_x_reg_n_0_[3] ),
        .I2(\u_ras/u_ras_state/r_v1_x_reg_n_0_[3] ),
        .I3(\u_ras/u_ras_state/r_state [1]),
        .I4(\u_ras/u_ras_state/r_v2_x_reg_n_0_[3] ),
        .I5(\u_ras/u_ras_state/r_state [0]),
        .O(w_err__0_carry_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair0" *) 
  LUT3 #(
    .INIT(8'hD4)) 
    w_err__0_carry_i_2
       (.I0(\u_ras/w_dy [1]),
        .I1(w_err__0_carry_i_9_n_0),
        .I2(\u_ras/p_2_in [1]),
        .O(w_err__0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair8" *) 
  LUT3 #(
    .INIT(8'hD4)) 
    w_err__0_carry_i_3
       (.I0(\u_ras/w_dy [0]),
        .I1(w_err__0_carry_i_10_n_0),
        .I2(\u_ras/p_2_in [0]),
        .O(w_err__0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair2" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    w_err__0_carry_i_4
       (.I0(\u_ras/w_dy [3]),
        .I1(w_err__0_carry_i_11_n_0),
        .I2(\u_ras/p_2_in [3]),
        .I3(w_err__0_carry_i_1_n_0),
        .O(w_err__0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair1" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    w_err__0_carry_i_5
       (.I0(\u_ras/w_dy [2]),
        .I1(w_err__0_carry_i_8_n_0),
        .I2(\u_ras/p_2_in [2]),
        .I3(w_err__0_carry_i_2_n_0),
        .O(w_err__0_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair0" *) 
  LUT4 #(
    .INIT(16'h9669)) 
    w_err__0_carry_i_6
       (.I0(\u_ras/w_dy [1]),
        .I1(w_err__0_carry_i_9_n_0),
        .I2(\u_ras/p_2_in [1]),
        .I3(w_err__0_carry_i_3_n_0),
        .O(w_err__0_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair8" *) 
  LUT3 #(
    .INIT(8'h96)) 
    w_err__0_carry_i_7
       (.I0(\u_ras/w_dy [0]),
        .I1(w_err__0_carry_i_10_n_0),
        .I2(\u_ras/p_2_in [0]),
        .O(w_err__0_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    w_err__0_carry_i_8
       (.I0(\u_ras/u_ras_line/r_x1 [2]),
        .I1(_inferred__5_carry_i_9_n_0_repN),
        .I2(\u_ras/u_ras_line/r_x0 [2]),
        .I3(w_err__0_carry_i_12_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(w_err__0_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    w_err__0_carry_i_9
       (.I0(\u_ras/u_ras_line/r_x1 [1]),
        .I1(_inferred__5_carry_i_9_n_0),
        .I2(\u_ras/u_ras_line/r_x0 [1]),
        .I3(w_err__0_carry_i_13_n_0),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .O(w_err__0_carry_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_1
       (.I0(\u_geo/u_geo_matrix/w_m1_out [7]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [7]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [6]),
        .I3(\u_geo/u_geo_matrix/w_m0_out [6]),
        .O(w_mag_frac_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_10
       (.I0(\u_geo/w_vw_mvp [5]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [5]),
        .O(\u_geo/u_geo_clip/w_add_in_a [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_10__0
       (.I0(\u_geo/w_vw_mvp [13]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [13]),
        .O(\u_geo/u_geo_clip/w_add_in_a [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_11
       (.I0(\u_geo/w_vw_mvp [3]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [3]),
        .O(\u_geo/u_geo_clip/w_add_in_a [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_11__0
       (.I0(\u_geo/w_vw_mvp [11]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [11]),
        .O(\u_geo/u_geo_clip/w_add_in_a [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_12
       (.I0(\u_geo/w_vw_mvp [1]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [1]),
        .O(\u_geo/u_geo_clip/w_add_in_a [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_12__0
       (.I0(\u_geo/w_vw_mvp [9]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [9]),
        .O(\u_geo/u_geo_clip/w_add_in_a [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_13
       (.I0(\u_geo/w_vw_mvp [6]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [6]),
        .O(\u_geo/u_geo_clip/w_add_in_a [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_13__0
       (.I0(\u_geo/w_vw_mvp [14]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [14]),
        .O(\u_geo/u_geo_clip/w_add_in_a [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_14
       (.I0(\u_geo/w_vw_mvp [4]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [4]),
        .O(\u_geo/u_geo_clip/w_add_in_a [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_14__0
       (.I0(\u_geo/w_vw_mvp [12]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [12]),
        .O(\u_geo/u_geo_clip/w_add_in_a [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_15
       (.I0(\u_geo/w_vw_mvp [2]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [2]),
        .O(\u_geo/u_geo_clip/w_add_in_a [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_15__0
       (.I0(\u_geo/w_vw_mvp [10]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [10]),
        .O(\u_geo/u_geo_clip/w_add_in_a [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_16
       (.I0(\u_geo/w_vw_mvp [0]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [0]),
        .O(\u_geo/u_geo_clip/w_add_in_a [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_16__0
       (.I0(\u_geo/w_vw_mvp [8]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [8]),
        .O(\u_geo/u_geo_clip/w_add_in_a [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_1__0
       (.I0(\u_geo/u_geo_matrix/w_m1_out [15]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [15]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [14]),
        .I3(\u_geo/u_geo_matrix/w_m0_out [14]),
        .O(w_mag_frac_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_1__1
       (.I0(\u_geo/u_geo_matrix/w_m3_out [7]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [7]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [6]),
        .I3(\u_geo/u_geo_matrix/w_m2_out [6]),
        .O(w_mag_frac_carry_i_1__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_1__2
       (.I0(\u_geo/u_geo_matrix/w_m3_out [15]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [15]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [14]),
        .I3(\u_geo/u_geo_matrix/w_m2_out [14]),
        .O(w_mag_frac_carry_i_1__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_1__3
       (.I0(\u_geo/u_geo_matrix/w_add23_out [7]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [7]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [6]),
        .I3(\u_geo/u_geo_matrix/w_add01_out [6]),
        .O(w_mag_frac_carry_i_1__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_1__4
       (.I0(\u_geo/u_geo_matrix/w_add23_out [15]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [15]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [14]),
        .I3(\u_geo/u_geo_matrix/w_add01_out [14]),
        .O(w_mag_frac_carry_i_1__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h222222B2B2B222B2)) 
    w_mag_frac_carry_i_1__5
       (.I0(\r_f0[7]_i_2_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [7]),
        .I2(\r_f0[6]_i_2_n_0 ),
        .I3(\u_geo/w_vw_clip [6]),
        .I4(\u_geo/w_state_clip ),
        .I5(\u_geo/w_vw_mvp [6]),
        .O(w_mag_frac_carry_i_1__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h222222B2B2B222B2)) 
    w_mag_frac_carry_i_1__6
       (.I0(\r_f0[15]_i_3__2_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [15]),
        .I2(\r_f0[14]_i_2_n_0 ),
        .I3(\u_geo/w_vw_clip [14]),
        .I4(\u_geo/w_state_clip ),
        .I5(\u_geo/w_vw_mvp [14]),
        .O(w_mag_frac_carry_i_1__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_2
       (.I0(\u_geo/u_geo_matrix/w_m1_out [5]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [5]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [4]),
        .I3(\u_geo/u_geo_matrix/w_m0_out [4]),
        .O(w_mag_frac_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_2__0
       (.I0(\u_geo/u_geo_matrix/w_m1_out [13]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [13]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [12]),
        .I3(\u_geo/u_geo_matrix/w_m0_out [12]),
        .O(w_mag_frac_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_2__1
       (.I0(\u_geo/u_geo_matrix/w_m3_out [5]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [5]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [4]),
        .I3(\u_geo/u_geo_matrix/w_m2_out [4]),
        .O(w_mag_frac_carry_i_2__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_2__2
       (.I0(\u_geo/u_geo_matrix/w_m3_out [13]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [13]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [12]),
        .I3(\u_geo/u_geo_matrix/w_m2_out [12]),
        .O(w_mag_frac_carry_i_2__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_2__3
       (.I0(\u_geo/u_geo_matrix/w_add23_out [5]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [5]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [4]),
        .I3(\u_geo/u_geo_matrix/w_add01_out [4]),
        .O(w_mag_frac_carry_i_2__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_2__4
       (.I0(\u_geo/u_geo_matrix/w_add23_out [13]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [13]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [12]),
        .I3(\u_geo/u_geo_matrix/w_add01_out [12]),
        .O(w_mag_frac_carry_i_2__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h222222B2B2B222B2)) 
    w_mag_frac_carry_i_2__5
       (.I0(\r_f0[5]_i_2_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [5]),
        .I2(\r_f0[4]_i_2_n_0 ),
        .I3(\u_geo/w_vw_clip [4]),
        .I4(\u_geo/w_state_clip ),
        .I5(\u_geo/w_vw_mvp [4]),
        .O(w_mag_frac_carry_i_2__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h222222B2B2B222B2)) 
    w_mag_frac_carry_i_2__6
       (.I0(\r_f0[13]_i_2_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [13]),
        .I2(\r_f0[12]_i_2_n_0 ),
        .I3(\u_geo/w_vw_clip [12]),
        .I4(\u_geo/w_state_clip ),
        .I5(\u_geo/w_vw_mvp [12]),
        .O(w_mag_frac_carry_i_2__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_3
       (.I0(\u_geo/u_geo_matrix/w_m1_out [3]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [3]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [2]),
        .I3(\u_geo/u_geo_matrix/w_m0_out [2]),
        .O(w_mag_frac_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_3__0
       (.I0(\u_geo/u_geo_matrix/w_m1_out [11]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [11]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [10]),
        .I3(\u_geo/u_geo_matrix/w_m0_out [10]),
        .O(w_mag_frac_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_3__1
       (.I0(\u_geo/u_geo_matrix/w_m3_out [3]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [3]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [2]),
        .I3(\u_geo/u_geo_matrix/w_m2_out [2]),
        .O(w_mag_frac_carry_i_3__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_3__2
       (.I0(\u_geo/u_geo_matrix/w_m3_out [11]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [11]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [10]),
        .I3(\u_geo/u_geo_matrix/w_m2_out [10]),
        .O(w_mag_frac_carry_i_3__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_3__3
       (.I0(\u_geo/u_geo_matrix/w_add23_out [3]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [3]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [2]),
        .I3(\u_geo/u_geo_matrix/w_add01_out [2]),
        .O(w_mag_frac_carry_i_3__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_3__4
       (.I0(\u_geo/u_geo_matrix/w_add23_out [11]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [11]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [10]),
        .I3(\u_geo/u_geo_matrix/w_add01_out [10]),
        .O(w_mag_frac_carry_i_3__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h222222B2B2B222B2)) 
    w_mag_frac_carry_i_3__5
       (.I0(\r_f0[3]_i_2_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [3]),
        .I2(\r_f0[2]_i_2_n_0 ),
        .I3(\u_geo/w_vw_clip [2]),
        .I4(\u_geo/w_state_clip ),
        .I5(\u_geo/w_vw_mvp [2]),
        .O(w_mag_frac_carry_i_3__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h222222B2B2B222B2)) 
    w_mag_frac_carry_i_3__6
       (.I0(\r_f0[11]_i_2_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [11]),
        .I2(\r_f0[10]_i_2_n_0 ),
        .I3(\u_geo/w_vw_clip [10]),
        .I4(\u_geo/w_state_clip ),
        .I5(\u_geo/w_vw_mvp [10]),
        .O(w_mag_frac_carry_i_3__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_4
       (.I0(\u_geo/u_geo_matrix/w_m1_out [1]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [1]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [0]),
        .I3(\u_geo/u_geo_matrix/w_m0_out [0]),
        .O(w_mag_frac_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_4__0
       (.I0(\u_geo/u_geo_matrix/w_m1_out [9]),
        .I1(\u_geo/u_geo_matrix/w_m0_out [9]),
        .I2(\u_geo/u_geo_matrix/w_m1_out [8]),
        .I3(\u_geo/u_geo_matrix/w_m0_out [8]),
        .O(w_mag_frac_carry_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_4__1
       (.I0(\u_geo/u_geo_matrix/w_m3_out [1]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [1]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [0]),
        .I3(\u_geo/u_geo_matrix/w_m2_out [0]),
        .O(w_mag_frac_carry_i_4__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_4__2
       (.I0(\u_geo/u_geo_matrix/w_m3_out [9]),
        .I1(\u_geo/u_geo_matrix/w_m2_out [9]),
        .I2(\u_geo/u_geo_matrix/w_m3_out [8]),
        .I3(\u_geo/u_geo_matrix/w_m2_out [8]),
        .O(w_mag_frac_carry_i_4__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_4__3
       (.I0(\u_geo/u_geo_matrix/w_add23_out [1]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [1]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [0]),
        .I3(\u_geo/u_geo_matrix/w_add01_out [0]),
        .O(w_mag_frac_carry_i_4__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h22B2)) 
    w_mag_frac_carry_i_4__4
       (.I0(\u_geo/u_geo_matrix/w_add23_out [9]),
        .I1(\u_geo/u_geo_matrix/w_add01_out [9]),
        .I2(\u_geo/u_geo_matrix/w_add23_out [8]),
        .I3(\u_geo/u_geo_matrix/w_add01_out [8]),
        .O(w_mag_frac_carry_i_4__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h222222B2B2B222B2)) 
    w_mag_frac_carry_i_4__5
       (.I0(\r_f0[1]_i_2_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [1]),
        .I2(r_f0),
        .I3(\u_geo/w_vw_clip [0]),
        .I4(\u_geo/w_state_clip ),
        .I5(\u_geo/w_vw_mvp [0]),
        .O(w_mag_frac_carry_i_4__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h222222B2B2B222B2)) 
    w_mag_frac_carry_i_4__6
       (.I0(\r_f0[9]_i_2_n_0 ),
        .I1(\u_geo/u_geo_clip/w_add_in_a [9]),
        .I2(\r_f0[8]_i_2_n_0 ),
        .I3(\u_geo/w_vw_clip [8]),
        .I4(\u_geo/w_state_clip ),
        .I5(\u_geo/w_vw_mvp [8]),
        .O(w_mag_frac_carry_i_4__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_5
       (.I0(\u_geo/u_geo_matrix/w_m0_out [7]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [7]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [6]),
        .I3(\u_geo/u_geo_matrix/w_m1_out [6]),
        .O(w_mag_frac_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_5__0
       (.I0(\u_geo/u_geo_matrix/w_m0_out [15]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [15]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [14]),
        .I3(\u_geo/u_geo_matrix/w_m1_out [14]),
        .O(w_mag_frac_carry_i_5__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_5__1
       (.I0(\u_geo/u_geo_matrix/w_m2_out [7]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [7]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [6]),
        .I3(\u_geo/u_geo_matrix/w_m3_out [6]),
        .O(w_mag_frac_carry_i_5__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_5__2
       (.I0(\u_geo/u_geo_matrix/w_m2_out [15]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [15]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [14]),
        .I3(\u_geo/u_geo_matrix/w_m3_out [14]),
        .O(w_mag_frac_carry_i_5__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_5__3
       (.I0(\u_geo/u_geo_matrix/w_add01_out [7]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [7]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [6]),
        .I3(\u_geo/u_geo_matrix/w_add23_out [6]),
        .O(w_mag_frac_carry_i_5__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_5__4
       (.I0(\u_geo/u_geo_matrix/w_add01_out [15]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [15]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [14]),
        .I3(\u_geo/u_geo_matrix/w_add23_out [14]),
        .O(w_mag_frac_carry_i_5__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB84700000000B847)) 
    w_mag_frac_carry_i_5__5
       (.I0(\u_geo/w_vw_mvp [7]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [7]),
        .I3(\r_f0[7]_i_2_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [6]),
        .I5(\r_f0[6]_i_2_n_0 ),
        .O(w_mag_frac_carry_i_5__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB84700000000B847)) 
    w_mag_frac_carry_i_5__6
       (.I0(\u_geo/w_vw_mvp [15]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/u_geo_clip/r_vw_reg_n_0_ ),
        .I3(\r_f0[15]_i_3__2_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [14]),
        .I5(\r_f0[14]_i_2_n_0 ),
        .O(w_mag_frac_carry_i_5__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_6
       (.I0(\u_geo/u_geo_matrix/w_m0_out [5]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [5]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [4]),
        .I3(\u_geo/u_geo_matrix/w_m1_out [4]),
        .O(w_mag_frac_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_6__0
       (.I0(\u_geo/u_geo_matrix/w_m0_out [13]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [13]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [12]),
        .I3(\u_geo/u_geo_matrix/w_m1_out [12]),
        .O(w_mag_frac_carry_i_6__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_6__1
       (.I0(\u_geo/u_geo_matrix/w_m2_out [5]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [5]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [4]),
        .I3(\u_geo/u_geo_matrix/w_m3_out [4]),
        .O(w_mag_frac_carry_i_6__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_6__2
       (.I0(\u_geo/u_geo_matrix/w_m2_out [13]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [13]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [12]),
        .I3(\u_geo/u_geo_matrix/w_m3_out [12]),
        .O(w_mag_frac_carry_i_6__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_6__3
       (.I0(\u_geo/u_geo_matrix/w_add01_out [5]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [5]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [4]),
        .I3(\u_geo/u_geo_matrix/w_add23_out [4]),
        .O(w_mag_frac_carry_i_6__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_6__4
       (.I0(\u_geo/u_geo_matrix/w_add01_out [13]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [13]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [12]),
        .I3(\u_geo/u_geo_matrix/w_add23_out [12]),
        .O(w_mag_frac_carry_i_6__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB84700000000B847)) 
    w_mag_frac_carry_i_6__5
       (.I0(\u_geo/w_vw_mvp [5]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [5]),
        .I3(\r_f0[5]_i_2_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [4]),
        .I5(\r_f0[4]_i_2_n_0 ),
        .O(w_mag_frac_carry_i_6__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB84700000000B847)) 
    w_mag_frac_carry_i_6__6
       (.I0(\u_geo/w_vw_mvp [13]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [13]),
        .I3(\r_f0[13]_i_2_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [12]),
        .I5(\r_f0[12]_i_2_n_0 ),
        .O(w_mag_frac_carry_i_6__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_7
       (.I0(\u_geo/u_geo_matrix/w_m0_out [3]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [3]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [2]),
        .I3(\u_geo/u_geo_matrix/w_m1_out [2]),
        .O(w_mag_frac_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_7__0
       (.I0(\u_geo/u_geo_matrix/w_m0_out [11]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [11]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [10]),
        .I3(\u_geo/u_geo_matrix/w_m1_out [10]),
        .O(w_mag_frac_carry_i_7__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_7__1
       (.I0(\u_geo/u_geo_matrix/w_m2_out [3]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [3]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [2]),
        .I3(\u_geo/u_geo_matrix/w_m3_out [2]),
        .O(w_mag_frac_carry_i_7__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_7__2
       (.I0(\u_geo/u_geo_matrix/w_m2_out [11]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [11]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [10]),
        .I3(\u_geo/u_geo_matrix/w_m3_out [10]),
        .O(w_mag_frac_carry_i_7__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_7__3
       (.I0(\u_geo/u_geo_matrix/w_add01_out [3]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [3]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [2]),
        .I3(\u_geo/u_geo_matrix/w_add23_out [2]),
        .O(w_mag_frac_carry_i_7__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_7__4
       (.I0(\u_geo/u_geo_matrix/w_add01_out [11]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [11]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [10]),
        .I3(\u_geo/u_geo_matrix/w_add23_out [10]),
        .O(w_mag_frac_carry_i_7__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB84700000000B847)) 
    w_mag_frac_carry_i_7__5
       (.I0(\u_geo/w_vw_mvp [3]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [3]),
        .I3(\r_f0[3]_i_2_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [2]),
        .I5(\r_f0[2]_i_2_n_0 ),
        .O(w_mag_frac_carry_i_7__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB84700000000B847)) 
    w_mag_frac_carry_i_7__6
       (.I0(\u_geo/w_vw_mvp [11]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [11]),
        .I3(\r_f0[11]_i_2_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [10]),
        .I5(\r_f0[10]_i_2_n_0 ),
        .O(w_mag_frac_carry_i_7__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_8
       (.I0(\u_geo/u_geo_matrix/w_m0_out [1]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [1]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [0]),
        .I3(\u_geo/u_geo_matrix/w_m1_out [0]),
        .O(w_mag_frac_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_8__0
       (.I0(\u_geo/u_geo_matrix/w_m0_out [9]),
        .I1(\u_geo/u_geo_matrix/w_m1_out [9]),
        .I2(\u_geo/u_geo_matrix/w_m0_out [8]),
        .I3(\u_geo/u_geo_matrix/w_m1_out [8]),
        .O(w_mag_frac_carry_i_8__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_8__1
       (.I0(\u_geo/u_geo_matrix/w_m2_out [1]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [1]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [0]),
        .I3(\u_geo/u_geo_matrix/w_m3_out [0]),
        .O(w_mag_frac_carry_i_8__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_8__2
       (.I0(\u_geo/u_geo_matrix/w_m2_out [9]),
        .I1(\u_geo/u_geo_matrix/w_m3_out [9]),
        .I2(\u_geo/u_geo_matrix/w_m2_out [8]),
        .I3(\u_geo/u_geo_matrix/w_m3_out [8]),
        .O(w_mag_frac_carry_i_8__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_8__3
       (.I0(\u_geo/u_geo_matrix/w_add01_out [1]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [1]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [0]),
        .I3(\u_geo/u_geo_matrix/w_add23_out [0]),
        .O(w_mag_frac_carry_i_8__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_mag_frac_carry_i_8__4
       (.I0(\u_geo/u_geo_matrix/w_add01_out [9]),
        .I1(\u_geo/u_geo_matrix/w_add23_out [9]),
        .I2(\u_geo/u_geo_matrix/w_add01_out [8]),
        .I3(\u_geo/u_geo_matrix/w_add23_out [8]),
        .O(w_mag_frac_carry_i_8__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB84700000000B847)) 
    w_mag_frac_carry_i_8__5
       (.I0(\u_geo/w_vw_mvp [1]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [1]),
        .I3(\r_f0[1]_i_2_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [0]),
        .I5(r_f0),
        .O(w_mag_frac_carry_i_8__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB84700000000B847)) 
    w_mag_frac_carry_i_8__6
       (.I0(\u_geo/w_vw_mvp [9]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [9]),
        .I3(\r_f0[9]_i_2_n_0 ),
        .I4(\u_geo/u_geo_clip/w_add_in_a [8]),
        .I5(\r_f0[8]_i_2_n_0 ),
        .O(w_mag_frac_carry_i_8__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_9
       (.I0(\u_geo/w_vw_mvp [7]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/w_vw_clip [7]),
        .O(\u_geo/u_geo_clip/w_add_in_a [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    w_mag_frac_carry_i_9__0
       (.I0(\u_geo/w_vw_mvp [15]),
        .I1(\u_geo/w_state_clip ),
        .I2(\u_geo/u_geo_clip/r_vw_reg_n_0_ ),
        .O(\u_geo/u_geo_clip/w_add_in_a [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    w_reject0_carry__0_i_1
       (.I0(w_scr_h_m1[10]),
        .I1(\u_ras/r_y [10]),
        .I2(w_scr_h_m1[11]),
        .O(w_reject0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    w_reject0_carry__0_i_2
       (.I0(\u_ras/r_y [8]),
        .I1(w_scr_h_m1[8]),
        .I2(w_scr_h_m1[9]),
        .I3(\u_ras/r_y [9]),
        .O(w_reject0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    w_reject0_carry__0_i_3
       (.I0(w_scr_h_m1[14]),
        .I1(w_scr_h_m1[15]),
        .O(w_reject0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    w_reject0_carry__0_i_4
       (.I0(w_scr_h_m1[12]),
        .I1(w_scr_h_m1[13]),
        .O(w_reject0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h09)) 
    w_reject0_carry__0_i_5
       (.I0(\u_ras/r_y [10]),
        .I1(w_scr_h_m1[10]),
        .I2(w_scr_h_m1[11]),
        .O(w_reject0_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_reject0_carry__0_i_6
       (.I0(\u_ras/r_y [8]),
        .I1(w_scr_h_m1[8]),
        .I2(\u_ras/r_y [9]),
        .I3(w_scr_h_m1[9]),
        .O(w_reject0_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    w_reject0_carry_i_1
       (.I0(\u_ras/r_y [6]),
        .I1(w_scr_h_m1[6]),
        .I2(w_scr_h_m1[7]),
        .I3(\u_ras/r_y [7]),
        .O(w_reject0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    w_reject0_carry_i_2
       (.I0(\u_ras/r_y [4]),
        .I1(w_scr_h_m1[4]),
        .I2(w_scr_h_m1[5]),
        .I3(\u_ras/r_y [5]),
        .O(w_reject0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    w_reject0_carry_i_3
       (.I0(\u_ras/r_y [2]),
        .I1(w_scr_h_m1[2]),
        .I2(w_scr_h_m1[3]),
        .I3(\u_ras/r_y [3]),
        .O(w_reject0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    w_reject0_carry_i_4
       (.I0(\u_ras/r_y [0]),
        .I1(w_scr_h_m1[0]),
        .I2(w_scr_h_m1[1]),
        .I3(\u_ras/r_y [1]),
        .O(w_reject0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_reject0_carry_i_5
       (.I0(\u_ras/r_y [6]),
        .I1(w_scr_h_m1[6]),
        .I2(\u_ras/r_y [7]),
        .I3(w_scr_h_m1[7]),
        .O(w_reject0_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_reject0_carry_i_6
       (.I0(\u_ras/r_y [4]),
        .I1(w_scr_h_m1[4]),
        .I2(\u_ras/r_y [5]),
        .I3(w_scr_h_m1[5]),
        .O(w_reject0_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_reject0_carry_i_7
       (.I0(\u_ras/r_y [2]),
        .I1(w_scr_h_m1[2]),
        .I2(\u_ras/r_y [3]),
        .I3(w_scr_h_m1[3]),
        .O(w_reject0_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_reject0_carry_i_8
       (.I0(\u_ras/r_y [0]),
        .I1(w_scr_h_m1[0]),
        .I2(\u_ras/r_y [1]),
        .I3(w_scr_h_m1[1]),
        .O(w_reject0_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    w_reject1_carry__0_i_1
       (.I0(w_scr_w_m1[10]),
        .I1(\u_ras/u_ras_line/r_x_reg_n_0_[10] ),
        .I2(w_scr_w_m1[11]),
        .O(w_reject1_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    w_reject1_carry__0_i_2
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[8] ),
        .I1(w_scr_w_m1[8]),
        .I2(w_scr_w_m1[9]),
        .I3(\u_ras/u_ras_line/r_x_reg_n_0_[9] ),
        .O(w_reject1_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    w_reject1_carry__0_i_3
       (.I0(w_scr_w_m1[14]),
        .I1(w_scr_w_m1[15]),
        .O(w_reject1_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    w_reject1_carry__0_i_4
       (.I0(w_scr_w_m1[12]),
        .I1(w_scr_w_m1[13]),
        .O(w_reject1_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h09)) 
    w_reject1_carry__0_i_5
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[10] ),
        .I1(w_scr_w_m1[10]),
        .I2(w_scr_w_m1[11]),
        .O(w_reject1_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_reject1_carry__0_i_6
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[8] ),
        .I1(w_scr_w_m1[8]),
        .I2(\u_ras/u_ras_line/r_x_reg_n_0_[9] ),
        .I3(w_scr_w_m1[9]),
        .O(w_reject1_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    w_reject1_carry_i_1
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[6] ),
        .I1(w_scr_w_m1[6]),
        .I2(w_scr_w_m1[7]),
        .I3(\u_ras/u_ras_line/r_x_reg_n_0_[7] ),
        .O(w_reject1_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    w_reject1_carry_i_2
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[4] ),
        .I1(w_scr_w_m1[4]),
        .I2(w_scr_w_m1[5]),
        .I3(\u_ras/u_ras_line/r_x_reg_n_0_[5] ),
        .O(w_reject1_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    w_reject1_carry_i_3
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[2] ),
        .I1(w_scr_w_m1[2]),
        .I2(w_scr_w_m1[3]),
        .I3(\u_ras/u_ras_line/r_x_reg_n_0_[3] ),
        .O(w_reject1_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    w_reject1_carry_i_4
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_ ),
        .I1(w_scr_w_m1[0]),
        .I2(w_scr_w_m1[1]),
        .I3(\u_ras/u_ras_line/r_x_reg_n_0_[1] ),
        .O(w_reject1_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_reject1_carry_i_5
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[6] ),
        .I1(w_scr_w_m1[6]),
        .I2(\u_ras/u_ras_line/r_x_reg_n_0_[7] ),
        .I3(w_scr_w_m1[7]),
        .O(w_reject1_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_reject1_carry_i_6
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[4] ),
        .I1(w_scr_w_m1[4]),
        .I2(\u_ras/u_ras_line/r_x_reg_n_0_[5] ),
        .I3(w_scr_w_m1[5]),
        .O(w_reject1_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_reject1_carry_i_7
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_[2] ),
        .I1(w_scr_w_m1[2]),
        .I2(\u_ras/u_ras_line/r_x_reg_n_0_[3] ),
        .I3(w_scr_w_m1[3]),
        .O(w_reject1_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    w_reject1_carry_i_8
       (.I0(\u_ras/u_ras_line/r_x_reg_n_0_ ),
        .I1(w_scr_w_m1[0]),
        .I2(\u_ras/u_ras_line/r_x_reg_n_0_[1] ),
        .I3(w_scr_w_m1[1]),
        .O(w_reject1_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    w_rom_correct_i_1
       (.I0(g0_b8_n_0),
        .I1(\u_geo/w_vw_clip [14]),
        .O(w_rom_correct_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F2F22FF02020022)) 
    w_sx_flag1_carry__0_i_1
       (.I0(\u_ras/w_x1 [10]),
        .I1(\u_ras/w_x0 [10]),
        .I2(\u_ras/u_ras_line/r_x0 [11]),
        .I3(\u_ras/w_v0_x [11]),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .I5(\u_ras/w_x1 [11]),
        .O(w_sx_flag1_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry__0_i_10
       (.I0(\u_ras/u_ras_line/r_x1 [9]),
        .I1(\u_ras/w_v1_x [9]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    w_sx_flag1_carry__0_i_11
       (.I0(\u_ras/w_v0_x [11]),
        .I1(\u_ras/u_ras_line/r_x0 [11]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/w_v1_x [11]),
        .I4(\u_ras/u_ras_line/r_x1 [11]),
        .O(w_sx_flag1_carry__0_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    w_sx_flag1_carry__0_i_12
       (.I0(\u_ras/w_v0_x [9]),
        .I1(\u_ras/u_ras_line/r_x0 [9]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/w_v1_x [9]),
        .I4(\u_ras/u_ras_line/r_x1 [9]),
        .O(w_sx_flag1_carry__0_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h028AFFFF0000028A)) 
    w_sx_flag1_carry__0_i_2
       (.I0(\u_ras/w_x1 [8]),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(\u_ras/w_v0_x [8]),
        .I3(\u_ras/u_ras_line/r_x0 [8]),
        .I4(\u_ras/w_x0 [9]),
        .I5(\u_ras/w_x1 [9]),
        .O(w_sx_flag1_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC5CA35300000000)) 
    w_sx_flag1_carry__0_i_3
       (.I0(\u_ras/u_ras_line/r_x1 [10]),
        .I1(\u_ras/w_v1_x [10]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_x0 [10]),
        .I4(\u_ras/w_v0_x [10]),
        .I5(w_sx_flag1_carry__0_i_11_n_0),
        .O(w_sx_flag1_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC5CA35300000000)) 
    w_sx_flag1_carry__0_i_4
       (.I0(\u_ras/u_ras_line/r_x1 [8]),
        .I1(\u_ras/w_v1_x [8]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_x0 [8]),
        .I4(\u_ras/w_v0_x [8]),
        .I5(w_sx_flag1_carry__0_i_12_n_0),
        .O(w_sx_flag1_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry__0_i_5
       (.I0(\u_ras/u_ras_line/r_x1 [10]),
        .I1(\u_ras/w_v1_x [10]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry__0_i_6
       (.I0(\u_ras/u_ras_line/r_x0 [10]),
        .I1(\u_ras/w_v0_x[10]_repN ),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x0 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry__0_i_7
       (.I0(\u_ras/u_ras_line/r_x1 [11]),
        .I1(\u_ras/w_v1_x [11]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry__0_i_8
       (.I0(\u_ras/u_ras_line/r_x1 [8]),
        .I1(\u_ras/w_v1_x [8]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry__0_i_9
       (.I0(\u_ras/u_ras_line/r_x0 [9]),
        .I1(\u_ras/w_v0_x [9]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x0 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h028AFFFF0000028A)) 
    w_sx_flag1_carry_i_1
       (.I0(\u_ras/w_x1 [6]),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(\u_ras/w_v0_x [6]),
        .I3(\u_ras/u_ras_line/r_x0 [6]),
        .I4(\u_ras/w_x0 [7]),
        .I5(\u_ras/w_x1 [7]),
        .O(w_sx_flag1_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry_i_10
       (.I0(\u_ras/u_ras_line/r_x0 [7]),
        .I1(\u_ras/w_v0_x [7]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x0 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry_i_11
       (.I0(\u_ras/u_ras_line/r_x1 [7]),
        .I1(\u_ras/w_v1_x [7]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry_i_12
       (.I0(\u_ras/u_ras_line/r_x1 [4]),
        .I1(\u_ras/w_v1_x [4]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry_i_13
       (.I0(\u_ras/u_ras_line/r_x0 [5]),
        .I1(\u_ras/w_v0_x [5]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x0 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry_i_14
       (.I0(\u_ras/u_ras_line/r_x1 [5]),
        .I1(\u_ras/w_v1_x [5]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry_i_15
       (.I0(\u_ras/u_ras_line/r_x1 [2]),
        .I1(\u_ras/w_v1_x [2]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry_i_16
       (.I0(\u_ras/u_ras_line/r_x0 [3]),
        .I1(\u_ras/w_v0_x [3]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry_i_17
       (.I0(\u_ras/u_ras_line/r_x1 [3]),
        .I1(\u_ras/w_v1_x [3]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry_i_18
       (.I0(\u_ras/u_ras_line/r_x1 [0]),
        .I1(\u_ras/w_v1_x [0]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x1 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry_i_19
       (.I0(\u_ras/u_ras_line/r_x0 [1]),
        .I1(\u_ras/w_v0_x [1]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h028AFFFF0000028A)) 
    w_sx_flag1_carry_i_2
       (.I0(\u_ras/w_x1 [4]),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(\u_ras/w_v0_x [4]),
        .I3(\u_ras/u_ras_line/r_x0 [4]),
        .I4(\u_ras/w_x0 [5]),
        .I5(\u_ras/w_x1 [5]),
        .O(w_sx_flag1_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry_i_20
       (.I0(\u_ras/u_ras_line/r_x1 [1]),
        .I1(\u_ras/w_v1_x [1]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    w_sx_flag1_carry_i_21
       (.I0(\u_ras/w_v0_x [7]),
        .I1(\u_ras/u_ras_line/r_x0 [7]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/w_v1_x [7]),
        .I4(\u_ras/u_ras_line/r_x1 [7]),
        .O(w_sx_flag1_carry_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    w_sx_flag1_carry_i_22
       (.I0(\u_ras/w_v0_x [5]),
        .I1(\u_ras/u_ras_line/r_x0 [5]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/w_v1_x [5]),
        .I4(\u_ras/u_ras_line/r_x1 [5]),
        .O(w_sx_flag1_carry_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    w_sx_flag1_carry_i_23
       (.I0(\u_ras/w_v0_x [3]),
        .I1(\u_ras/u_ras_line/r_x0 [3]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/w_v1_x [3]),
        .I4(\u_ras/u_ras_line/r_x1 [3]),
        .O(w_sx_flag1_carry_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    w_sx_flag1_carry_i_24
       (.I0(\u_ras/w_v0_x [1]),
        .I1(\u_ras/u_ras_line/r_x0 [1]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/w_v1_x [1]),
        .I4(\u_ras/u_ras_line/r_x1 [1]),
        .O(w_sx_flag1_carry_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h028AFFFF0000028A)) 
    w_sx_flag1_carry_i_3
       (.I0(\u_ras/w_x1 [2]),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(\u_ras/w_v0_x [2]),
        .I3(\u_ras/u_ras_line/r_x0 [2]),
        .I4(\u_ras/w_x0 [3]),
        .I5(\u_ras/w_x1 [3]),
        .O(w_sx_flag1_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h028AFFFF0000028A)) 
    w_sx_flag1_carry_i_4
       (.I0(\u_ras/w_x1 [0]),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(\u_ras/w_v0_x [0]),
        .I3(\u_ras/u_ras_line/r_x0 [0]),
        .I4(\u_ras/w_x0 [1]),
        .I5(\u_ras/w_x1 [1]),
        .O(w_sx_flag1_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC5CA35300000000)) 
    w_sx_flag1_carry_i_5
       (.I0(\u_ras/u_ras_line/r_x1 [6]),
        .I1(\u_ras/w_v1_x [6]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_x0 [6]),
        .I4(\u_ras/w_v0_x [6]),
        .I5(w_sx_flag1_carry_i_21_n_0),
        .O(w_sx_flag1_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC5CA35300000000)) 
    w_sx_flag1_carry_i_6
       (.I0(\u_ras/u_ras_line/r_x1 [4]),
        .I1(\u_ras/w_v1_x [4]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_x0 [4]),
        .I4(\u_ras/w_v0_x [4]),
        .I5(w_sx_flag1_carry_i_22_n_0),
        .O(w_sx_flag1_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC5CA35300000000)) 
    w_sx_flag1_carry_i_7
       (.I0(\u_ras/u_ras_line/r_x1 [2]),
        .I1(\u_ras/w_v1_x [2]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_x0 [2]),
        .I4(\u_ras/w_v0_x [2]),
        .I5(w_sx_flag1_carry_i_23_n_0),
        .O(w_sx_flag1_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC5CA35300000000)) 
    w_sx_flag1_carry_i_8
       (.I0(\u_ras/u_ras_line/r_x1 [0]),
        .I1(\u_ras/w_v1_x [0]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_x0 [0]),
        .I4(\u_ras/w_v0_x [0]),
        .I5(w_sx_flag1_carry_i_24_n_0),
        .O(w_sx_flag1_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sx_flag1_carry_i_9
       (.I0(\u_ras/u_ras_line/r_x1 [6]),
        .I1(\u_ras/w_v1_x [6]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_x1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2F2F22FF02020022)) 
    w_sy_flag1_carry__0_i_1
       (.I0(\u_ras/w_y1 [10]),
        .I1(\u_ras/w_y0 [10]),
        .I2(\u_ras/u_ras_line/r_y0 [11]),
        .I3(\u_ras/w_v0_y [11]),
        .I4(w_sy_flag1_carry_i_10_n_0),
        .I5(\u_ras/w_y1 [11]),
        .O(w_sy_flag1_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry__0_i_10
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[9] ),
        .I1(\u_ras/w_v1_y [9]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    w_sy_flag1_carry__0_i_11
       (.I0(\u_ras/w_v0_y [11]),
        .I1(\u_ras/u_ras_line/r_y0 [11]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/w_v1_y [11]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[11] ),
        .O(w_sy_flag1_carry__0_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    w_sy_flag1_carry__0_i_12
       (.I0(\u_ras/w_v0_y [9]),
        .I1(\u_ras/u_ras_line/r_y0 [9]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/w_v1_y [9]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[9] ),
        .O(w_sy_flag1_carry__0_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h028AFFFF0000028A)) 
    w_sy_flag1_carry__0_i_2
       (.I0(\u_ras/w_y1 [8]),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(\u_ras/w_v0_y [8]),
        .I3(\u_ras/u_ras_line/r_y0 [8]),
        .I4(\u_ras/w_y0 [9]),
        .I5(\u_ras/w_y1 [9]),
        .O(w_sy_flag1_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC5CA35300000000)) 
    w_sy_flag1_carry__0_i_3
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[10] ),
        .I1(\u_ras/w_v1_y [10]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [10]),
        .I4(\u_ras/w_v0_y [10]),
        .I5(w_sy_flag1_carry__0_i_11_n_0),
        .O(w_sy_flag1_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC5CA35300000000)) 
    w_sy_flag1_carry__0_i_4
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[8] ),
        .I1(\u_ras/w_v1_y [8]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [8]),
        .I4(\u_ras/w_v0_y [8]),
        .I5(w_sy_flag1_carry__0_i_12_n_0),
        .O(w_sy_flag1_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry__0_i_5
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[10] ),
        .I1(\u_ras/w_v1_y [10]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry__0_i_6
       (.I0(\u_ras/u_ras_line/r_y0 [10]),
        .I1(\u_ras/w_v0_y[10]_repN ),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y0 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry__0_i_7
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[11] ),
        .I1(\u_ras/w_v1_y [11]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry__0_i_8
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[8] ),
        .I1(\u_ras/w_v1_y [8]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry__0_i_9
       (.I0(\u_ras/u_ras_line/r_y0 [9]),
        .I1(\u_ras/w_v0_y [9]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y0 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h028AFFFF0000028A)) 
    w_sy_flag1_carry_i_1
       (.I0(\u_ras/w_y1[6]_repN ),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(\u_ras/w_v0_y [6]),
        .I3(\u_ras/u_ras_line/r_y0 [6]),
        .I4(\u_ras/w_y0 [7]),
        .I5(\u_ras/w_y1 [7]),
        .O(w_sy_flag1_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    w_sy_flag1_carry_i_10
       (.I0(\u_ras/u_ras_line/r_state_reg_n_0_[1] ),
        .I1(\u_ras/u_ras_line/r_state_reg_n_0_ ),
        .O(w_sy_flag1_carry_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_11
       (.I0(\u_ras/u_ras_line/r_y0 [7]),
        .I1(\u_ras/w_v0_y [7]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y0 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_12
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[7] ),
        .I1(\u_ras/w_v1_y [7]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_13
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[4] ),
        .I1(\u_ras/w_v1_y [4]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_14
       (.I0(\u_ras/u_ras_line/r_y0 [5]),
        .I1(\u_ras/w_v0_y [5]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y0 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_15
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[5] ),
        .I1(\u_ras/w_v1_y [5]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_16
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[2] ),
        .I1(\u_ras/w_v1_y [2]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_17
       (.I0(\u_ras/u_ras_line/r_y0 [3]),
        .I1(\u_ras/w_v0_y [3]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_18
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[3] ),
        .I1(\u_ras/w_v1_y [3]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_19
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_ ),
        .I1(\u_ras/w_v1_y [0]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h028AFFFF0000028A)) 
    w_sy_flag1_carry_i_2
       (.I0(\u_ras/w_y1 [4]),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(\u_ras/w_v0_y [4]),
        .I3(\u_ras/u_ras_line/r_y0 [4]),
        .I4(\u_ras/w_y0 [5]),
        .I5(\u_ras/w_y1 [5]),
        .O(w_sy_flag1_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_20
       (.I0(\u_ras/u_ras_line/r_y0 [1]),
        .I1(\u_ras/w_v0_y [1]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_21
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[1] ),
        .I1(\u_ras/w_v1_y [1]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "w_sy_flag1_carry_i_21" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_21_replica
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[1] ),
        .I1(\u_ras/w_v1_y [1]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1[1]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    w_sy_flag1_carry_i_22
       (.I0(\u_ras/w_v0_y [7]),
        .I1(\u_ras/u_ras_line/r_y0 [7]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/w_v1_y [7]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[7] ),
        .O(w_sy_flag1_carry_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    w_sy_flag1_carry_i_23
       (.I0(\u_ras/w_v0_y [5]),
        .I1(\u_ras/u_ras_line/r_y0 [5]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/w_v1_y [5]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[5] ),
        .O(w_sy_flag1_carry_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    w_sy_flag1_carry_i_24
       (.I0(\u_ras/w_v0_y [3]),
        .I1(\u_ras/u_ras_line/r_y0 [3]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/w_v1_y [3]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[3] ),
        .O(w_sy_flag1_carry_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    w_sy_flag1_carry_i_25
       (.I0(\u_ras/w_v0_y [1]),
        .I1(\u_ras/u_ras_line/r_y0 [1]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/w_v1_y [1]),
        .I4(\u_ras/u_ras_line/r_y1_reg_n_0_[1] ),
        .O(w_sy_flag1_carry_i_25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h028AFFFF0000028A)) 
    w_sy_flag1_carry_i_3
       (.I0(\u_ras/w_y1 [2]),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(\u_ras/w_v0_y [2]),
        .I3(\u_ras/u_ras_line/r_y0 [2]),
        .I4(\u_ras/w_y0 [3]),
        .I5(\u_ras/w_y1 [3]),
        .O(w_sy_flag1_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h028AFFFF0000028A)) 
    w_sy_flag1_carry_i_4
       (.I0(\u_ras/w_y1 [0]),
        .I1(w_sy_flag1_carry_i_10_n_0),
        .I2(\u_ras/w_v0_y [0]),
        .I3(\u_ras/u_ras_line/r_y0 [0]),
        .I4(\u_ras/w_y0 [1]),
        .I5(\u_ras/w_y1[1]_repN ),
        .O(w_sy_flag1_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC5CA35300000000)) 
    w_sy_flag1_carry_i_5
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[6] ),
        .I1(\u_ras/w_v1_y [6]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [6]),
        .I4(\u_ras/w_v0_y [6]),
        .I5(w_sy_flag1_carry_i_22_n_0),
        .O(w_sy_flag1_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC5CA35300000000)) 
    w_sy_flag1_carry_i_6
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[4] ),
        .I1(\u_ras/w_v1_y [4]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [4]),
        .I4(\u_ras/w_v0_y [4]),
        .I5(w_sy_flag1_carry_i_23_n_0),
        .O(w_sy_flag1_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC5CA35300000000)) 
    w_sy_flag1_carry_i_7
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[2] ),
        .I1(\u_ras/w_v1_y [2]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [2]),
        .I4(\u_ras/w_v0_y [2]),
        .I5(w_sy_flag1_carry_i_24_n_0),
        .O(w_sy_flag1_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAC5CA35300000000)) 
    w_sy_flag1_carry_i_8
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_ ),
        .I1(\u_ras/w_v1_y [0]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .I3(\u_ras/u_ras_line/r_y0 [0]),
        .I4(\u_ras/w_v0_y [0]),
        .I5(w_sy_flag1_carry_i_25_n_0),
        .O(w_sy_flag1_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_9
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[6] ),
        .I1(\u_ras/w_v1_y [6]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "w_sy_flag1_carry_i_9" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    w_sy_flag1_carry_i_9_replica
       (.I0(\u_ras/u_ras_line/r_y1_reg_n_0_[6] ),
        .I1(\u_ras/w_v1_y [6]),
        .I2(w_sy_flag1_carry_i_10_n_0),
        .O(\u_ras/w_y1[6]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_y0_carry_i_1
       (.I0(w_scr_h_m1[11]),
        .I1(\u_ras/w_y ),
        .O(w_y0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_y0_carry_i_1__0
       (.I0(w_scr_h_m1[7]),
        .I1(\u_ras/r_y [7]),
        .O(w_y0_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_y0_carry_i_1__1
       (.I0(w_scr_h_m1[3]),
        .I1(\u_ras/r_y [3]),
        .O(w_y0_carry_i_1__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_y0_carry_i_2
       (.I0(w_scr_h_m1[10]),
        .I1(\u_ras/r_y [10]),
        .O(w_y0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_y0_carry_i_2__0
       (.I0(w_scr_h_m1[6]),
        .I1(\u_ras/r_y [6]),
        .O(w_y0_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_y0_carry_i_2__1
       (.I0(w_scr_h_m1[2]),
        .I1(\u_ras/r_y [2]),
        .O(w_y0_carry_i_2__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_y0_carry_i_3
       (.I0(w_scr_h_m1[9]),
        .I1(\u_ras/r_y [9]),
        .O(w_y0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_y0_carry_i_3__0
       (.I0(w_scr_h_m1[5]),
        .I1(\u_ras/r_y [5]),
        .O(w_y0_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_y0_carry_i_3__1
       (.I0(w_scr_h_m1[1]),
        .I1(\u_ras/r_y [1]),
        .O(w_y0_carry_i_3__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_y0_carry_i_4
       (.I0(w_scr_h_m1[8]),
        .I1(\u_ras/r_y [8]),
        .O(w_y0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_y0_carry_i_4__0
       (.I0(w_scr_h_m1[4]),
        .I1(\u_ras/r_y [4]),
        .O(w_y0_carry_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    w_y0_carry_i_4__1
       (.I0(w_scr_h_m1[0]),
        .I1(\u_ras/r_y [0]),
        .O(w_y0_carry_i_4__1_n_0));
endmodule
