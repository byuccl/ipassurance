// This holds the blackbox module definitions for the dfadd

module dfadd
	(
input clk,
input reset,
input start,
output finish,
input waitrequest,
output [31:0] return_val);
endmodule // dfadd