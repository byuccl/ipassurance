module basicrsa
   (indata,
    inExp,
    inMod,
    cypher,
    clk,
    ds,
    reset,
    backdoor,
    ready);
  output backdoor;
  input [31:0]indata;
  input [31:0]inExp;
  input [31:0]inMod;
  output [31:0]cypher;
  input clk;
  input ds;
  input reset;
  output ready;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire count;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire count_reg_n_0_;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \count_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]cypher;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[31]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[31]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[31]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[31]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cypher[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire done_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ds;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire first_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire first_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]inExp;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]inMod;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]indata;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [33:0]mcreg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[0]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[10]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[11]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[12]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[12]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[12]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[12]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[12]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[12]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[13]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[14]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[15]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[16]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[16]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[16]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[16]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[16]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[16]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[17]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[18]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[19]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[1]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[20]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[20]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[20]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[20]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[20]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[20]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[20]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[21]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[22]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[23]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[24]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[24]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[24]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[24]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[24]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[24]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[24]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[25]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[26]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[27]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[28]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[28]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[28]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[28]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[28]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[28]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[28]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[29]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[2]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[30]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[31]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[32]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[32]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[32]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[32]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[32]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[32]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[32]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[32]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[32]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[32]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[33]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[33]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[33]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[33]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[3]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[4]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[4]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[4]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[4]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[4]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[5]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[6]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[7]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[8]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[8]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[8]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[8]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[8]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[9]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]mcreg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[12]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[12]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[12]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[12]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[12]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[12]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[12]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[16]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[16]_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[16]_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[16]_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[16]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[16]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[16]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[16]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[16]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[16]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[16]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[20]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[20]_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[20]_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[20]_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[20]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[20]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[20]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[20]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[20]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[20]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[20]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[24]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[24]_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[24]_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[24]_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[24]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[24]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[24]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[24]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[24]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[24]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[24]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[28]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[28]_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[28]_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[28]_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[28]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[28]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[28]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[28]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[28]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[28]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[28]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[32]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[32]_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[32]_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[32]_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[32]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[32]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[32]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[32]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[32]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[32]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[32]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[32]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[33]_i_2__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[33]_i_2__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[33]_i_2__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[33]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[33]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[33]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[33]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[4]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[4]_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[4]_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[4]_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[4]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[4]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[4]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[4]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[4]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[4]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[4]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[8]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[8]_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[8]_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[8]_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[8]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[8]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[8]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[8]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[8]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[8]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mcreg_reg[8]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [32:0]minusOp;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [33:0]minusOp0_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__0_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__0_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__0_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__0_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__1_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__1_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__1_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__1_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__2_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__2_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__2_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__2_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__2_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__2_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__2_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__2_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__3_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__3_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__3_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__3_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__3_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__3_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__3_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__3_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__4_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__4_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__4_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__4_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__4_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__4_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__4_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__4_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__5_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__5_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__5_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__5_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__5_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__5_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__5_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__5_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__6_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__6_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__6_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__6_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__6_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__6_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__6_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__6_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__7_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__7_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__7_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__7_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__0_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__0_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__0_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__0_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__1_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__1_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__1_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__1_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__2_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__2_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__2_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__2_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__2_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__2_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__2_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__2_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__3_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__3_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__3_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__3_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__3_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__3_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__3_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__3_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__4_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__4_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__4_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__4_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__4_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__4_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__4_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__4_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__5_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__5_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__5_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__5_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__5_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__5_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__5_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__5_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__6_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__6_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__6_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__6_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__6_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__6_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__6_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__6_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__7_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__7_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__7_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry__7_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__1_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__5_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__5_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__5_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__5_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__6_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__6_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__6_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__6_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__7_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__7_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__7_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry__7_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__0_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__7_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry__7_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/minusOp_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/mpreg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__7_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry__7_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/plusOp_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modmultiply/prodreg0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]modreg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:1]modreg1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modreg2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modreg[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mcreg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__5_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__5_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__5_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__5_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__6_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__6_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__6_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__6_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__7_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__7_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__7_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry__7_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__0_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__5_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__5_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__5_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__5_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__6_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__6_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__6_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__6_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__7_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__7_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__7_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry__7_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/minusOp_inferred__1_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg1_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/modreg2_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/mpreg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__5_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__5_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__5_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__5_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__6_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__6_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__6_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__6_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__7_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__7_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__7_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry__7_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/plusOp_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \modsqr/prodreg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire mpreg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[10]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[11]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[12]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[13]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[14]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[15]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[16]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[17]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[18]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[19]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[1]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[20]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[21]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[22]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[23]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[24]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[25]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[26]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[27]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[28]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[29]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[2]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[30]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_10__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_11__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_4__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_5__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_6__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_7__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_8__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_9__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[31]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[3]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[4]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[5]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[6]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[7]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[8]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[9]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \mpreg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multgo_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multgo_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multgo_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multgo_reg_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multrdy;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__0_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__0_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__0_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__0_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__1_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__1_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__1_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__1_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__2_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__2_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__2_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__2_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__2_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__2_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__2_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__2_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__3_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__3_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__3_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__3_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__3_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__3_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__3_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__3_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__4_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__4_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__4_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__4_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__4_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__4_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__4_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__4_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__5_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__5_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__5_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__5_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__5_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__5_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__5_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__5_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__6_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__6_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__6_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__6_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__6_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__6_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__6_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__6_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__7_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__7_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__7_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry__7_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [33:0]prodreg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [33:0]prodreg1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[32]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[32]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[33]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[33]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[33]_i_3__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[33]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \prodreg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ready;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire reset;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]root;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \root[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sqrin;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sqrin_reg_n_0_;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sqrin_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sqrrdy;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]tempin;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \tempin[9]_i_1_n_0 ;

  assign backdoor =  sqrrdy ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[0]_i_1 
       (.I0(inExp[1]),
        .I1(ready),
        .I2(\count_reg_n_0_[1] ),
        .O(count));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[10]_i_1 
       (.I0(inExp[11]),
        .I1(ready),
        .I2(\count_reg_n_0_[11] ),
        .O(\count[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[11]_i_1 
       (.I0(inExp[12]),
        .I1(ready),
        .I2(\count_reg_n_0_[12] ),
        .O(\count[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[12]_i_1 
       (.I0(inExp[13]),
        .I1(ready),
        .I2(\count_reg_n_0_[13] ),
        .O(\count[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[13]_i_1 
       (.I0(inExp[14]),
        .I1(ready),
        .I2(\count_reg_n_0_[14] ),
        .O(\count[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[14]_i_1 
       (.I0(inExp[15]),
        .I1(ready),
        .I2(\count_reg_n_0_[15] ),
        .O(\count[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[15]_i_1 
       (.I0(inExp[16]),
        .I1(ready),
        .I2(\count_reg_n_0_[16] ),
        .O(\count[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[16]_i_1 
       (.I0(inExp[17]),
        .I1(ready),
        .I2(\count_reg_n_0_[17] ),
        .O(\count[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[17]_i_1 
       (.I0(inExp[18]),
        .I1(ready),
        .I2(\count_reg_n_0_[18] ),
        .O(\count[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[18]_i_1 
       (.I0(inExp[19]),
        .I1(ready),
        .I2(\count_reg_n_0_[19] ),
        .O(\count[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[19]_i_1 
       (.I0(inExp[20]),
        .I1(ready),
        .I2(\count_reg_n_0_[20] ),
        .O(\count[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[1]_i_1 
       (.I0(inExp[2]),
        .I1(ready),
        .I2(\count_reg_n_0_[2] ),
        .O(\count[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[20]_i_1 
       (.I0(inExp[21]),
        .I1(ready),
        .I2(\count_reg_n_0_[21] ),
        .O(\count[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[21]_i_1 
       (.I0(inExp[22]),
        .I1(ready),
        .I2(\count_reg_n_0_[22] ),
        .O(\count[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[22]_i_1 
       (.I0(inExp[23]),
        .I1(ready),
        .I2(\count_reg_n_0_[23] ),
        .O(\count[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[23]_i_1 
       (.I0(inExp[24]),
        .I1(ready),
        .I2(\count_reg_n_0_[24] ),
        .O(\count[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[24]_i_1 
       (.I0(inExp[25]),
        .I1(ready),
        .I2(\count_reg_n_0_[25] ),
        .O(\count[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[25]_i_1 
       (.I0(inExp[26]),
        .I1(ready),
        .I2(\count_reg_n_0_[26] ),
        .O(\count[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[26]_i_1 
       (.I0(inExp[27]),
        .I1(ready),
        .I2(\count_reg_n_0_[27] ),
        .O(\count[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[27]_i_1 
       (.I0(inExp[28]),
        .I1(ready),
        .I2(\count_reg_n_0_[28] ),
        .O(\count[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[28]_i_1 
       (.I0(inExp[29]),
        .I1(ready),
        .I2(\count_reg_n_0_[29] ),
        .O(\count[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[29]_i_1 
       (.I0(inExp[30]),
        .I1(ready),
        .I2(\count_reg_n_0_[30] ),
        .O(\count[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[2]_i_1 
       (.I0(inExp[3]),
        .I1(ready),
        .I2(\count_reg_n_0_[3] ),
        .O(\count[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFF8F88888888)) 
    \count[30]_i_1 
       (.I0(ds),
        .I1(ready),
        .I2(\cypher[31]_i_3_n_0 ),
        .I3(\cypher[31]_i_4_n_0 ),
        .I4(\cypher[31]_i_5_n_0 ),
        .I5(\cypher[31]_i_6_n_0 ),
        .O(\count[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \count[30]_i_2 
       (.I0(ready),
        .I1(inExp[31]),
        .O(\count[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[3]_i_1 
       (.I0(inExp[4]),
        .I1(ready),
        .I2(\count_reg_n_0_[4] ),
        .O(\count[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[4]_i_1 
       (.I0(inExp[5]),
        .I1(ready),
        .I2(\count_reg_n_0_[5] ),
        .O(\count[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[5]_i_1 
       (.I0(inExp[6]),
        .I1(ready),
        .I2(\count_reg_n_0_[6] ),
        .O(\count[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[6]_i_1 
       (.I0(inExp[7]),
        .I1(ready),
        .I2(\count_reg_n_0_[7] ),
        .O(\count[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[7]_i_1 
       (.I0(inExp[8]),
        .I1(ready),
        .I2(\count_reg_n_0_[8] ),
        .O(\count[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[8]_i_1 
       (.I0(inExp[9]),
        .I1(ready),
        .I2(\count_reg_n_0_[9] ),
        .O(\count[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \count[9]_i_1 
       (.I0(inExp[10]),
        .I1(ready),
        .I2(\count_reg_n_0_[10] ),
        .O(\count[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[0] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(count),
        .Q(count_reg_n_0_));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[10] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[10]_i_1_n_0 ),
        .Q(\count_reg_n_0_[10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[11] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[11]_i_1_n_0 ),
        .Q(\count_reg_n_0_[11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[12] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[12]_i_1_n_0 ),
        .Q(\count_reg_n_0_[12] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[13] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[13]_i_1_n_0 ),
        .Q(\count_reg_n_0_[13] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[14] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[14]_i_1_n_0 ),
        .Q(\count_reg_n_0_[14] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[15] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[15]_i_1_n_0 ),
        .Q(\count_reg_n_0_[15] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[16] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[16]_i_1_n_0 ),
        .Q(\count_reg_n_0_[16] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[17] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[17]_i_1_n_0 ),
        .Q(\count_reg_n_0_[17] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[18] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[18]_i_1_n_0 ),
        .Q(\count_reg_n_0_[18] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[19] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[19]_i_1_n_0 ),
        .Q(\count_reg_n_0_[19] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[1] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[1]_i_1_n_0 ),
        .Q(\count_reg_n_0_[1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[20] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[20]_i_1_n_0 ),
        .Q(\count_reg_n_0_[20] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[21] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[21]_i_1_n_0 ),
        .Q(\count_reg_n_0_[21] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[22] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[22]_i_1_n_0 ),
        .Q(\count_reg_n_0_[22] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[23] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[23]_i_1_n_0 ),
        .Q(\count_reg_n_0_[23] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[24] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[24]_i_1_n_0 ),
        .Q(\count_reg_n_0_[24] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[25] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[25]_i_1_n_0 ),
        .Q(\count_reg_n_0_[25] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[26] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[26]_i_1_n_0 ),
        .Q(\count_reg_n_0_[26] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[27] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[27]_i_1_n_0 ),
        .Q(\count_reg_n_0_[27] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[28] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[28]_i_1_n_0 ),
        .Q(\count_reg_n_0_[28] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[29] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[29]_i_1_n_0 ),
        .Q(\count_reg_n_0_[29] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[2] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[2]_i_1_n_0 ),
        .Q(\count_reg_n_0_[2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[30] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[30]_i_2_n_0 ),
        .Q(\count_reg_n_0_[30] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[3] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[3]_i_1_n_0 ),
        .Q(\count_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[4] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[4]_i_1_n_0 ),
        .Q(\count_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[5] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[5]_i_1_n_0 ),
        .Q(\count_reg_n_0_[5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[6] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[6]_i_1_n_0 ),
        .Q(\count_reg_n_0_[6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[7] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[7]_i_1_n_0 ),
        .Q(\count_reg_n_0_[7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[8] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[8]_i_1_n_0 ),
        .Q(\count_reg_n_0_[8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \count_reg[9] 
       (.C(clk),
        .CE(\count[30]_i_1_n_0 ),
        .CLR(reset),
        .D(\count[9]_i_1_n_0 ),
        .Q(\count_reg_n_0_[9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[0]_i_1 
       (.I0(prodreg1[0]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry_n_7 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[0]),
        .O(\cypher[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[10]_i_1 
       (.I0(prodreg1[10]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__1_n_5 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[10]),
        .O(\cypher[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[11]_i_1 
       (.I0(prodreg1[11]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__1_n_4 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[11]),
        .O(\cypher[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[12]_i_1 
       (.I0(prodreg1[12]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__2_n_7 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[12]),
        .O(\cypher[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[13]_i_1 
       (.I0(prodreg1[13]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__2_n_6 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[13]),
        .O(\cypher[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[14]_i_1 
       (.I0(prodreg1[14]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__2_n_5 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[14]),
        .O(\cypher[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[15]_i_1 
       (.I0(prodreg1[15]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__2_n_4 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[15]),
        .O(\cypher[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[16]_i_1 
       (.I0(prodreg1[16]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__3_n_7 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[16]),
        .O(\cypher[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[17]_i_1 
       (.I0(prodreg1[17]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__3_n_6 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[17]),
        .O(\cypher[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[18]_i_1 
       (.I0(prodreg1[18]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__3_n_5 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[18]),
        .O(\cypher[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[19]_i_1 
       (.I0(prodreg1[19]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__3_n_4 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[19]),
        .O(\cypher[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[1]_i_1 
       (.I0(prodreg1[1]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry_n_6 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[1]),
        .O(\cypher[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[20]_i_1 
       (.I0(prodreg1[20]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__4_n_7 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[20]),
        .O(\cypher[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[21]_i_1 
       (.I0(prodreg1[21]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__4_n_6 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[21]),
        .O(\cypher[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[22]_i_1 
       (.I0(prodreg1[22]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__4_n_5 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[22]),
        .O(\cypher[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[23]_i_1 
       (.I0(prodreg1[23]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__4_n_4 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[23]),
        .O(\cypher[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[24]_i_1 
       (.I0(prodreg1[24]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__5_n_7 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[24]),
        .O(\cypher[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[25]_i_1 
       (.I0(prodreg1[25]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__5_n_6 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[25]),
        .O(\cypher[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[26]_i_1 
       (.I0(prodreg1[26]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__5_n_5 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[26]),
        .O(\cypher[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[27]_i_1 
       (.I0(prodreg1[27]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__5_n_4 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[27]),
        .O(\cypher[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[28]_i_1 
       (.I0(prodreg1[28]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__6_n_7 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[28]),
        .O(\cypher[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[29]_i_1 
       (.I0(prodreg1[29]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__6_n_6 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[29]),
        .O(\cypher[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[2]_i_1 
       (.I0(prodreg1[2]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry_n_5 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[2]),
        .O(\cypher[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[30]_i_1 
       (.I0(prodreg1[30]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__6_n_5 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[30]),
        .O(\cypher[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \cypher[31]_i_1 
       (.I0(reset),
        .I1(\cypher[31]_i_3_n_0 ),
        .I2(\cypher[31]_i_4_n_0 ),
        .I3(\cypher[31]_i_5_n_0 ),
        .I4(\cypher[31]_i_6_n_0 ),
        .O(\cypher[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \cypher[31]_i_10 
       (.I0(\count_reg_n_0_[27] ),
        .I1(\count_reg_n_0_[17] ),
        .I2(\count_reg_n_0_[19] ),
        .I3(\count_reg_n_0_[15] ),
        .O(\cypher[31]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \cypher[31]_i_11 
       (.I0(\count_reg_n_0_[26] ),
        .I1(\count_reg_n_0_[10] ),
        .I2(\count_reg_n_0_[25] ),
        .I3(\count_reg_n_0_[18] ),
        .O(\cypher[31]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[31]_i_2 
       (.I0(prodreg1[31]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__6_n_4 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[31]),
        .O(\cypher[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \cypher[31]_i_3 
       (.I0(\cypher[31]_i_7_n_0 ),
        .I1(\cypher[31]_i_8_n_0 ),
        .I2(\cypher[31]_i_9_n_0 ),
        .I3(\count_reg_n_0_[13] ),
        .I4(\count_reg_n_0_[24] ),
        .I5(\count_reg_n_0_[8] ),
        .O(\cypher[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \cypher[31]_i_4 
       (.I0(\count_reg_n_0_[11] ),
        .I1(\count_reg_n_0_[21] ),
        .I2(\count_reg_n_0_[9] ),
        .I3(\count_reg_n_0_[22] ),
        .I4(\cypher[31]_i_10_n_0 ),
        .O(\cypher[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \cypher[31]_i_5 
       (.I0(\count_reg_n_0_[5] ),
        .I1(\count_reg_n_0_[6] ),
        .I2(\count_reg_n_0_[4] ),
        .I3(\count_reg_n_0_[7] ),
        .I4(\cypher[31]_i_11_n_0 ),
        .O(\cypher[31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \cypher[31]_i_6 
       (.I0(multgo_reg_n_0),
        .I1(multrdy),
        .I2(sqrrdy),
        .I3(ready),
        .O(\cypher[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \cypher[31]_i_7 
       (.I0(\count_reg_n_0_[20] ),
        .I1(\count_reg_n_0_[3] ),
        .I2(\count_reg_n_0_[28] ),
        .I3(\count_reg_n_0_[14] ),
        .O(\cypher[31]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \cypher[31]_i_8 
       (.I0(\count_reg_n_0_[30] ),
        .I1(\count_reg_n_0_[23] ),
        .I2(\count_reg_n_0_[29] ),
        .I3(\count_reg_n_0_[2] ),
        .O(\cypher[31]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \cypher[31]_i_9 
       (.I0(\count_reg_n_0_[16] ),
        .I1(\count_reg_n_0_[1] ),
        .I2(\count_reg_n_0_[12] ),
        .I3(count_reg_n_0_),
        .O(\cypher[31]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[3]_i_1 
       (.I0(prodreg1[3]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry_n_4 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[3]),
        .O(\cypher[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[4]_i_1 
       (.I0(prodreg1[4]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__0_n_7 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[4]),
        .O(\cypher[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[5]_i_1 
       (.I0(prodreg1[5]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__0_n_6 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[5]),
        .O(\cypher[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[6]_i_1 
       (.I0(prodreg1[6]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__0_n_5 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[6]),
        .O(\cypher[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[7]_i_1 
       (.I0(prodreg1[7]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__0_n_4 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[7]),
        .O(\cypher[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[8]_i_1 
       (.I0(prodreg1[8]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__1_n_7 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[8]),
        .O(\cypher[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cypher[9]_i_1 
       (.I0(prodreg1[9]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__1_n_6 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[9]),
        .O(\cypher[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[0] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[0]_i_1_n_0 ),
        .Q(cypher[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[10] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[10]_i_1_n_0 ),
        .Q(cypher[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[11] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[11]_i_1_n_0 ),
        .Q(cypher[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[12] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[12]_i_1_n_0 ),
        .Q(cypher[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[13] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[13]_i_1_n_0 ),
        .Q(cypher[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[14] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[14]_i_1_n_0 ),
        .Q(cypher[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[15] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[15]_i_1_n_0 ),
        .Q(cypher[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[16] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[16]_i_1_n_0 ),
        .Q(cypher[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[17] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[17]_i_1_n_0 ),
        .Q(cypher[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[18] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[18]_i_1_n_0 ),
        .Q(cypher[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[19] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[19]_i_1_n_0 ),
        .Q(cypher[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[1] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[1]_i_1_n_0 ),
        .Q(cypher[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[20] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[20]_i_1_n_0 ),
        .Q(cypher[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[21] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[21]_i_1_n_0 ),
        .Q(cypher[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[22] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[22]_i_1_n_0 ),
        .Q(cypher[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[23] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[23]_i_1_n_0 ),
        .Q(cypher[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[24] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[24]_i_1_n_0 ),
        .Q(cypher[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[25] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[25]_i_1_n_0 ),
        .Q(cypher[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[26] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[26]_i_1_n_0 ),
        .Q(cypher[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[27] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[27]_i_1_n_0 ),
        .Q(cypher[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[28] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[28]_i_1_n_0 ),
        .Q(cypher[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[29] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[29]_i_1_n_0 ),
        .Q(cypher[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[2] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[2]_i_1_n_0 ),
        .Q(cypher[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[30] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[30]_i_1_n_0 ),
        .Q(cypher[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[31] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[31]_i_2_n_0 ),
        .Q(cypher[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[3] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[3]_i_1_n_0 ),
        .Q(cypher[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[4] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[4]_i_1_n_0 ),
        .Q(cypher[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[5] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[5]_i_1_n_0 ),
        .Q(cypher[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[6] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[6]_i_1_n_0 ),
        .Q(cypher[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[7] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[7]_i_1_n_0 ),
        .Q(cypher[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[8] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[8]_i_1_n_0 ),
        .Q(cypher[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \cypher_reg[9] 
       (.C(clk),
        .CE(\cypher[31]_i_1_n_0 ),
        .D(\cypher[9]_i_1_n_0 ),
        .Q(cypher[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCCCCFC44444444)) 
    done_i_1
       (.I0(ds),
        .I1(ready),
        .I2(\cypher[31]_i_3_n_0 ),
        .I3(\cypher[31]_i_4_n_0 ),
        .I4(\cypher[31]_i_5_n_0 ),
        .I5(\cypher[31]_i_6_n_0 ),
        .O(done_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    done_reg
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(done_i_1_n_0),
        .PRE(reset),
        .Q(ready));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT3 #(
    .INIT(8'h35)) 
    first_i_1
       (.I0(\mpreg[31]_i_3_n_0 ),
        .I1(multgo_reg_n_0),
        .I2(multrdy),
        .O(first_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT3 #(
    .INIT(8'h1D)) 
    first_i_1__0
       (.I0(\mpreg[31]_i_3__0_n_0 ),
        .I1(sqrrdy),
        .I2(multgo_reg_n_0),
        .O(first_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \mcreg[0]_i_1 
       (.I0(sqrrdy),
        .I1(root[0]),
        .O(\mcreg[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \mcreg[0]_i_1__0 
       (.I0(multrdy),
        .I1(tempin[0]),
        .O(\mcreg[0]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[10]_i_1 
       (.I0(root[10]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[9] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[12]_i_2_n_6 ),
        .O(\mcreg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[10]_i_1__0 
       (.I0(tempin[10]),
        .I1(multrdy),
        .I2(mcreg[9]),
        .I3(minusOp[32]),
        .I4(minusOp[9]),
        .O(\mcreg[10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[11]_i_1 
       (.I0(root[11]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[10] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[12]_i_2_n_5 ),
        .O(\mcreg[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[11]_i_1__0 
       (.I0(tempin[11]),
        .I1(multrdy),
        .I2(mcreg[10]),
        .I3(minusOp[32]),
        .I4(minusOp[10]),
        .O(\mcreg[11]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[12]_i_1 
       (.I0(root[12]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[11] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[12]_i_2_n_4 ),
        .O(\mcreg[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[12]_i_1__0 
       (.I0(tempin[12]),
        .I1(multrdy),
        .I2(mcreg[11]),
        .I3(minusOp[32]),
        .I4(minusOp[11]),
        .O(\mcreg[12]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[12]_i_3 
       (.I0(\modsqr/mcreg_reg_n_0_[11] ),
        .I1(\modsqr/modreg1_reg_n_0_[11] ),
        .O(\mcreg[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[12]_i_3__0 
       (.I0(mcreg[11]),
        .I1(modreg1[11]),
        .O(\mcreg[12]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[12]_i_4 
       (.I0(\modsqr/mcreg_reg_n_0_[10] ),
        .I1(\modsqr/modreg1_reg_n_0_ ),
        .O(\mcreg[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[12]_i_4__0 
       (.I0(mcreg[10]),
        .I1(modreg1[10]),
        .O(\mcreg[12]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[12]_i_5 
       (.I0(\modsqr/mcreg_reg_n_0_[9] ),
        .I1(\modsqr/modreg1_reg_n_0_[9] ),
        .O(\mcreg[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[12]_i_5__0 
       (.I0(mcreg[9]),
        .I1(modreg1[9]),
        .O(\mcreg[12]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[12]_i_6 
       (.I0(\modsqr/mcreg_reg_n_0_[8] ),
        .I1(\modsqr/modreg1_reg_n_0_[8] ),
        .O(\mcreg[12]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[12]_i_6__0 
       (.I0(mcreg[8]),
        .I1(modreg1[8]),
        .O(\mcreg[12]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[13]_i_1 
       (.I0(root[13]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[12] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[16]_i_2_n_7 ),
        .O(\mcreg[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[13]_i_1__0 
       (.I0(tempin[13]),
        .I1(multrdy),
        .I2(mcreg[12]),
        .I3(minusOp[32]),
        .I4(minusOp[12]),
        .O(\mcreg[13]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[14]_i_1 
       (.I0(root[14]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[13] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[16]_i_2_n_6 ),
        .O(\mcreg[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[14]_i_1__0 
       (.I0(tempin[14]),
        .I1(multrdy),
        .I2(mcreg[13]),
        .I3(minusOp[32]),
        .I4(minusOp[13]),
        .O(\mcreg[14]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[15]_i_1 
       (.I0(root[15]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[14] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[16]_i_2_n_5 ),
        .O(\mcreg[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[15]_i_1__0 
       (.I0(tempin[15]),
        .I1(multrdy),
        .I2(mcreg[14]),
        .I3(minusOp[32]),
        .I4(minusOp[14]),
        .O(\mcreg[15]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[16]_i_1 
       (.I0(root[16]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[15] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[16]_i_2_n_4 ),
        .O(\mcreg[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[16]_i_1__0 
       (.I0(tempin[16]),
        .I1(multrdy),
        .I2(mcreg[15]),
        .I3(minusOp[32]),
        .I4(minusOp[15]),
        .O(\mcreg[16]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[16]_i_3 
       (.I0(\modsqr/mcreg_reg_n_0_[15] ),
        .I1(\modsqr/modreg1_reg_n_0_[15] ),
        .O(\mcreg[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[16]_i_3__0 
       (.I0(mcreg[15]),
        .I1(modreg1[15]),
        .O(\mcreg[16]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[16]_i_4 
       (.I0(\modsqr/mcreg_reg_n_0_[14] ),
        .I1(\modsqr/modreg1_reg_n_0_[14] ),
        .O(\mcreg[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[16]_i_4__0 
       (.I0(mcreg[14]),
        .I1(modreg1[14]),
        .O(\mcreg[16]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[16]_i_5 
       (.I0(\modsqr/mcreg_reg_n_0_[13] ),
        .I1(\modsqr/modreg1_reg_n_0_[13] ),
        .O(\mcreg[16]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[16]_i_5__0 
       (.I0(mcreg[13]),
        .I1(modreg1[13]),
        .O(\mcreg[16]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[16]_i_6 
       (.I0(\modsqr/mcreg_reg_n_0_[12] ),
        .I1(\modsqr/modreg1_reg_n_0_[12] ),
        .O(\mcreg[16]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[16]_i_6__0 
       (.I0(mcreg[12]),
        .I1(modreg1[12]),
        .O(\mcreg[16]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[17]_i_1 
       (.I0(root[17]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[16] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[20]_i_2_n_7 ),
        .O(\mcreg[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[17]_i_1__0 
       (.I0(tempin[17]),
        .I1(multrdy),
        .I2(mcreg[16]),
        .I3(minusOp[32]),
        .I4(minusOp[16]),
        .O(\mcreg[17]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[18]_i_1 
       (.I0(root[18]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[17] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[20]_i_2_n_6 ),
        .O(\mcreg[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[18]_i_1__0 
       (.I0(tempin[18]),
        .I1(multrdy),
        .I2(mcreg[17]),
        .I3(minusOp[32]),
        .I4(minusOp[17]),
        .O(\mcreg[18]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[19]_i_1 
       (.I0(root[19]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[18] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[20]_i_2_n_5 ),
        .O(\mcreg[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[19]_i_1__0 
       (.I0(tempin[19]),
        .I1(multrdy),
        .I2(mcreg[18]),
        .I3(minusOp[32]),
        .I4(minusOp[18]),
        .O(\mcreg[19]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[1]_i_1 
       (.I0(root[1]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_ ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[4]_i_2_n_7 ),
        .O(\mcreg[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[1]_i_1__0 
       (.I0(tempin[1]),
        .I1(multrdy),
        .I2(mcreg[0]),
        .I3(minusOp[32]),
        .I4(minusOp[0]),
        .O(\mcreg[1]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[20]_i_1 
       (.I0(root[20]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[19] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[20]_i_2_n_4 ),
        .O(\mcreg[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[20]_i_1__0 
       (.I0(tempin[20]),
        .I1(multrdy),
        .I2(mcreg[19]),
        .I3(minusOp[32]),
        .I4(minusOp[19]),
        .O(\mcreg[20]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[20]_i_3 
       (.I0(\modsqr/mcreg_reg_n_0_[19] ),
        .I1(\modsqr/modreg1_reg_n_0_[19] ),
        .O(\mcreg[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[20]_i_3__0 
       (.I0(mcreg[19]),
        .I1(modreg1[19]),
        .O(\mcreg[20]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[20]_i_4 
       (.I0(\modsqr/mcreg_reg_n_0_[18] ),
        .I1(\modsqr/modreg1_reg_n_0_[18] ),
        .O(\mcreg[20]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[20]_i_4__0 
       (.I0(mcreg[18]),
        .I1(modreg1[18]),
        .O(\mcreg[20]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[20]_i_5 
       (.I0(\modsqr/mcreg_reg_n_0_[17] ),
        .I1(\modsqr/modreg1_reg_n_0_[17] ),
        .O(\mcreg[20]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[20]_i_5__0 
       (.I0(mcreg[17]),
        .I1(modreg1[17]),
        .O(\mcreg[20]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[20]_i_6 
       (.I0(\modsqr/mcreg_reg_n_0_[16] ),
        .I1(\modsqr/modreg1_reg_n_0_[16] ),
        .O(\mcreg[20]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[20]_i_6__0 
       (.I0(mcreg[16]),
        .I1(modreg1[16]),
        .O(\mcreg[20]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[21]_i_1 
       (.I0(root[21]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[20] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[24]_i_2_n_7 ),
        .O(\mcreg[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[21]_i_1__0 
       (.I0(tempin[21]),
        .I1(multrdy),
        .I2(mcreg[20]),
        .I3(minusOp[32]),
        .I4(minusOp[20]),
        .O(\mcreg[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[22]_i_1 
       (.I0(root[22]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[21] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[24]_i_2_n_6 ),
        .O(\mcreg[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[22]_i_1__0 
       (.I0(tempin[22]),
        .I1(multrdy),
        .I2(mcreg[21]),
        .I3(minusOp[32]),
        .I4(minusOp[21]),
        .O(\mcreg[22]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[23]_i_1 
       (.I0(root[23]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[22] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[24]_i_2_n_5 ),
        .O(\mcreg[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[23]_i_1__0 
       (.I0(tempin[23]),
        .I1(multrdy),
        .I2(mcreg[22]),
        .I3(minusOp[32]),
        .I4(minusOp[22]),
        .O(\mcreg[23]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[24]_i_1 
       (.I0(root[24]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[23] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[24]_i_2_n_4 ),
        .O(\mcreg[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[24]_i_1__0 
       (.I0(tempin[24]),
        .I1(multrdy),
        .I2(mcreg[23]),
        .I3(minusOp[32]),
        .I4(minusOp[23]),
        .O(\mcreg[24]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[24]_i_3 
       (.I0(\modsqr/mcreg_reg_n_0_[23] ),
        .I1(\modsqr/modreg1_reg_n_0_[23] ),
        .O(\mcreg[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[24]_i_3__0 
       (.I0(mcreg[23]),
        .I1(modreg1[23]),
        .O(\mcreg[24]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[24]_i_4 
       (.I0(\modsqr/mcreg_reg_n_0_[22] ),
        .I1(\modsqr/modreg1_reg_n_0_[22] ),
        .O(\mcreg[24]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[24]_i_4__0 
       (.I0(mcreg[22]),
        .I1(modreg1[22]),
        .O(\mcreg[24]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[24]_i_5 
       (.I0(\modsqr/mcreg_reg_n_0_[21] ),
        .I1(\modsqr/modreg1_reg_n_0_[21] ),
        .O(\mcreg[24]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[24]_i_5__0 
       (.I0(mcreg[21]),
        .I1(modreg1[21]),
        .O(\mcreg[24]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[24]_i_6 
       (.I0(\modsqr/mcreg_reg_n_0_[20] ),
        .I1(\modsqr/modreg1_reg_n_0_[20] ),
        .O(\mcreg[24]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[24]_i_6__0 
       (.I0(mcreg[20]),
        .I1(modreg1[20]),
        .O(\mcreg[24]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[25]_i_1 
       (.I0(root[25]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[24] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[28]_i_2_n_7 ),
        .O(\mcreg[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[25]_i_1__0 
       (.I0(tempin[25]),
        .I1(multrdy),
        .I2(mcreg[24]),
        .I3(minusOp[32]),
        .I4(minusOp[24]),
        .O(\mcreg[25]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[26]_i_1 
       (.I0(root[26]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[25] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[28]_i_2_n_6 ),
        .O(\mcreg[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[26]_i_1__0 
       (.I0(tempin[26]),
        .I1(multrdy),
        .I2(mcreg[25]),
        .I3(minusOp[32]),
        .I4(minusOp[25]),
        .O(\mcreg[26]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[27]_i_1 
       (.I0(root[27]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[26] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[28]_i_2_n_5 ),
        .O(\mcreg[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[27]_i_1__0 
       (.I0(tempin[27]),
        .I1(multrdy),
        .I2(mcreg[26]),
        .I3(minusOp[32]),
        .I4(minusOp[26]),
        .O(\mcreg[27]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[28]_i_1 
       (.I0(root[28]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[27] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[28]_i_2_n_4 ),
        .O(\mcreg[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[28]_i_1__0 
       (.I0(tempin[28]),
        .I1(multrdy),
        .I2(mcreg[27]),
        .I3(minusOp[32]),
        .I4(minusOp[27]),
        .O(\mcreg[28]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[28]_i_3 
       (.I0(\modsqr/mcreg_reg_n_0_[27] ),
        .I1(\modsqr/modreg1_reg_n_0_[27] ),
        .O(\mcreg[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[28]_i_3__0 
       (.I0(mcreg[27]),
        .I1(modreg1[27]),
        .O(\mcreg[28]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[28]_i_4 
       (.I0(\modsqr/mcreg_reg_n_0_[26] ),
        .I1(\modsqr/modreg1_reg_n_0_[26] ),
        .O(\mcreg[28]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[28]_i_4__0 
       (.I0(mcreg[26]),
        .I1(modreg1[26]),
        .O(\mcreg[28]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[28]_i_5 
       (.I0(\modsqr/mcreg_reg_n_0_[25] ),
        .I1(\modsqr/modreg1_reg_n_0_[25] ),
        .O(\mcreg[28]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[28]_i_5__0 
       (.I0(mcreg[25]),
        .I1(modreg1[25]),
        .O(\mcreg[28]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[28]_i_6 
       (.I0(\modsqr/mcreg_reg_n_0_[24] ),
        .I1(\modsqr/modreg1_reg_n_0_[24] ),
        .O(\mcreg[28]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[28]_i_6__0 
       (.I0(mcreg[24]),
        .I1(modreg1[24]),
        .O(\mcreg[28]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[29]_i_1 
       (.I0(root[29]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[28] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[32]_i_2_n_7 ),
        .O(\mcreg[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[29]_i_1__0 
       (.I0(tempin[29]),
        .I1(multrdy),
        .I2(mcreg[28]),
        .I3(minusOp[32]),
        .I4(minusOp[28]),
        .O(\mcreg[29]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[2]_i_1 
       (.I0(root[2]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[1] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[4]_i_2_n_6 ),
        .O(\mcreg[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[2]_i_1__0 
       (.I0(tempin[2]),
        .I1(multrdy),
        .I2(mcreg[1]),
        .I3(minusOp[32]),
        .I4(minusOp[1]),
        .O(\mcreg[2]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[30]_i_1 
       (.I0(root[30]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[29] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[32]_i_2_n_6 ),
        .O(\mcreg[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[30]_i_1__0 
       (.I0(tempin[30]),
        .I1(multrdy),
        .I2(mcreg[29]),
        .I3(minusOp[32]),
        .I4(minusOp[29]),
        .O(\mcreg[30]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[31]_i_1 
       (.I0(root[31]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[30] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[32]_i_2_n_5 ),
        .O(\mcreg[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[31]_i_1__0 
       (.I0(tempin[31]),
        .I1(multrdy),
        .I2(mcreg[30]),
        .I3(minusOp[32]),
        .I4(minusOp[30]),
        .O(\mcreg[31]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \mcreg[32]_i_1 
       (.I0(\mcreg_reg[32]_i_2_n_4 ),
        .I1(\mcreg_reg[33]_i_2_n_7 ),
        .I2(\modsqr/mcreg_reg_n_0_[31] ),
        .I3(sqrrdy),
        .O(\mcreg[32]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \mcreg[32]_i_1__0 
       (.I0(minusOp[31]),
        .I1(minusOp[32]),
        .I2(mcreg[31]),
        .I3(multrdy),
        .O(\mcreg[32]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[32]_i_3 
       (.I0(\modsqr/mcreg_reg_n_0_[31] ),
        .I1(\modsqr/modreg1_reg_n_0_[31] ),
        .O(\mcreg[32]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[32]_i_3__0 
       (.I0(mcreg[31]),
        .I1(modreg1[31]),
        .O(\mcreg[32]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[32]_i_4 
       (.I0(\modsqr/mcreg_reg_n_0_[30] ),
        .I1(\modsqr/modreg1_reg_n_0_[30] ),
        .O(\mcreg[32]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[32]_i_4__0 
       (.I0(mcreg[30]),
        .I1(modreg1[30]),
        .O(\mcreg[32]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[32]_i_5 
       (.I0(\modsqr/mcreg_reg_n_0_[29] ),
        .I1(\modsqr/modreg1_reg_n_0_[29] ),
        .O(\mcreg[32]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[32]_i_5__0 
       (.I0(mcreg[29]),
        .I1(modreg1[29]),
        .O(\mcreg[32]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[32]_i_6 
       (.I0(\modsqr/mcreg_reg_n_0_[28] ),
        .I1(\modsqr/modreg1_reg_n_0_[28] ),
        .O(\mcreg[32]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[32]_i_6__0 
       (.I0(mcreg[28]),
        .I1(modreg1[28]),
        .O(\mcreg[32]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \mcreg[33]_i_1 
       (.I0(sqrrdy),
        .I1(\mcreg_reg[33]_i_2_n_7 ),
        .I2(\modsqr/mcreg_reg_n_0_[32] ),
        .O(\mcreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \mcreg[33]_i_1__0 
       (.I0(multrdy),
        .I1(minusOp[32]),
        .I2(mcreg[32]),
        .O(\mcreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \mcreg[33]_i_3 
       (.I0(mcreg[32]),
        .O(\mcreg[33]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \mcreg[33]_i_3__0 
       (.I0(\modsqr/mcreg_reg_n_0_[32] ),
        .O(\mcreg[33]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[3]_i_1 
       (.I0(root[3]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[2] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[4]_i_2_n_5 ),
        .O(\mcreg[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[3]_i_1__0 
       (.I0(tempin[3]),
        .I1(multrdy),
        .I2(mcreg[2]),
        .I3(minusOp[32]),
        .I4(minusOp[2]),
        .O(\mcreg[3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[4]_i_1 
       (.I0(root[4]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[3] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[4]_i_2_n_4 ),
        .O(\mcreg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[4]_i_1__0 
       (.I0(tempin[4]),
        .I1(multrdy),
        .I2(mcreg[3]),
        .I3(minusOp[32]),
        .I4(minusOp[3]),
        .O(\mcreg[4]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[4]_i_3 
       (.I0(\modsqr/mcreg_reg_n_0_[3] ),
        .I1(\modsqr/modreg1_reg_n_0_[3] ),
        .O(\mcreg[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[4]_i_3__0 
       (.I0(mcreg[3]),
        .I1(modreg1[3]),
        .O(\mcreg[4]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[4]_i_4 
       (.I0(\modsqr/mcreg_reg_n_0_[2] ),
        .I1(\modsqr/modreg1_reg_n_0_[2] ),
        .O(\mcreg[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[4]_i_4__0 
       (.I0(mcreg[2]),
        .I1(modreg1[2]),
        .O(\mcreg[4]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[4]_i_5 
       (.I0(\modsqr/mcreg_reg_n_0_[1] ),
        .I1(\modsqr/modreg1_reg_n_0_[1] ),
        .O(\mcreg[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[4]_i_5__0 
       (.I0(mcreg[1]),
        .I1(modreg1[1]),
        .O(\mcreg[4]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[4]_i_6 
       (.I0(\modsqr/mcreg_reg_n_0_ ),
        .I1(\modsqr/modreg2_reg_n_0_ ),
        .O(\mcreg[4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[4]_i_6__0 
       (.I0(mcreg[0]),
        .I1(modreg2),
        .O(\mcreg[4]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[5]_i_1 
       (.I0(root[5]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[4] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[8]_i_2_n_7 ),
        .O(\mcreg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[5]_i_1__0 
       (.I0(tempin[5]),
        .I1(multrdy),
        .I2(mcreg[4]),
        .I3(minusOp[32]),
        .I4(minusOp[4]),
        .O(\mcreg[5]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[6]_i_1 
       (.I0(root[6]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[5] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[8]_i_2_n_6 ),
        .O(\mcreg[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[6]_i_1__0 
       (.I0(tempin[6]),
        .I1(multrdy),
        .I2(mcreg[5]),
        .I3(minusOp[32]),
        .I4(minusOp[5]),
        .O(\mcreg[6]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[7]_i_1 
       (.I0(root[7]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[6] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[8]_i_2_n_5 ),
        .O(\mcreg[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[7]_i_1__0 
       (.I0(tempin[7]),
        .I1(multrdy),
        .I2(mcreg[6]),
        .I3(minusOp[32]),
        .I4(minusOp[6]),
        .O(\mcreg[7]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[8]_i_1 
       (.I0(root[8]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[7] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[8]_i_2_n_4 ),
        .O(\mcreg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[8]_i_1__0 
       (.I0(tempin[8]),
        .I1(multrdy),
        .I2(mcreg[7]),
        .I3(minusOp[32]),
        .I4(minusOp[7]),
        .O(\mcreg[8]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[8]_i_3 
       (.I0(\modsqr/mcreg_reg_n_0_[7] ),
        .I1(\modsqr/modreg1_reg_n_0_[7] ),
        .O(\mcreg[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[8]_i_3__0 
       (.I0(mcreg[7]),
        .I1(modreg1[7]),
        .O(\mcreg[8]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[8]_i_4 
       (.I0(\modsqr/mcreg_reg_n_0_[6] ),
        .I1(\modsqr/modreg1_reg_n_0_[6] ),
        .O(\mcreg[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[8]_i_4__0 
       (.I0(mcreg[6]),
        .I1(modreg1[6]),
        .O(\mcreg[8]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[8]_i_5 
       (.I0(\modsqr/mcreg_reg_n_0_[5] ),
        .I1(\modsqr/modreg1_reg_n_0_[5] ),
        .O(\mcreg[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[8]_i_5__0 
       (.I0(mcreg[5]),
        .I1(modreg1[5]),
        .O(\mcreg[8]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[8]_i_6 
       (.I0(\modsqr/mcreg_reg_n_0_[4] ),
        .I1(\modsqr/modreg1_reg_n_0_[4] ),
        .O(\mcreg[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \mcreg[8]_i_6__0 
       (.I0(mcreg[4]),
        .I1(modreg1[4]),
        .O(\mcreg[8]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[9]_i_1 
       (.I0(root[9]),
        .I1(sqrrdy),
        .I2(\modsqr/mcreg_reg_n_0_[8] ),
        .I3(\mcreg_reg[33]_i_2_n_7 ),
        .I4(\mcreg_reg[12]_i_2_n_7 ),
        .O(\mcreg[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \mcreg[9]_i_1__0 
       (.I0(tempin[9]),
        .I1(multrdy),
        .I2(mcreg[8]),
        .I3(minusOp[32]),
        .I4(minusOp[8]),
        .O(\mcreg[9]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[12]_i_2 
       (.CI(\mcreg_reg[8]_i_2_n_0 ),
        .CO({\mcreg_reg[12]_i_2_n_0 ,\mcreg_reg[12]_i_2_n_1 ,\mcreg_reg[12]_i_2_n_2 ,\mcreg_reg[12]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/mcreg_reg_n_0_[11] ,\modsqr/mcreg_reg_n_0_[10] ,\modsqr/mcreg_reg_n_0_[9] ,\modsqr/mcreg_reg_n_0_[8] }),
        .O({\mcreg_reg[12]_i_2_n_4 ,\mcreg_reg[12]_i_2_n_5 ,\mcreg_reg[12]_i_2_n_6 ,\mcreg_reg[12]_i_2_n_7 }),
        .S({\mcreg[12]_i_3_n_0 ,\mcreg[12]_i_4_n_0 ,\mcreg[12]_i_5_n_0 ,\mcreg[12]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[12]_i_2__0 
       (.CI(\mcreg_reg[8]_i_2__0_n_0 ),
        .CO(mcreg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI(mcreg[11:8]),
        .O(minusOp[11:8]),
        .S({\mcreg[12]_i_3__0_n_0 ,\mcreg[12]_i_4__0_n_0 ,\mcreg[12]_i_5__0_n_0 ,\mcreg[12]_i_6__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[16]_i_2 
       (.CI(\mcreg_reg[12]_i_2_n_0 ),
        .CO({\mcreg_reg[16]_i_2_n_0 ,\mcreg_reg[16]_i_2_n_1 ,\mcreg_reg[16]_i_2_n_2 ,\mcreg_reg[16]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/mcreg_reg_n_0_[15] ,\modsqr/mcreg_reg_n_0_[14] ,\modsqr/mcreg_reg_n_0_[13] ,\modsqr/mcreg_reg_n_0_[12] }),
        .O({\mcreg_reg[16]_i_2_n_4 ,\mcreg_reg[16]_i_2_n_5 ,\mcreg_reg[16]_i_2_n_6 ,\mcreg_reg[16]_i_2_n_7 }),
        .S({\mcreg[16]_i_3_n_0 ,\mcreg[16]_i_4_n_0 ,\mcreg[16]_i_5_n_0 ,\mcreg[16]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[16]_i_2__0 
       (.CI(mcreg_reg[3]),
        .CO({\mcreg_reg[16]_i_2__0_n_0 ,\mcreg_reg[16]_i_2__0_n_1 ,\mcreg_reg[16]_i_2__0_n_2 ,\mcreg_reg[16]_i_2__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(mcreg[15:12]),
        .O(minusOp[15:12]),
        .S({\mcreg[16]_i_3__0_n_0 ,\mcreg[16]_i_4__0_n_0 ,\mcreg[16]_i_5__0_n_0 ,\mcreg[16]_i_6__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[20]_i_2 
       (.CI(\mcreg_reg[16]_i_2_n_0 ),
        .CO({\mcreg_reg[20]_i_2_n_0 ,\mcreg_reg[20]_i_2_n_1 ,\mcreg_reg[20]_i_2_n_2 ,\mcreg_reg[20]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/mcreg_reg_n_0_[19] ,\modsqr/mcreg_reg_n_0_[18] ,\modsqr/mcreg_reg_n_0_[17] ,\modsqr/mcreg_reg_n_0_[16] }),
        .O({\mcreg_reg[20]_i_2_n_4 ,\mcreg_reg[20]_i_2_n_5 ,\mcreg_reg[20]_i_2_n_6 ,\mcreg_reg[20]_i_2_n_7 }),
        .S({\mcreg[20]_i_3_n_0 ,\mcreg[20]_i_4_n_0 ,\mcreg[20]_i_5_n_0 ,\mcreg[20]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[20]_i_2__0 
       (.CI(\mcreg_reg[16]_i_2__0_n_0 ),
        .CO({\mcreg_reg[20]_i_2__0_n_0 ,\mcreg_reg[20]_i_2__0_n_1 ,\mcreg_reg[20]_i_2__0_n_2 ,\mcreg_reg[20]_i_2__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(mcreg[19:16]),
        .O(minusOp[19:16]),
        .S({\mcreg[20]_i_3__0_n_0 ,\mcreg[20]_i_4__0_n_0 ,\mcreg[20]_i_5__0_n_0 ,\mcreg[20]_i_6__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[24]_i_2 
       (.CI(\mcreg_reg[20]_i_2_n_0 ),
        .CO({\mcreg_reg[24]_i_2_n_0 ,\mcreg_reg[24]_i_2_n_1 ,\mcreg_reg[24]_i_2_n_2 ,\mcreg_reg[24]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/mcreg_reg_n_0_[23] ,\modsqr/mcreg_reg_n_0_[22] ,\modsqr/mcreg_reg_n_0_[21] ,\modsqr/mcreg_reg_n_0_[20] }),
        .O({\mcreg_reg[24]_i_2_n_4 ,\mcreg_reg[24]_i_2_n_5 ,\mcreg_reg[24]_i_2_n_6 ,\mcreg_reg[24]_i_2_n_7 }),
        .S({\mcreg[24]_i_3_n_0 ,\mcreg[24]_i_4_n_0 ,\mcreg[24]_i_5_n_0 ,\mcreg[24]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[24]_i_2__0 
       (.CI(\mcreg_reg[20]_i_2__0_n_0 ),
        .CO({\mcreg_reg[24]_i_2__0_n_0 ,\mcreg_reg[24]_i_2__0_n_1 ,\mcreg_reg[24]_i_2__0_n_2 ,\mcreg_reg[24]_i_2__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(mcreg[23:20]),
        .O(minusOp[23:20]),
        .S({\mcreg[24]_i_3__0_n_0 ,\mcreg[24]_i_4__0_n_0 ,\mcreg[24]_i_5__0_n_0 ,\mcreg[24]_i_6__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[28]_i_2 
       (.CI(\mcreg_reg[24]_i_2_n_0 ),
        .CO({\mcreg_reg[28]_i_2_n_0 ,\mcreg_reg[28]_i_2_n_1 ,\mcreg_reg[28]_i_2_n_2 ,\mcreg_reg[28]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/mcreg_reg_n_0_[27] ,\modsqr/mcreg_reg_n_0_[26] ,\modsqr/mcreg_reg_n_0_[25] ,\modsqr/mcreg_reg_n_0_[24] }),
        .O({\mcreg_reg[28]_i_2_n_4 ,\mcreg_reg[28]_i_2_n_5 ,\mcreg_reg[28]_i_2_n_6 ,\mcreg_reg[28]_i_2_n_7 }),
        .S({\mcreg[28]_i_3_n_0 ,\mcreg[28]_i_4_n_0 ,\mcreg[28]_i_5_n_0 ,\mcreg[28]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[28]_i_2__0 
       (.CI(\mcreg_reg[24]_i_2__0_n_0 ),
        .CO({\mcreg_reg[28]_i_2__0_n_0 ,\mcreg_reg[28]_i_2__0_n_1 ,\mcreg_reg[28]_i_2__0_n_2 ,\mcreg_reg[28]_i_2__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(mcreg[27:24]),
        .O(minusOp[27:24]),
        .S({\mcreg[28]_i_3__0_n_0 ,\mcreg[28]_i_4__0_n_0 ,\mcreg[28]_i_5__0_n_0 ,\mcreg[28]_i_6__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[32]_i_2 
       (.CI(\mcreg_reg[28]_i_2_n_0 ),
        .CO({\mcreg_reg[32]_i_2_n_0 ,\mcreg_reg[32]_i_2_n_1 ,\mcreg_reg[32]_i_2_n_2 ,\mcreg_reg[32]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/mcreg_reg_n_0_[31] ,\modsqr/mcreg_reg_n_0_[30] ,\modsqr/mcreg_reg_n_0_[29] ,\modsqr/mcreg_reg_n_0_[28] }),
        .O({\mcreg_reg[32]_i_2_n_4 ,\mcreg_reg[32]_i_2_n_5 ,\mcreg_reg[32]_i_2_n_6 ,\mcreg_reg[32]_i_2_n_7 }),
        .S({\mcreg[32]_i_3_n_0 ,\mcreg[32]_i_4_n_0 ,\mcreg[32]_i_5_n_0 ,\mcreg[32]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[32]_i_2__0 
       (.CI(\mcreg_reg[28]_i_2__0_n_0 ),
        .CO({\mcreg_reg[32]_i_2__0_n_0 ,\mcreg_reg[32]_i_2__0_n_1 ,\mcreg_reg[32]_i_2__0_n_2 ,\mcreg_reg[32]_i_2__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(mcreg[31:28]),
        .O(minusOp[31:28]),
        .S({\mcreg[32]_i_3__0_n_0 ,\mcreg[32]_i_4__0_n_0 ,\mcreg[32]_i_5__0_n_0 ,\mcreg[32]_i_6__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[33]_i_2 
       (.CI(\mcreg_reg[32]_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\mcreg_reg[33]_i_2_n_4 ,\mcreg_reg[33]_i_2_n_5 ,\mcreg_reg[33]_i_2_n_6 ,\mcreg_reg[33]_i_2_n_7 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\mcreg[33]_i_3__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[33]_i_2__0 
       (.CI(\mcreg_reg[32]_i_2__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\mcreg_reg[33]_i_2__0_n_4 ,\mcreg_reg[33]_i_2__0_n_5 ,\mcreg_reg[33]_i_2__0_n_6 ,minusOp[32]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\mcreg[33]_i_3_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[4]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\mcreg_reg[4]_i_2_n_0 ,\mcreg_reg[4]_i_2_n_1 ,\mcreg_reg[4]_i_2_n_2 ,\mcreg_reg[4]_i_2_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\modsqr/mcreg_reg_n_0_[3] ,\modsqr/mcreg_reg_n_0_[2] ,\modsqr/mcreg_reg_n_0_[1] ,\modsqr/mcreg_reg_n_0_ }),
        .O({\mcreg_reg[4]_i_2_n_4 ,\mcreg_reg[4]_i_2_n_5 ,\mcreg_reg[4]_i_2_n_6 ,\mcreg_reg[4]_i_2_n_7 }),
        .S({\mcreg[4]_i_3_n_0 ,\mcreg[4]_i_4_n_0 ,\mcreg[4]_i_5_n_0 ,\mcreg[4]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[4]_i_2__0 
       (.CI(\<const0>__0__0 ),
        .CO({\mcreg_reg[4]_i_2__0_n_0 ,\mcreg_reg[4]_i_2__0_n_1 ,\mcreg_reg[4]_i_2__0_n_2 ,\mcreg_reg[4]_i_2__0_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI(mcreg[3:0]),
        .O(minusOp[3:0]),
        .S({\mcreg[4]_i_3__0_n_0 ,\mcreg[4]_i_4__0_n_0 ,\mcreg[4]_i_5__0_n_0 ,\mcreg[4]_i_6__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[8]_i_2 
       (.CI(\mcreg_reg[4]_i_2_n_0 ),
        .CO({\mcreg_reg[8]_i_2_n_0 ,\mcreg_reg[8]_i_2_n_1 ,\mcreg_reg[8]_i_2_n_2 ,\mcreg_reg[8]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/mcreg_reg_n_0_[7] ,\modsqr/mcreg_reg_n_0_[6] ,\modsqr/mcreg_reg_n_0_[5] ,\modsqr/mcreg_reg_n_0_[4] }),
        .O({\mcreg_reg[8]_i_2_n_4 ,\mcreg_reg[8]_i_2_n_5 ,\mcreg_reg[8]_i_2_n_6 ,\mcreg_reg[8]_i_2_n_7 }),
        .S({\mcreg[8]_i_3_n_0 ,\mcreg[8]_i_4_n_0 ,\mcreg[8]_i_5_n_0 ,\mcreg[8]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \mcreg_reg[8]_i_2__0 
       (.CI(\mcreg_reg[4]_i_2__0_n_0 ),
        .CO({\mcreg_reg[8]_i_2__0_n_0 ,\mcreg_reg[8]_i_2__0_n_1 ,\mcreg_reg[8]_i_2__0_n_2 ,\mcreg_reg[8]_i_2__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(mcreg[7:4]),
        .O(minusOp[7:4]),
        .S({\mcreg[8]_i_3__0_n_0 ,\mcreg[8]_i_4__0_n_0 ,\mcreg[8]_i_5__0_n_0 ,\mcreg[8]_i_6__0_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__0_i_1
       (.I0(\modsqr/plusOp_carry__0_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[7] ),
        .O(minusOp_inferred__0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__0_i_1__0
       (.I0(prodreg1[7]),
        .I1(modreg1[7]),
        .O(minusOp_inferred__0_carry__0_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__0_i_2
       (.I0(\modsqr/plusOp_carry__0_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[6] ),
        .O(minusOp_inferred__0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__0_i_2__0
       (.I0(prodreg1[6]),
        .I1(modreg1[6]),
        .O(minusOp_inferred__0_carry__0_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__0_i_3
       (.I0(\modsqr/plusOp_carry__0_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[5] ),
        .O(minusOp_inferred__0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__0_i_3__0
       (.I0(prodreg1[5]),
        .I1(modreg1[5]),
        .O(minusOp_inferred__0_carry__0_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__0_i_4
       (.I0(\modsqr/plusOp_carry__0_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[4] ),
        .O(minusOp_inferred__0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__0_i_4__0
       (.I0(prodreg1[4]),
        .I1(modreg1[4]),
        .O(minusOp_inferred__0_carry__0_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__1_i_1
       (.I0(\modsqr/plusOp_carry__1_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[11] ),
        .O(minusOp_inferred__0_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__1_i_1__0
       (.I0(prodreg1[11]),
        .I1(modreg1[11]),
        .O(minusOp_inferred__0_carry__1_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__1_i_2
       (.I0(\modsqr/plusOp_carry__1_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_ ),
        .O(minusOp_inferred__0_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__1_i_2__0
       (.I0(prodreg1[10]),
        .I1(modreg1[10]),
        .O(minusOp_inferred__0_carry__1_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__1_i_3
       (.I0(\modsqr/plusOp_carry__1_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[9] ),
        .O(minusOp_inferred__0_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__1_i_3__0
       (.I0(prodreg1[9]),
        .I1(modreg1[9]),
        .O(minusOp_inferred__0_carry__1_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__1_i_4
       (.I0(\modsqr/plusOp_carry__1_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[8] ),
        .O(minusOp_inferred__0_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__1_i_4__0
       (.I0(prodreg1[8]),
        .I1(modreg1[8]),
        .O(minusOp_inferred__0_carry__1_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__2_i_1
       (.I0(\modsqr/plusOp_carry__2_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[15] ),
        .O(minusOp_inferred__0_carry__2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__2_i_1__0
       (.I0(prodreg1[15]),
        .I1(modreg1[15]),
        .O(minusOp_inferred__0_carry__2_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__2_i_2
       (.I0(\modsqr/plusOp_carry__2_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[14] ),
        .O(minusOp_inferred__0_carry__2_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__2_i_2__0
       (.I0(prodreg1[14]),
        .I1(modreg1[14]),
        .O(minusOp_inferred__0_carry__2_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__2_i_3
       (.I0(\modsqr/plusOp_carry__2_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[13] ),
        .O(minusOp_inferred__0_carry__2_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__2_i_3__0
       (.I0(prodreg1[13]),
        .I1(modreg1[13]),
        .O(minusOp_inferred__0_carry__2_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__2_i_4
       (.I0(\modsqr/plusOp_carry__2_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[12] ),
        .O(minusOp_inferred__0_carry__2_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__2_i_4__0
       (.I0(prodreg1[12]),
        .I1(modreg1[12]),
        .O(minusOp_inferred__0_carry__2_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__3_i_1
       (.I0(\modsqr/plusOp_carry__3_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[19] ),
        .O(minusOp_inferred__0_carry__3_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__3_i_1__0
       (.I0(prodreg1[19]),
        .I1(modreg1[19]),
        .O(minusOp_inferred__0_carry__3_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__3_i_2
       (.I0(\modsqr/plusOp_carry__3_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[18] ),
        .O(minusOp_inferred__0_carry__3_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__3_i_2__0
       (.I0(prodreg1[18]),
        .I1(modreg1[18]),
        .O(minusOp_inferred__0_carry__3_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__3_i_3
       (.I0(\modsqr/plusOp_carry__3_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[17] ),
        .O(minusOp_inferred__0_carry__3_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__3_i_3__0
       (.I0(prodreg1[17]),
        .I1(modreg1[17]),
        .O(minusOp_inferred__0_carry__3_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__3_i_4
       (.I0(\modsqr/plusOp_carry__3_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[16] ),
        .O(minusOp_inferred__0_carry__3_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__3_i_4__0
       (.I0(prodreg1[16]),
        .I1(modreg1[16]),
        .O(minusOp_inferred__0_carry__3_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__4_i_1
       (.I0(\modsqr/plusOp_carry__4_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[23] ),
        .O(minusOp_inferred__0_carry__4_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__4_i_1__0
       (.I0(prodreg1[23]),
        .I1(modreg1[23]),
        .O(minusOp_inferred__0_carry__4_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__4_i_2
       (.I0(\modsqr/plusOp_carry__4_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[22] ),
        .O(minusOp_inferred__0_carry__4_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__4_i_2__0
       (.I0(prodreg1[22]),
        .I1(modreg1[22]),
        .O(minusOp_inferred__0_carry__4_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__4_i_3
       (.I0(\modsqr/plusOp_carry__4_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[21] ),
        .O(minusOp_inferred__0_carry__4_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__4_i_3__0
       (.I0(prodreg1[21]),
        .I1(modreg1[21]),
        .O(minusOp_inferred__0_carry__4_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__4_i_4
       (.I0(\modsqr/plusOp_carry__4_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[20] ),
        .O(minusOp_inferred__0_carry__4_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__4_i_4__0
       (.I0(prodreg1[20]),
        .I1(modreg1[20]),
        .O(minusOp_inferred__0_carry__4_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__5_i_1
       (.I0(\modsqr/plusOp_carry__5_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[27] ),
        .O(minusOp_inferred__0_carry__5_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__5_i_1__0
       (.I0(prodreg1[27]),
        .I1(modreg1[27]),
        .O(minusOp_inferred__0_carry__5_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__5_i_2
       (.I0(\modsqr/plusOp_carry__5_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[26] ),
        .O(minusOp_inferred__0_carry__5_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__5_i_2__0
       (.I0(prodreg1[26]),
        .I1(modreg1[26]),
        .O(minusOp_inferred__0_carry__5_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__5_i_3
       (.I0(\modsqr/plusOp_carry__5_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[25] ),
        .O(minusOp_inferred__0_carry__5_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__5_i_3__0
       (.I0(prodreg1[25]),
        .I1(modreg1[25]),
        .O(minusOp_inferred__0_carry__5_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__5_i_4
       (.I0(\modsqr/plusOp_carry__5_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[24] ),
        .O(minusOp_inferred__0_carry__5_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__5_i_4__0
       (.I0(prodreg1[24]),
        .I1(modreg1[24]),
        .O(minusOp_inferred__0_carry__5_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__6_i_1
       (.I0(\modsqr/plusOp_carry__6_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[31] ),
        .O(minusOp_inferred__0_carry__6_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__6_i_1__0
       (.I0(prodreg1[31]),
        .I1(modreg1[31]),
        .O(minusOp_inferred__0_carry__6_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__6_i_2
       (.I0(\modsqr/plusOp_carry__6_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[30] ),
        .O(minusOp_inferred__0_carry__6_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__6_i_2__0
       (.I0(prodreg1[30]),
        .I1(modreg1[30]),
        .O(minusOp_inferred__0_carry__6_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__6_i_3
       (.I0(\modsqr/plusOp_carry__6_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[29] ),
        .O(minusOp_inferred__0_carry__6_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__6_i_3__0
       (.I0(prodreg1[29]),
        .I1(modreg1[29]),
        .O(minusOp_inferred__0_carry__6_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__6_i_4
       (.I0(\modsqr/plusOp_carry__6_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[28] ),
        .O(minusOp_inferred__0_carry__6_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__6_i_4__0
       (.I0(prodreg1[28]),
        .I1(modreg1[28]),
        .O(minusOp_inferred__0_carry__6_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    minusOp_inferred__0_carry__7_i_1
       (.I0(\modsqr/plusOp_carry__7_n_6 ),
        .O(minusOp_inferred__0_carry__7_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    minusOp_inferred__0_carry__7_i_1__0
       (.I0(prodreg1[33]),
        .O(minusOp_inferred__0_carry__7_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    minusOp_inferred__0_carry__7_i_2
       (.I0(\modsqr/plusOp_carry__7_n_7 ),
        .O(minusOp_inferred__0_carry__7_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    minusOp_inferred__0_carry__7_i_2__0
       (.I0(prodreg1[32]),
        .O(minusOp_inferred__0_carry__7_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry_i_1
       (.I0(\modsqr/plusOp_carry_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[3] ),
        .O(minusOp_inferred__0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry_i_1__0
       (.I0(prodreg1[3]),
        .I1(modreg1[3]),
        .O(minusOp_inferred__0_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry_i_2
       (.I0(\modsqr/plusOp_carry_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[2] ),
        .O(minusOp_inferred__0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry_i_2__0
       (.I0(prodreg1[2]),
        .I1(modreg1[2]),
        .O(minusOp_inferred__0_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry_i_3
       (.I0(\modsqr/plusOp_carry_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[1] ),
        .O(minusOp_inferred__0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry_i_3__0
       (.I0(prodreg1[1]),
        .I1(modreg1[1]),
        .O(minusOp_inferred__0_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry_i_4
       (.I0(\modsqr/plusOp_carry_n_7 ),
        .I1(\modsqr/modreg2_reg_n_0_ ),
        .O(minusOp_inferred__0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry_i_4__0
       (.I0(prodreg1[0]),
        .I1(modreg2),
        .O(minusOp_inferred__0_carry_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__0_i_1
       (.I0(\modsqr/plusOp_carry__0_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[6] ),
        .O(minusOp_inferred__1_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__0_i_1__0
       (.I0(prodreg1[7]),
        .I1(modreg1[6]),
        .O(minusOp_inferred__1_carry__0_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__0_i_2
       (.I0(\modsqr/plusOp_carry__0_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[5] ),
        .O(minusOp_inferred__1_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__0_i_2__0
       (.I0(prodreg1[6]),
        .I1(modreg1[5]),
        .O(minusOp_inferred__1_carry__0_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__0_i_3
       (.I0(\modsqr/plusOp_carry__0_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[4] ),
        .O(minusOp_inferred__1_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__0_i_3__0
       (.I0(prodreg1[5]),
        .I1(modreg1[4]),
        .O(minusOp_inferred__1_carry__0_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__0_i_4
       (.I0(\modsqr/plusOp_carry__0_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[3] ),
        .O(minusOp_inferred__1_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__0_i_4__0
       (.I0(prodreg1[4]),
        .I1(modreg1[3]),
        .O(minusOp_inferred__1_carry__0_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__1_i_1
       (.I0(\modsqr/plusOp_carry__1_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_ ),
        .O(minusOp_inferred__1_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__1_i_1__0
       (.I0(prodreg1[11]),
        .I1(modreg1[10]),
        .O(minusOp_inferred__1_carry__1_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__1_i_2
       (.I0(\modsqr/plusOp_carry__1_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[9] ),
        .O(minusOp_inferred__1_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__1_i_2__0
       (.I0(prodreg1[10]),
        .I1(modreg1[9]),
        .O(minusOp_inferred__1_carry__1_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__1_i_3
       (.I0(\modsqr/plusOp_carry__1_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[8] ),
        .O(minusOp_inferred__1_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__1_i_3__0
       (.I0(prodreg1[9]),
        .I1(modreg1[8]),
        .O(minusOp_inferred__1_carry__1_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__1_i_4
       (.I0(\modsqr/plusOp_carry__1_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[7] ),
        .O(minusOp_inferred__1_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__1_i_4__0
       (.I0(prodreg1[8]),
        .I1(modreg1[7]),
        .O(minusOp_inferred__1_carry__1_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__2_i_1
       (.I0(\modsqr/plusOp_carry__2_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[14] ),
        .O(minusOp_inferred__1_carry__2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__2_i_1__0
       (.I0(prodreg1[15]),
        .I1(modreg1[14]),
        .O(minusOp_inferred__1_carry__2_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__2_i_2
       (.I0(\modsqr/plusOp_carry__2_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[13] ),
        .O(minusOp_inferred__1_carry__2_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__2_i_2__0
       (.I0(prodreg1[14]),
        .I1(modreg1[13]),
        .O(minusOp_inferred__1_carry__2_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__2_i_3
       (.I0(\modsqr/plusOp_carry__2_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[12] ),
        .O(minusOp_inferred__1_carry__2_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__2_i_3__0
       (.I0(prodreg1[13]),
        .I1(modreg1[12]),
        .O(minusOp_inferred__1_carry__2_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__2_i_4
       (.I0(\modsqr/plusOp_carry__2_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[11] ),
        .O(minusOp_inferred__1_carry__2_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__2_i_4__0
       (.I0(prodreg1[12]),
        .I1(modreg1[11]),
        .O(minusOp_inferred__1_carry__2_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__3_i_1
       (.I0(\modsqr/plusOp_carry__3_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[18] ),
        .O(minusOp_inferred__1_carry__3_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__3_i_1__0
       (.I0(prodreg1[19]),
        .I1(modreg1[18]),
        .O(minusOp_inferred__1_carry__3_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__3_i_2
       (.I0(\modsqr/plusOp_carry__3_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[17] ),
        .O(minusOp_inferred__1_carry__3_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__3_i_2__0
       (.I0(prodreg1[18]),
        .I1(modreg1[17]),
        .O(minusOp_inferred__1_carry__3_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__3_i_3
       (.I0(\modsqr/plusOp_carry__3_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[16] ),
        .O(minusOp_inferred__1_carry__3_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__3_i_3__0
       (.I0(prodreg1[17]),
        .I1(modreg1[16]),
        .O(minusOp_inferred__1_carry__3_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__3_i_4
       (.I0(\modsqr/plusOp_carry__3_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[15] ),
        .O(minusOp_inferred__1_carry__3_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__3_i_4__0
       (.I0(prodreg1[16]),
        .I1(modreg1[15]),
        .O(minusOp_inferred__1_carry__3_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__4_i_1
       (.I0(\modsqr/plusOp_carry__4_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[22] ),
        .O(minusOp_inferred__1_carry__4_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__4_i_1__0
       (.I0(prodreg1[23]),
        .I1(modreg1[22]),
        .O(minusOp_inferred__1_carry__4_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__4_i_2
       (.I0(\modsqr/plusOp_carry__4_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[21] ),
        .O(minusOp_inferred__1_carry__4_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__4_i_2__0
       (.I0(prodreg1[22]),
        .I1(modreg1[21]),
        .O(minusOp_inferred__1_carry__4_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__4_i_3
       (.I0(\modsqr/plusOp_carry__4_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[20] ),
        .O(minusOp_inferred__1_carry__4_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__4_i_3__0
       (.I0(prodreg1[21]),
        .I1(modreg1[20]),
        .O(minusOp_inferred__1_carry__4_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__4_i_4
       (.I0(\modsqr/plusOp_carry__4_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[19] ),
        .O(minusOp_inferred__1_carry__4_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__4_i_4__0
       (.I0(prodreg1[20]),
        .I1(modreg1[19]),
        .O(minusOp_inferred__1_carry__4_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__5_i_1
       (.I0(\modsqr/plusOp_carry__5_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[26] ),
        .O(minusOp_inferred__1_carry__5_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__5_i_1__0
       (.I0(prodreg1[27]),
        .I1(modreg1[26]),
        .O(minusOp_inferred__1_carry__5_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__5_i_2
       (.I0(\modsqr/plusOp_carry__5_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[25] ),
        .O(minusOp_inferred__1_carry__5_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__5_i_2__0
       (.I0(prodreg1[26]),
        .I1(modreg1[25]),
        .O(minusOp_inferred__1_carry__5_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__5_i_3
       (.I0(\modsqr/plusOp_carry__5_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[24] ),
        .O(minusOp_inferred__1_carry__5_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__5_i_3__0
       (.I0(prodreg1[25]),
        .I1(modreg1[24]),
        .O(minusOp_inferred__1_carry__5_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__5_i_4
       (.I0(\modsqr/plusOp_carry__5_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[23] ),
        .O(minusOp_inferred__1_carry__5_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__5_i_4__0
       (.I0(prodreg1[24]),
        .I1(modreg1[23]),
        .O(minusOp_inferred__1_carry__5_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__6_i_1
       (.I0(\modsqr/plusOp_carry__6_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[30] ),
        .O(minusOp_inferred__1_carry__6_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__6_i_1__0
       (.I0(prodreg1[31]),
        .I1(modreg1[30]),
        .O(minusOp_inferred__1_carry__6_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__6_i_2
       (.I0(\modsqr/plusOp_carry__6_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[29] ),
        .O(minusOp_inferred__1_carry__6_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__6_i_2__0
       (.I0(prodreg1[30]),
        .I1(modreg1[29]),
        .O(minusOp_inferred__1_carry__6_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__6_i_3
       (.I0(\modsqr/plusOp_carry__6_n_6 ),
        .I1(\modsqr/modreg1_reg_n_0_[28] ),
        .O(minusOp_inferred__1_carry__6_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__6_i_3__0
       (.I0(prodreg1[29]),
        .I1(modreg1[28]),
        .O(minusOp_inferred__1_carry__6_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__6_i_4
       (.I0(\modsqr/plusOp_carry__6_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[27] ),
        .O(minusOp_inferred__1_carry__6_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__6_i_4__0
       (.I0(prodreg1[28]),
        .I1(modreg1[27]),
        .O(minusOp_inferred__1_carry__6_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    minusOp_inferred__1_carry__7_i_1
       (.I0(prodreg1[33]),
        .O(minusOp_inferred__1_carry__7_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    minusOp_inferred__1_carry__7_i_1__0
       (.I0(\modsqr/plusOp_carry__7_n_6 ),
        .O(minusOp_inferred__1_carry__7_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__7_i_2
       (.I0(\modsqr/plusOp_carry__7_n_7 ),
        .I1(\modsqr/modreg1_reg_n_0_[31] ),
        .O(minusOp_inferred__1_carry__7_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry__7_i_2__0
       (.I0(prodreg1[32]),
        .I1(modreg1[31]),
        .O(minusOp_inferred__1_carry__7_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry_i_1
       (.I0(\modsqr/plusOp_carry_n_4 ),
        .I1(\modsqr/modreg1_reg_n_0_[2] ),
        .O(minusOp_inferred__1_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry_i_1__0
       (.I0(prodreg1[3]),
        .I1(modreg1[2]),
        .O(minusOp_inferred__1_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry_i_2
       (.I0(\modsqr/plusOp_carry_n_5 ),
        .I1(\modsqr/modreg1_reg_n_0_[1] ),
        .O(minusOp_inferred__1_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry_i_2__0
       (.I0(prodreg1[2]),
        .I1(modreg1[1]),
        .O(minusOp_inferred__1_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry_i_3
       (.I0(\modsqr/plusOp_carry_n_6 ),
        .I1(\modsqr/modreg2_reg_n_0_ ),
        .O(minusOp_inferred__1_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__1_carry_i_3__0
       (.I0(prodreg1[1]),
        .I1(modreg2),
        .O(minusOp_inferred__1_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    minusOp_inferred__1_carry_i_4
       (.I0(\modsqr/plusOp_carry_n_7 ),
        .O(minusOp_inferred__1_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    minusOp_inferred__1_carry_i_4__0
       (.I0(prodreg1[0]),
        .O(minusOp_inferred__1_carry_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \modmultiply/first_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(first_i_1_n_0),
        .PRE(reset),
        .Q(multrdy));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[0] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[0]_i_1__0_n_0 ),
        .Q(mcreg[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[10] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[10]_i_1__0_n_0 ),
        .Q(mcreg[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[11] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[11]_i_1__0_n_0 ),
        .Q(mcreg[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[12] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[12]_i_1__0_n_0 ),
        .Q(mcreg[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[13] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[13]_i_1__0_n_0 ),
        .Q(mcreg[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[14] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[14]_i_1__0_n_0 ),
        .Q(mcreg[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[15] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[15]_i_1__0_n_0 ),
        .Q(mcreg[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[16] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[16]_i_1__0_n_0 ),
        .Q(mcreg[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[17] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[17]_i_1__0_n_0 ),
        .Q(mcreg[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[18] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[18]_i_1__0_n_0 ),
        .Q(mcreg[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[19] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[19]_i_1__0_n_0 ),
        .Q(mcreg[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[1] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[1]_i_1__0_n_0 ),
        .Q(mcreg[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[20] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[20]_i_1__0_n_0 ),
        .Q(mcreg[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[21] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[21]_i_1__0_n_0 ),
        .Q(mcreg[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[22] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[22]_i_1__0_n_0 ),
        .Q(mcreg[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[23] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[23]_i_1__0_n_0 ),
        .Q(mcreg[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[24] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[24]_i_1__0_n_0 ),
        .Q(mcreg[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[25] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[25]_i_1__0_n_0 ),
        .Q(mcreg[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[26] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[26]_i_1__0_n_0 ),
        .Q(mcreg[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[27] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[27]_i_1__0_n_0 ),
        .Q(mcreg[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[28] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[28]_i_1__0_n_0 ),
        .Q(mcreg[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[29] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[29]_i_1__0_n_0 ),
        .Q(mcreg[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[2] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[2]_i_1__0_n_0 ),
        .Q(mcreg[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[30] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[30]_i_1__0_n_0 ),
        .Q(mcreg[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[31] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[31]_i_1__0_n_0 ),
        .Q(mcreg[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[32] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[32]_i_1__0_n_0 ),
        .Q(mcreg[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[33] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[33]_i_1__0_n_0 ),
        .Q(mcreg[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[3] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[3]_i_1__0_n_0 ),
        .Q(mcreg[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[4] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[4]_i_1__0_n_0 ),
        .Q(mcreg[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[5] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[5]_i_1__0_n_0 ),
        .Q(mcreg[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[6] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[6]_i_1__0_n_0 ),
        .Q(mcreg[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[7] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[7]_i_1__0_n_0 ),
        .Q(mcreg[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[8] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[8]_i_1__0_n_0 ),
        .Q(mcreg[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mcreg_reg[9] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mcreg[9]_i_1__0_n_0 ),
        .Q(mcreg[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\modmultiply/minusOp_inferred__0_carry_n_0 ,\modmultiply/minusOp_inferred__0_carry_n_1 ,\modmultiply/minusOp_inferred__0_carry_n_2 ,\modmultiply/minusOp_inferred__0_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI(prodreg1[3:0]),
        .O({\modmultiply/minusOp_inferred__0_carry_n_4 ,\modmultiply/minusOp_inferred__0_carry_n_5 ,\modmultiply/minusOp_inferred__0_carry_n_6 ,\modmultiply/minusOp_inferred__0_carry_n_7 }),
        .S({minusOp_inferred__0_carry_i_1__0_n_0,minusOp_inferred__0_carry_i_2__0_n_0,minusOp_inferred__0_carry_i_3__0_n_0,minusOp_inferred__0_carry_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__0_carry__0 
       (.CI(\modmultiply/minusOp_inferred__0_carry_n_0 ),
        .CO({\modmultiply/minusOp_inferred__0_carry__0_n_0 ,\modmultiply/minusOp_inferred__0_carry__0_n_1 ,\modmultiply/minusOp_inferred__0_carry__0_n_2 ,\modmultiply/minusOp_inferred__0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[7:4]),
        .O({\modmultiply/minusOp_inferred__0_carry__0_n_4 ,\modmultiply/minusOp_inferred__0_carry__0_n_5 ,\modmultiply/minusOp_inferred__0_carry__0_n_6 ,\modmultiply/minusOp_inferred__0_carry__0_n_7 }),
        .S({minusOp_inferred__0_carry__0_i_1__0_n_0,minusOp_inferred__0_carry__0_i_2__0_n_0,minusOp_inferred__0_carry__0_i_3__0_n_0,minusOp_inferred__0_carry__0_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__0_carry__1 
       (.CI(\modmultiply/minusOp_inferred__0_carry__0_n_0 ),
        .CO({\modmultiply/minusOp_inferred__0_carry__1_n_0 ,\modmultiply/minusOp_inferred__0_carry__1_n_1 ,\modmultiply/minusOp_inferred__0_carry__1_n_2 ,\modmultiply/minusOp_inferred__0_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[11:8]),
        .O({\modmultiply/minusOp_inferred__0_carry__1_n_4 ,\modmultiply/minusOp_inferred__0_carry__1_n_5 ,\modmultiply/minusOp_inferred__0_carry__1_n_6 ,\modmultiply/minusOp_inferred__0_carry__1_n_7 }),
        .S({minusOp_inferred__0_carry__1_i_1__0_n_0,minusOp_inferred__0_carry__1_i_2__0_n_0,minusOp_inferred__0_carry__1_i_3__0_n_0,minusOp_inferred__0_carry__1_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__0_carry__2 
       (.CI(\modmultiply/minusOp_inferred__0_carry__1_n_0 ),
        .CO({\modmultiply/minusOp_inferred__0_carry__2_n_0 ,\modmultiply/minusOp_inferred__0_carry__2_n_1 ,\modmultiply/minusOp_inferred__0_carry__2_n_2 ,\modmultiply/minusOp_inferred__0_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[15:12]),
        .O({\modmultiply/minusOp_inferred__0_carry__2_n_4 ,\modmultiply/minusOp_inferred__0_carry__2_n_5 ,\modmultiply/minusOp_inferred__0_carry__2_n_6 ,\modmultiply/minusOp_inferred__0_carry__2_n_7 }),
        .S({minusOp_inferred__0_carry__2_i_1__0_n_0,minusOp_inferred__0_carry__2_i_2__0_n_0,minusOp_inferred__0_carry__2_i_3__0_n_0,minusOp_inferred__0_carry__2_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__0_carry__3 
       (.CI(\modmultiply/minusOp_inferred__0_carry__2_n_0 ),
        .CO({\modmultiply/minusOp_inferred__0_carry__3_n_0 ,\modmultiply/minusOp_inferred__0_carry__3_n_1 ,\modmultiply/minusOp_inferred__0_carry__3_n_2 ,\modmultiply/minusOp_inferred__0_carry__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[19:16]),
        .O({\modmultiply/minusOp_inferred__0_carry__3_n_4 ,\modmultiply/minusOp_inferred__0_carry__3_n_5 ,\modmultiply/minusOp_inferred__0_carry__3_n_6 ,\modmultiply/minusOp_inferred__0_carry__3_n_7 }),
        .S({minusOp_inferred__0_carry__3_i_1__0_n_0,minusOp_inferred__0_carry__3_i_2__0_n_0,minusOp_inferred__0_carry__3_i_3__0_n_0,minusOp_inferred__0_carry__3_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__0_carry__4 
       (.CI(\modmultiply/minusOp_inferred__0_carry__3_n_0 ),
        .CO({\modmultiply/minusOp_inferred__0_carry__4_n_0 ,\modmultiply/minusOp_inferred__0_carry__4_n_1 ,\modmultiply/minusOp_inferred__0_carry__4_n_2 ,\modmultiply/minusOp_inferred__0_carry__4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[23:20]),
        .O({\modmultiply/minusOp_inferred__0_carry__4_n_4 ,\modmultiply/minusOp_inferred__0_carry__4_n_5 ,\modmultiply/minusOp_inferred__0_carry__4_n_6 ,\modmultiply/minusOp_inferred__0_carry__4_n_7 }),
        .S({minusOp_inferred__0_carry__4_i_1__0_n_0,minusOp_inferred__0_carry__4_i_2__0_n_0,minusOp_inferred__0_carry__4_i_3__0_n_0,minusOp_inferred__0_carry__4_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__0_carry__5 
       (.CI(\modmultiply/minusOp_inferred__0_carry__4_n_0 ),
        .CO({\modmultiply/minusOp_inferred__0_carry__5_n_0 ,\modmultiply/minusOp_inferred__0_carry__5_n_1 ,\modmultiply/minusOp_inferred__0_carry__5_n_2 ,\modmultiply/minusOp_inferred__0_carry__5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[27:24]),
        .O({\modmultiply/minusOp_inferred__0_carry__5_n_4 ,\modmultiply/minusOp_inferred__0_carry__5_n_5 ,\modmultiply/minusOp_inferred__0_carry__5_n_6 ,\modmultiply/minusOp_inferred__0_carry__5_n_7 }),
        .S({minusOp_inferred__0_carry__5_i_1__0_n_0,minusOp_inferred__0_carry__5_i_2__0_n_0,minusOp_inferred__0_carry__5_i_3__0_n_0,minusOp_inferred__0_carry__5_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__0_carry__6 
       (.CI(\modmultiply/minusOp_inferred__0_carry__5_n_0 ),
        .CO({\modmultiply/minusOp_inferred__0_carry__6_n_0 ,\modmultiply/minusOp_inferred__0_carry__6_n_1 ,\modmultiply/minusOp_inferred__0_carry__6_n_2 ,\modmultiply/minusOp_inferred__0_carry__6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[31:28]),
        .O({\modmultiply/minusOp_inferred__0_carry__6_n_4 ,\modmultiply/minusOp_inferred__0_carry__6_n_5 ,\modmultiply/minusOp_inferred__0_carry__6_n_6 ,\modmultiply/minusOp_inferred__0_carry__6_n_7 }),
        .S({minusOp_inferred__0_carry__6_i_1__0_n_0,minusOp_inferred__0_carry__6_i_2__0_n_0,minusOp_inferred__0_carry__6_i_3__0_n_0,minusOp_inferred__0_carry__6_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__0_carry__7 
       (.CI(\modmultiply/minusOp_inferred__0_carry__6_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,prodreg1[32]}),
        .O({\modmultiply/minusOp_inferred__0_carry__7_n_4 ,\modmultiply/minusOp_inferred__0_carry__7_n_5 ,\modmultiply/minusOp_inferred__0_carry__7_n_6 ,\modmultiply/minusOp_inferred__0_carry__7_n_7 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,minusOp_inferred__0_carry__7_i_1__0_n_0,minusOp_inferred__0_carry__7_i_2__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\modmultiply/minusOp_inferred__1_carry_n_0 ,\modmultiply/minusOp_inferred__1_carry_n_1 ,\modmultiply/minusOp_inferred__1_carry_n_2 ,\modmultiply/minusOp_inferred__1_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI(prodreg1[3:0]),
        .O(minusOp0_in[3:0]),
        .S({minusOp_inferred__1_carry_i_1__0_n_0,minusOp_inferred__1_carry_i_2__0_n_0,minusOp_inferred__1_carry_i_3__0_n_0,minusOp_inferred__1_carry_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__1_carry__0 
       (.CI(\modmultiply/minusOp_inferred__1_carry_n_0 ),
        .CO({\modmultiply/minusOp_inferred__1_carry__0_n_0 ,\modmultiply/minusOp_inferred__1_carry__0_n_1 ,\modmultiply/minusOp_inferred__1_carry__0_n_2 ,\modmultiply/minusOp_inferred__1_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[7:4]),
        .O(minusOp0_in[7:4]),
        .S({minusOp_inferred__1_carry__0_i_1__0_n_0,minusOp_inferred__1_carry__0_i_2__0_n_0,minusOp_inferred__1_carry__0_i_3__0_n_0,minusOp_inferred__1_carry__0_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__1_carry__1 
       (.CI(\modmultiply/minusOp_inferred__1_carry__0_n_0 ),
        .CO({\modmultiply/minusOp_inferred__1_carry__1_n_0 ,\modmultiply/minusOp_inferred__1_carry__1_n_1 ,\modmultiply/minusOp_inferred__1_carry__1_n_2 ,\modmultiply/minusOp_inferred__1_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[11:8]),
        .O(minusOp0_in[11:8]),
        .S({minusOp_inferred__1_carry__1_i_1__0_n_0,minusOp_inferred__1_carry__1_i_2__0_n_0,minusOp_inferred__1_carry__1_i_3__0_n_0,minusOp_inferred__1_carry__1_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__1_carry__2 
       (.CI(\modmultiply/minusOp_inferred__1_carry__1_n_0 ),
        .CO({\modmultiply/minusOp_inferred__1_carry__2_n_0 ,\modmultiply/minusOp_inferred__1_carry__2_n_1 ,\modmultiply/minusOp_inferred__1_carry__2_n_2 ,\modmultiply/minusOp_inferred__1_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[15:12]),
        .O(minusOp0_in[15:12]),
        .S({minusOp_inferred__1_carry__2_i_1__0_n_0,minusOp_inferred__1_carry__2_i_2__0_n_0,minusOp_inferred__1_carry__2_i_3__0_n_0,minusOp_inferred__1_carry__2_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__1_carry__3 
       (.CI(\modmultiply/minusOp_inferred__1_carry__2_n_0 ),
        .CO({\modmultiply/minusOp_inferred__1_carry__3_n_0 ,\modmultiply/minusOp_inferred__1_carry__3_n_1 ,\modmultiply/minusOp_inferred__1_carry__3_n_2 ,\modmultiply/minusOp_inferred__1_carry__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[19:16]),
        .O(minusOp0_in[19:16]),
        .S({minusOp_inferred__1_carry__3_i_1__0_n_0,minusOp_inferred__1_carry__3_i_2__0_n_0,minusOp_inferred__1_carry__3_i_3__0_n_0,minusOp_inferred__1_carry__3_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__1_carry__4 
       (.CI(\modmultiply/minusOp_inferred__1_carry__3_n_0 ),
        .CO({\modmultiply/minusOp_inferred__1_carry__4_n_0 ,\modmultiply/minusOp_inferred__1_carry__4_n_1 ,\modmultiply/minusOp_inferred__1_carry__4_n_2 ,\modmultiply/minusOp_inferred__1_carry__4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[23:20]),
        .O(minusOp0_in[23:20]),
        .S({minusOp_inferred__1_carry__4_i_1__0_n_0,minusOp_inferred__1_carry__4_i_2__0_n_0,minusOp_inferred__1_carry__4_i_3__0_n_0,minusOp_inferred__1_carry__4_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__1_carry__5 
       (.CI(\modmultiply/minusOp_inferred__1_carry__4_n_0 ),
        .CO({\modmultiply/minusOp_inferred__1_carry__5_n_0 ,\modmultiply/minusOp_inferred__1_carry__5_n_1 ,\modmultiply/minusOp_inferred__1_carry__5_n_2 ,\modmultiply/minusOp_inferred__1_carry__5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[27:24]),
        .O(minusOp0_in[27:24]),
        .S({minusOp_inferred__1_carry__5_i_1__0_n_0,minusOp_inferred__1_carry__5_i_2__0_n_0,minusOp_inferred__1_carry__5_i_3__0_n_0,minusOp_inferred__1_carry__5_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__1_carry__6 
       (.CI(\modmultiply/minusOp_inferred__1_carry__5_n_0 ),
        .CO({\modmultiply/minusOp_inferred__1_carry__6_n_0 ,\modmultiply/minusOp_inferred__1_carry__6_n_1 ,\modmultiply/minusOp_inferred__1_carry__6_n_2 ,\modmultiply/minusOp_inferred__1_carry__6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg1[31:28]),
        .O(minusOp0_in[31:28]),
        .S({minusOp_inferred__1_carry__6_i_1__0_n_0,minusOp_inferred__1_carry__6_i_2__0_n_0,minusOp_inferred__1_carry__6_i_3__0_n_0,minusOp_inferred__1_carry__6_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/minusOp_inferred__1_carry__7 
       (.CI(\modmultiply/minusOp_inferred__1_carry__6_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,prodreg1[32]}),
        .O({\modmultiply/minusOp_inferred__1_carry__7_n_4 ,\modmultiply/minusOp_inferred__1_carry__7_n_5 ,minusOp0_in[33:32]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,minusOp_inferred__1_carry__7_i_1_n_0,minusOp_inferred__1_carry__7_i_2__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[10] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[10]),
        .Q(modreg1[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[11] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[11]),
        .Q(modreg1[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[12] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[12]),
        .Q(modreg1[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[13] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[13]),
        .Q(modreg1[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[14] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[14]),
        .Q(modreg1[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[15] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[15]),
        .Q(modreg1[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[16] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[16]),
        .Q(modreg1[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[17] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[17]),
        .Q(modreg1[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[18] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[18]),
        .Q(modreg1[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[19] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[19]),
        .Q(modreg1[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[1] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[1]),
        .Q(modreg1[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[20] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[20]),
        .Q(modreg1[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[21] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[21]),
        .Q(modreg1[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[22] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[22]),
        .Q(modreg1[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[23] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[23]),
        .Q(modreg1[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[24] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[24]),
        .Q(modreg1[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[25] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[25]),
        .Q(modreg1[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[26] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[26]),
        .Q(modreg1[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[27] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[27]),
        .Q(modreg1[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[28] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[28]),
        .Q(modreg1[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[29] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[29]),
        .Q(modreg1[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[2] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[2]),
        .Q(modreg1[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[30] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[30]),
        .Q(modreg1[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[31] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[31]),
        .Q(modreg1[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[3] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[3]),
        .Q(modreg1[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[4] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[4]),
        .Q(modreg1[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[5] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[5]),
        .Q(modreg1[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[6] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[6]),
        .Q(modreg1[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[7] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[7]),
        .Q(modreg1[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[8] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[8]),
        .Q(modreg1[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg1_reg[9] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[9]),
        .Q(modreg1[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/modreg2_reg[1] 
       (.C(clk),
        .CE(\prodreg[33]_i_1_n_0 ),
        .D(modreg[0]),
        .Q(modreg2),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[0] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(mpreg),
        .Q(\modmultiply/mpreg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[10] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[10]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[11] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[11]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[12] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[12]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[13] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[13]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[14] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[14]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[15] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[15]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[16] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[16]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[17] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[17]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[18] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[18]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[19] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[19]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[1] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[1]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[20] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[20]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[21] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[21]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[22] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[22]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[23] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[23]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[24] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[24]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[25] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[25]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[26] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[26]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[27] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[27]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[28] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[28]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[29] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[29]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[2] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[2]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[30] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[30]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[31] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[31]_i_2__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[3] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[3]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[4] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[4]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[5] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[5]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[6] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[6]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[7] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[7]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[8] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[8]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/mpreg_reg[9] 
       (.C(clk),
        .CE(\modmultiply/mpreg0 ),
        .D(\mpreg[9]_i_1__0_n_0 ),
        .Q(\modmultiply/mpreg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/plusOp_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\modmultiply/plusOp_carry_n_0 ,\modmultiply/plusOp_carry_n_1 ,\modmultiply/plusOp_carry_n_2 ,\modmultiply/plusOp_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg[3:0]),
        .O(prodreg1[3:0]),
        .S({plusOp_carry_i_1__0_n_0,plusOp_carry_i_2__0_n_0,plusOp_carry_i_3__0_n_0,plusOp_carry_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/plusOp_carry__0 
       (.CI(\modmultiply/plusOp_carry_n_0 ),
        .CO({\modmultiply/plusOp_carry__0_n_0 ,\modmultiply/plusOp_carry__0_n_1 ,\modmultiply/plusOp_carry__0_n_2 ,\modmultiply/plusOp_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg[7:4]),
        .O(prodreg1[7:4]),
        .S({plusOp_carry__0_i_1__0_n_0,plusOp_carry__0_i_2__0_n_0,plusOp_carry__0_i_3__0_n_0,plusOp_carry__0_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/plusOp_carry__1 
       (.CI(\modmultiply/plusOp_carry__0_n_0 ),
        .CO({\modmultiply/plusOp_carry__1_n_0 ,\modmultiply/plusOp_carry__1_n_1 ,\modmultiply/plusOp_carry__1_n_2 ,\modmultiply/plusOp_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg[11:8]),
        .O(prodreg1[11:8]),
        .S({plusOp_carry__1_i_1__0_n_0,plusOp_carry__1_i_2__0_n_0,plusOp_carry__1_i_3__0_n_0,plusOp_carry__1_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/plusOp_carry__2 
       (.CI(\modmultiply/plusOp_carry__1_n_0 ),
        .CO({\modmultiply/plusOp_carry__2_n_0 ,\modmultiply/plusOp_carry__2_n_1 ,\modmultiply/plusOp_carry__2_n_2 ,\modmultiply/plusOp_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg[15:12]),
        .O(prodreg1[15:12]),
        .S({plusOp_carry__2_i_1__0_n_0,plusOp_carry__2_i_2__0_n_0,plusOp_carry__2_i_3__0_n_0,plusOp_carry__2_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/plusOp_carry__3 
       (.CI(\modmultiply/plusOp_carry__2_n_0 ),
        .CO({\modmultiply/plusOp_carry__3_n_0 ,\modmultiply/plusOp_carry__3_n_1 ,\modmultiply/plusOp_carry__3_n_2 ,\modmultiply/plusOp_carry__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg[19:16]),
        .O(prodreg1[19:16]),
        .S({plusOp_carry__3_i_1__0_n_0,plusOp_carry__3_i_2__0_n_0,plusOp_carry__3_i_3__0_n_0,plusOp_carry__3_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/plusOp_carry__4 
       (.CI(\modmultiply/plusOp_carry__3_n_0 ),
        .CO({\modmultiply/plusOp_carry__4_n_0 ,\modmultiply/plusOp_carry__4_n_1 ,\modmultiply/plusOp_carry__4_n_2 ,\modmultiply/plusOp_carry__4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg[23:20]),
        .O(prodreg1[23:20]),
        .S({plusOp_carry__4_i_1__0_n_0,plusOp_carry__4_i_2__0_n_0,plusOp_carry__4_i_3__0_n_0,plusOp_carry__4_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/plusOp_carry__5 
       (.CI(\modmultiply/plusOp_carry__4_n_0 ),
        .CO({\modmultiply/plusOp_carry__5_n_0 ,\modmultiply/plusOp_carry__5_n_1 ,\modmultiply/plusOp_carry__5_n_2 ,\modmultiply/plusOp_carry__5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg[27:24]),
        .O(prodreg1[27:24]),
        .S({plusOp_carry__5_i_1__0_n_0,plusOp_carry__5_i_2__0_n_0,plusOp_carry__5_i_3__0_n_0,plusOp_carry__5_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/plusOp_carry__6 
       (.CI(\modmultiply/plusOp_carry__5_n_0 ),
        .CO({\modmultiply/plusOp_carry__6_n_0 ,\modmultiply/plusOp_carry__6_n_1 ,\modmultiply/plusOp_carry__6_n_2 ,\modmultiply/plusOp_carry__6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(prodreg[31:28]),
        .O(prodreg1[31:28]),
        .S({plusOp_carry__6_i_1__0_n_0,plusOp_carry__6_i_2__0_n_0,plusOp_carry__6_i_3__0_n_0,plusOp_carry__6_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modmultiply/plusOp_carry__7 
       (.CI(\modmultiply/plusOp_carry__6_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,prodreg[32]}),
        .O({\modmultiply/plusOp_carry__7_n_4 ,\modmultiply/plusOp_carry__7_n_5 ,prodreg1[33:32]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,plusOp_carry__7_i_1__0_n_0,plusOp_carry__7_i_2__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[0] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[0]_i_1_n_0 ),
        .Q(prodreg[0]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[10] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[10]_i_1_n_0 ),
        .Q(prodreg[10]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[11] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[11]_i_1_n_0 ),
        .Q(prodreg[11]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[12] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[12]_i_1_n_0 ),
        .Q(prodreg[12]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[13] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[13]_i_1_n_0 ),
        .Q(prodreg[13]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[14] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[14]_i_1_n_0 ),
        .Q(prodreg[14]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[15] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[15]_i_1_n_0 ),
        .Q(prodreg[15]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[16] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[16]_i_1_n_0 ),
        .Q(prodreg[16]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[17] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[17]_i_1_n_0 ),
        .Q(prodreg[17]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[18] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[18]_i_1_n_0 ),
        .Q(prodreg[18]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[19] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[19]_i_1_n_0 ),
        .Q(prodreg[19]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[1] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[1]_i_1_n_0 ),
        .Q(prodreg[1]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[20] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[20]_i_1_n_0 ),
        .Q(prodreg[20]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[21] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[21]_i_1_n_0 ),
        .Q(prodreg[21]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[22] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[22]_i_1_n_0 ),
        .Q(prodreg[22]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[23] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[23]_i_1_n_0 ),
        .Q(prodreg[23]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[24] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[24]_i_1_n_0 ),
        .Q(prodreg[24]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[25] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[25]_i_1_n_0 ),
        .Q(prodreg[25]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[26] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[26]_i_1_n_0 ),
        .Q(prodreg[26]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[27] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[27]_i_1_n_0 ),
        .Q(prodreg[27]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[28] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[28]_i_1_n_0 ),
        .Q(prodreg[28]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[29] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[29]_i_1_n_0 ),
        .Q(prodreg[29]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[2] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[2]_i_1_n_0 ),
        .Q(prodreg[2]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[30] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[30]_i_1_n_0 ),
        .Q(prodreg[30]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[31] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[31]_i_2_n_0 ),
        .Q(prodreg[31]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[32] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\prodreg[32]_i_1__0_n_0 ),
        .Q(prodreg[32]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[33] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\prodreg[33]_i_3__0_n_0 ),
        .Q(prodreg[33]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[3] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[3]_i_1_n_0 ),
        .Q(prodreg[3]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[4] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[4]_i_1_n_0 ),
        .Q(prodreg[4]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[5] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[5]_i_1_n_0 ),
        .Q(prodreg[5]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[6] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[6]_i_1_n_0 ),
        .Q(prodreg[6]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[7] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[7]_i_1_n_0 ),
        .Q(prodreg[7]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[8] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[8]_i_1_n_0 ),
        .Q(prodreg[8]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modmultiply/prodreg_reg[9] 
       (.C(clk),
        .CE(\modmultiply/prodreg0 ),
        .D(\cypher[9]_i_1_n_0 ),
        .Q(prodreg[9]),
        .R(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \modreg[31]_i_1 
       (.I0(ready),
        .I1(ds),
        .O(\modreg[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[0] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[0]),
        .Q(modreg[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[10] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[10]),
        .Q(modreg[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[11] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[11]),
        .Q(modreg[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[12] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[12]),
        .Q(modreg[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[13] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[13]),
        .Q(modreg[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[14] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[14]),
        .Q(modreg[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[15] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[15]),
        .Q(modreg[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[16] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[16]),
        .Q(modreg[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[17] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[17]),
        .Q(modreg[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[18] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[18]),
        .Q(modreg[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[19] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[19]),
        .Q(modreg[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[1] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[1]),
        .Q(modreg[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[20] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[20]),
        .Q(modreg[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[21] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[21]),
        .Q(modreg[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[22] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[22]),
        .Q(modreg[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[23] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[23]),
        .Q(modreg[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[24] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[24]),
        .Q(modreg[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[25] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[25]),
        .Q(modreg[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[26] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[26]),
        .Q(modreg[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[27] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[27]),
        .Q(modreg[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[28] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[28]),
        .Q(modreg[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[29] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[29]),
        .Q(modreg[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[2] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[2]),
        .Q(modreg[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[30] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[30]),
        .Q(modreg[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[31] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[31]),
        .Q(modreg[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[3] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[3]),
        .Q(modreg[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[4] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[4]),
        .Q(modreg[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[5] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[5]),
        .Q(modreg[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[6] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[6]),
        .Q(modreg[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[7] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[7]),
        .Q(modreg[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[8] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[8]),
        .Q(modreg[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \modreg_reg[9] 
       (.C(clk),
        .CE(\modreg[31]_i_1_n_0 ),
        .CLR(reset),
        .D(inMod[9]),
        .Q(modreg[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \modsqr/first_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(first_i_1__0_n_0),
        .PRE(reset),
        .Q(sqrrdy));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[0] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[0]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[10] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[10]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[11] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[11]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[12] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[12]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[13] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[13]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[14] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[14]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[15] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[15]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[16] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[16]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[17] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[17]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[18] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[18]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[19] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[19]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[1] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[1]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[20] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[20]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[21] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[21]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[22] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[22]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[23] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[23]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[24] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[24]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[25] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[25]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[26] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[26]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[27] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[27]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[28] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[28]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[29] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[29]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[2] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[2]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[30] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[30]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[31] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[31]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[32] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[32]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[33] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[33]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[3] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[3]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[4] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[4]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[5] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[5]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[6] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[6]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[7] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[7]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[8] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[8]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mcreg_reg[9] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mcreg[9]_i_1_n_0 ),
        .Q(\modsqr/mcreg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\modsqr/minusOp_inferred__0_carry_n_0 ,\modsqr/minusOp_inferred__0_carry_n_1 ,\modsqr/minusOp_inferred__0_carry_n_2 ,\modsqr/minusOp_inferred__0_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\modsqr/plusOp_carry_n_4 ,\modsqr/plusOp_carry_n_5 ,\modsqr/plusOp_carry_n_6 ,\modsqr/plusOp_carry_n_7 }),
        .O({\modsqr/minusOp_inferred__0_carry_n_4 ,\modsqr/minusOp_inferred__0_carry_n_5 ,\modsqr/minusOp_inferred__0_carry_n_6 ,\modsqr/minusOp_inferred__0_carry_n_7 }),
        .S({minusOp_inferred__0_carry_i_1_n_0,minusOp_inferred__0_carry_i_2_n_0,minusOp_inferred__0_carry_i_3_n_0,minusOp_inferred__0_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__0_carry__0 
       (.CI(\modsqr/minusOp_inferred__0_carry_n_0 ),
        .CO({\modsqr/minusOp_inferred__0_carry__0_n_0 ,\modsqr/minusOp_inferred__0_carry__0_n_1 ,\modsqr/minusOp_inferred__0_carry__0_n_2 ,\modsqr/minusOp_inferred__0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__0_n_4 ,\modsqr/plusOp_carry__0_n_5 ,\modsqr/plusOp_carry__0_n_6 ,\modsqr/plusOp_carry__0_n_7 }),
        .O({\modsqr/minusOp_inferred__0_carry__0_n_4 ,\modsqr/minusOp_inferred__0_carry__0_n_5 ,\modsqr/minusOp_inferred__0_carry__0_n_6 ,\modsqr/minusOp_inferred__0_carry__0_n_7 }),
        .S({minusOp_inferred__0_carry__0_i_1_n_0,minusOp_inferred__0_carry__0_i_2_n_0,minusOp_inferred__0_carry__0_i_3_n_0,minusOp_inferred__0_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__0_carry__1 
       (.CI(\modsqr/minusOp_inferred__0_carry__0_n_0 ),
        .CO({\modsqr/minusOp_inferred__0_carry__1_n_0 ,\modsqr/minusOp_inferred__0_carry__1_n_1 ,\modsqr/minusOp_inferred__0_carry__1_n_2 ,\modsqr/minusOp_inferred__0_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__1_n_4 ,\modsqr/plusOp_carry__1_n_5 ,\modsqr/plusOp_carry__1_n_6 ,\modsqr/plusOp_carry__1_n_7 }),
        .O({\modsqr/minusOp_inferred__0_carry__1_n_4 ,\modsqr/minusOp_inferred__0_carry__1_n_5 ,\modsqr/minusOp_inferred__0_carry__1_n_6 ,\modsqr/minusOp_inferred__0_carry__1_n_7 }),
        .S({minusOp_inferred__0_carry__1_i_1_n_0,minusOp_inferred__0_carry__1_i_2_n_0,minusOp_inferred__0_carry__1_i_3_n_0,minusOp_inferred__0_carry__1_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__0_carry__2 
       (.CI(\modsqr/minusOp_inferred__0_carry__1_n_0 ),
        .CO({\modsqr/minusOp_inferred__0_carry__2_n_0 ,\modsqr/minusOp_inferred__0_carry__2_n_1 ,\modsqr/minusOp_inferred__0_carry__2_n_2 ,\modsqr/minusOp_inferred__0_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__2_n_4 ,\modsqr/plusOp_carry__2_n_5 ,\modsqr/plusOp_carry__2_n_6 ,\modsqr/plusOp_carry__2_n_7 }),
        .O({\modsqr/minusOp_inferred__0_carry__2_n_4 ,\modsqr/minusOp_inferred__0_carry__2_n_5 ,\modsqr/minusOp_inferred__0_carry__2_n_6 ,\modsqr/minusOp_inferred__0_carry__2_n_7 }),
        .S({minusOp_inferred__0_carry__2_i_1_n_0,minusOp_inferred__0_carry__2_i_2_n_0,minusOp_inferred__0_carry__2_i_3_n_0,minusOp_inferred__0_carry__2_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__0_carry__3 
       (.CI(\modsqr/minusOp_inferred__0_carry__2_n_0 ),
        .CO({\modsqr/minusOp_inferred__0_carry__3_n_0 ,\modsqr/minusOp_inferred__0_carry__3_n_1 ,\modsqr/minusOp_inferred__0_carry__3_n_2 ,\modsqr/minusOp_inferred__0_carry__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__3_n_4 ,\modsqr/plusOp_carry__3_n_5 ,\modsqr/plusOp_carry__3_n_6 ,\modsqr/plusOp_carry__3_n_7 }),
        .O({\modsqr/minusOp_inferred__0_carry__3_n_4 ,\modsqr/minusOp_inferred__0_carry__3_n_5 ,\modsqr/minusOp_inferred__0_carry__3_n_6 ,\modsqr/minusOp_inferred__0_carry__3_n_7 }),
        .S({minusOp_inferred__0_carry__3_i_1_n_0,minusOp_inferred__0_carry__3_i_2_n_0,minusOp_inferred__0_carry__3_i_3_n_0,minusOp_inferred__0_carry__3_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__0_carry__4 
       (.CI(\modsqr/minusOp_inferred__0_carry__3_n_0 ),
        .CO({\modsqr/minusOp_inferred__0_carry__4_n_0 ,\modsqr/minusOp_inferred__0_carry__4_n_1 ,\modsqr/minusOp_inferred__0_carry__4_n_2 ,\modsqr/minusOp_inferred__0_carry__4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__4_n_4 ,\modsqr/plusOp_carry__4_n_5 ,\modsqr/plusOp_carry__4_n_6 ,\modsqr/plusOp_carry__4_n_7 }),
        .O({\modsqr/minusOp_inferred__0_carry__4_n_4 ,\modsqr/minusOp_inferred__0_carry__4_n_5 ,\modsqr/minusOp_inferred__0_carry__4_n_6 ,\modsqr/minusOp_inferred__0_carry__4_n_7 }),
        .S({minusOp_inferred__0_carry__4_i_1_n_0,minusOp_inferred__0_carry__4_i_2_n_0,minusOp_inferred__0_carry__4_i_3_n_0,minusOp_inferred__0_carry__4_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__0_carry__5 
       (.CI(\modsqr/minusOp_inferred__0_carry__4_n_0 ),
        .CO({\modsqr/minusOp_inferred__0_carry__5_n_0 ,\modsqr/minusOp_inferred__0_carry__5_n_1 ,\modsqr/minusOp_inferred__0_carry__5_n_2 ,\modsqr/minusOp_inferred__0_carry__5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__5_n_4 ,\modsqr/plusOp_carry__5_n_5 ,\modsqr/plusOp_carry__5_n_6 ,\modsqr/plusOp_carry__5_n_7 }),
        .O({\modsqr/minusOp_inferred__0_carry__5_n_4 ,\modsqr/minusOp_inferred__0_carry__5_n_5 ,\modsqr/minusOp_inferred__0_carry__5_n_6 ,\modsqr/minusOp_inferred__0_carry__5_n_7 }),
        .S({minusOp_inferred__0_carry__5_i_1_n_0,minusOp_inferred__0_carry__5_i_2_n_0,minusOp_inferred__0_carry__5_i_3_n_0,minusOp_inferred__0_carry__5_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__0_carry__6 
       (.CI(\modsqr/minusOp_inferred__0_carry__5_n_0 ),
        .CO({\modsqr/minusOp_inferred__0_carry__6_n_0 ,\modsqr/minusOp_inferred__0_carry__6_n_1 ,\modsqr/minusOp_inferred__0_carry__6_n_2 ,\modsqr/minusOp_inferred__0_carry__6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__6_n_4 ,\modsqr/plusOp_carry__6_n_5 ,\modsqr/plusOp_carry__6_n_6 ,\modsqr/plusOp_carry__6_n_7 }),
        .O({\modsqr/minusOp_inferred__0_carry__6_n_4 ,\modsqr/minusOp_inferred__0_carry__6_n_5 ,\modsqr/minusOp_inferred__0_carry__6_n_6 ,\modsqr/minusOp_inferred__0_carry__6_n_7 }),
        .S({minusOp_inferred__0_carry__6_i_1_n_0,minusOp_inferred__0_carry__6_i_2_n_0,minusOp_inferred__0_carry__6_i_3_n_0,minusOp_inferred__0_carry__6_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__0_carry__7 
       (.CI(\modsqr/minusOp_inferred__0_carry__6_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\modsqr/plusOp_carry__7_n_7 }),
        .O({\modsqr/minusOp_inferred__0_carry__7_n_4 ,\modsqr/minusOp_inferred__0_carry__7_n_5 ,\modsqr/minusOp_inferred__0_carry__7_n_6 ,\modsqr/minusOp_inferred__0_carry__7_n_7 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,minusOp_inferred__0_carry__7_i_1_n_0,minusOp_inferred__0_carry__7_i_2_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\modsqr/minusOp_inferred__1_carry_n_0 ,\modsqr/minusOp_inferred__1_carry_n_1 ,\modsqr/minusOp_inferred__1_carry_n_2 ,\modsqr/minusOp_inferred__1_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\modsqr/plusOp_carry_n_4 ,\modsqr/plusOp_carry_n_5 ,\modsqr/plusOp_carry_n_6 ,\modsqr/plusOp_carry_n_7 }),
        .O({\modsqr/minusOp_inferred__1_carry_n_4 ,\modsqr/minusOp_inferred__1_carry_n_5 ,\modsqr/minusOp_inferred__1_carry_n_6 ,\modsqr/minusOp_inferred__1_carry_n_7 }),
        .S({minusOp_inferred__1_carry_i_1_n_0,minusOp_inferred__1_carry_i_2_n_0,minusOp_inferred__1_carry_i_3_n_0,minusOp_inferred__1_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__1_carry__0 
       (.CI(\modsqr/minusOp_inferred__1_carry_n_0 ),
        .CO({\modsqr/minusOp_inferred__1_carry__0_n_0 ,\modsqr/minusOp_inferred__1_carry__0_n_1 ,\modsqr/minusOp_inferred__1_carry__0_n_2 ,\modsqr/minusOp_inferred__1_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__0_n_4 ,\modsqr/plusOp_carry__0_n_5 ,\modsqr/plusOp_carry__0_n_6 ,\modsqr/plusOp_carry__0_n_7 }),
        .O({\modsqr/minusOp_inferred__1_carry__0_n_4 ,\modsqr/minusOp_inferred__1_carry__0_n_5 ,\modsqr/minusOp_inferred__1_carry__0_n_6 ,\modsqr/minusOp_inferred__1_carry__0_n_7 }),
        .S({minusOp_inferred__1_carry__0_i_1_n_0,minusOp_inferred__1_carry__0_i_2_n_0,minusOp_inferred__1_carry__0_i_3_n_0,minusOp_inferred__1_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__1_carry__1 
       (.CI(\modsqr/minusOp_inferred__1_carry__0_n_0 ),
        .CO({\modsqr/minusOp_inferred__1_carry__1_n_0 ,\modsqr/minusOp_inferred__1_carry__1_n_1 ,\modsqr/minusOp_inferred__1_carry__1_n_2 ,\modsqr/minusOp_inferred__1_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__1_n_4 ,\modsqr/plusOp_carry__1_n_5 ,\modsqr/plusOp_carry__1_n_6 ,\modsqr/plusOp_carry__1_n_7 }),
        .O({\modsqr/minusOp_inferred__1_carry__1_n_4 ,\modsqr/minusOp_inferred__1_carry__1_n_5 ,\modsqr/minusOp_inferred__1_carry__1_n_6 ,\modsqr/minusOp_inferred__1_carry__1_n_7 }),
        .S({minusOp_inferred__1_carry__1_i_1_n_0,minusOp_inferred__1_carry__1_i_2_n_0,minusOp_inferred__1_carry__1_i_3_n_0,minusOp_inferred__1_carry__1_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__1_carry__2 
       (.CI(\modsqr/minusOp_inferred__1_carry__1_n_0 ),
        .CO({\modsqr/minusOp_inferred__1_carry__2_n_0 ,\modsqr/minusOp_inferred__1_carry__2_n_1 ,\modsqr/minusOp_inferred__1_carry__2_n_2 ,\modsqr/minusOp_inferred__1_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__2_n_4 ,\modsqr/plusOp_carry__2_n_5 ,\modsqr/plusOp_carry__2_n_6 ,\modsqr/plusOp_carry__2_n_7 }),
        .O({\modsqr/minusOp_inferred__1_carry__2_n_4 ,\modsqr/minusOp_inferred__1_carry__2_n_5 ,\modsqr/minusOp_inferred__1_carry__2_n_6 ,\modsqr/minusOp_inferred__1_carry__2_n_7 }),
        .S({minusOp_inferred__1_carry__2_i_1_n_0,minusOp_inferred__1_carry__2_i_2_n_0,minusOp_inferred__1_carry__2_i_3_n_0,minusOp_inferred__1_carry__2_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__1_carry__3 
       (.CI(\modsqr/minusOp_inferred__1_carry__2_n_0 ),
        .CO({\modsqr/minusOp_inferred__1_carry__3_n_0 ,\modsqr/minusOp_inferred__1_carry__3_n_1 ,\modsqr/minusOp_inferred__1_carry__3_n_2 ,\modsqr/minusOp_inferred__1_carry__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__3_n_4 ,\modsqr/plusOp_carry__3_n_5 ,\modsqr/plusOp_carry__3_n_6 ,\modsqr/plusOp_carry__3_n_7 }),
        .O({\modsqr/minusOp_inferred__1_carry__3_n_4 ,\modsqr/minusOp_inferred__1_carry__3_n_5 ,\modsqr/minusOp_inferred__1_carry__3_n_6 ,\modsqr/minusOp_inferred__1_carry__3_n_7 }),
        .S({minusOp_inferred__1_carry__3_i_1_n_0,minusOp_inferred__1_carry__3_i_2_n_0,minusOp_inferred__1_carry__3_i_3_n_0,minusOp_inferred__1_carry__3_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__1_carry__4 
       (.CI(\modsqr/minusOp_inferred__1_carry__3_n_0 ),
        .CO({\modsqr/minusOp_inferred__1_carry__4_n_0 ,\modsqr/minusOp_inferred__1_carry__4_n_1 ,\modsqr/minusOp_inferred__1_carry__4_n_2 ,\modsqr/minusOp_inferred__1_carry__4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__4_n_4 ,\modsqr/plusOp_carry__4_n_5 ,\modsqr/plusOp_carry__4_n_6 ,\modsqr/plusOp_carry__4_n_7 }),
        .O({\modsqr/minusOp_inferred__1_carry__4_n_4 ,\modsqr/minusOp_inferred__1_carry__4_n_5 ,\modsqr/minusOp_inferred__1_carry__4_n_6 ,\modsqr/minusOp_inferred__1_carry__4_n_7 }),
        .S({minusOp_inferred__1_carry__4_i_1_n_0,minusOp_inferred__1_carry__4_i_2_n_0,minusOp_inferred__1_carry__4_i_3_n_0,minusOp_inferred__1_carry__4_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__1_carry__5 
       (.CI(\modsqr/minusOp_inferred__1_carry__4_n_0 ),
        .CO({\modsqr/minusOp_inferred__1_carry__5_n_0 ,\modsqr/minusOp_inferred__1_carry__5_n_1 ,\modsqr/minusOp_inferred__1_carry__5_n_2 ,\modsqr/minusOp_inferred__1_carry__5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__5_n_4 ,\modsqr/plusOp_carry__5_n_5 ,\modsqr/plusOp_carry__5_n_6 ,\modsqr/plusOp_carry__5_n_7 }),
        .O({\modsqr/minusOp_inferred__1_carry__5_n_4 ,\modsqr/minusOp_inferred__1_carry__5_n_5 ,\modsqr/minusOp_inferred__1_carry__5_n_6 ,\modsqr/minusOp_inferred__1_carry__5_n_7 }),
        .S({minusOp_inferred__1_carry__5_i_1_n_0,minusOp_inferred__1_carry__5_i_2_n_0,minusOp_inferred__1_carry__5_i_3_n_0,minusOp_inferred__1_carry__5_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__1_carry__6 
       (.CI(\modsqr/minusOp_inferred__1_carry__5_n_0 ),
        .CO({\modsqr/minusOp_inferred__1_carry__6_n_0 ,\modsqr/minusOp_inferred__1_carry__6_n_1 ,\modsqr/minusOp_inferred__1_carry__6_n_2 ,\modsqr/minusOp_inferred__1_carry__6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/plusOp_carry__6_n_4 ,\modsqr/plusOp_carry__6_n_5 ,\modsqr/plusOp_carry__6_n_6 ,\modsqr/plusOp_carry__6_n_7 }),
        .O({\modsqr/minusOp_inferred__1_carry__6_n_4 ,\modsqr/minusOp_inferred__1_carry__6_n_5 ,\modsqr/minusOp_inferred__1_carry__6_n_6 ,\modsqr/minusOp_inferred__1_carry__6_n_7 }),
        .S({minusOp_inferred__1_carry__6_i_1_n_0,minusOp_inferred__1_carry__6_i_2_n_0,minusOp_inferred__1_carry__6_i_3_n_0,minusOp_inferred__1_carry__6_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/minusOp_inferred__1_carry__7 
       (.CI(\modsqr/minusOp_inferred__1_carry__6_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\modsqr/plusOp_carry__7_n_7 }),
        .O({\modsqr/minusOp_inferred__1_carry__7_n_4 ,\modsqr/minusOp_inferred__1_carry__7_n_5 ,\modsqr/minusOp_inferred__1_carry__7_n_6 ,\modsqr/minusOp_inferred__1_carry__7_n_7 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,minusOp_inferred__1_carry__7_i_1__0_n_0,minusOp_inferred__1_carry__7_i_2_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[10] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[10]),
        .Q(\modsqr/modreg1_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[11] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[11]),
        .Q(\modsqr/modreg1_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[12] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[12]),
        .Q(\modsqr/modreg1_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[13] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[13]),
        .Q(\modsqr/modreg1_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[14] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[14]),
        .Q(\modsqr/modreg1_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[15] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[15]),
        .Q(\modsqr/modreg1_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[16] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[16]),
        .Q(\modsqr/modreg1_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[17] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[17]),
        .Q(\modsqr/modreg1_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[18] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[18]),
        .Q(\modsqr/modreg1_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[19] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[19]),
        .Q(\modsqr/modreg1_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[1] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[1]),
        .Q(\modsqr/modreg1_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[20] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[20]),
        .Q(\modsqr/modreg1_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[21] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[21]),
        .Q(\modsqr/modreg1_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[22] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[22]),
        .Q(\modsqr/modreg1_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[23] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[23]),
        .Q(\modsqr/modreg1_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[24] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[24]),
        .Q(\modsqr/modreg1_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[25] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[25]),
        .Q(\modsqr/modreg1_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[26] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[26]),
        .Q(\modsqr/modreg1_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[27] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[27]),
        .Q(\modsqr/modreg1_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[28] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[28]),
        .Q(\modsqr/modreg1_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[29] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[29]),
        .Q(\modsqr/modreg1_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[2] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[2]),
        .Q(\modsqr/modreg1_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[30] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[30]),
        .Q(\modsqr/modreg1_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[31] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[31]),
        .Q(\modsqr/modreg1_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[3] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[3]),
        .Q(\modsqr/modreg1_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[4] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[4]),
        .Q(\modsqr/modreg1_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[5] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[5]),
        .Q(\modsqr/modreg1_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[6] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[6]),
        .Q(\modsqr/modreg1_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[7] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[7]),
        .Q(\modsqr/modreg1_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[8] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[8]),
        .Q(\modsqr/modreg1_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg1_reg[9] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[9]),
        .Q(\modsqr/modreg1_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/modreg2_reg[1] 
       (.C(clk),
        .CE(\prodreg[33]_i_1__0_n_0 ),
        .D(modreg[0]),
        .Q(\modsqr/modreg2_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[0] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[0]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[10] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[10]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[11] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[11]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[12] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[12]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[13] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[13]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[14] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[14]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[15] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[15]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[16] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[16]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[17] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[17]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[18] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[18]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[19] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[19]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[1] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[1]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[20] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[20]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[21] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[21]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[22] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[22]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[23] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[23]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[24] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[24]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[25] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[25]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[26] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[26]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[27] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[27]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[28] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[28]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[29] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[29]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[2] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[2]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[30] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[30]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[31] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[31]_i_2_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[3] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[3]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[4] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[4]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[5] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[5]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[6] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[6]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[7] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[7]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[8] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[8]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/mpreg_reg[9] 
       (.C(clk),
        .CE(\modsqr/mpreg0 ),
        .D(\mpreg[9]_i_1_n_0 ),
        .Q(\modsqr/mpreg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/plusOp_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\modsqr/plusOp_carry_n_0 ,\modsqr/plusOp_carry_n_1 ,\modsqr/plusOp_carry_n_2 ,\modsqr/plusOp_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/prodreg_reg_n_0_[3] ,\modsqr/prodreg_reg_n_0_[2] ,\modsqr/prodreg_reg_n_0_[1] ,\modsqr/prodreg_reg_n_0_ }),
        .O({\modsqr/plusOp_carry_n_4 ,\modsqr/plusOp_carry_n_5 ,\modsqr/plusOp_carry_n_6 ,\modsqr/plusOp_carry_n_7 }),
        .S({plusOp_carry_i_1_n_0,plusOp_carry_i_2_n_0,plusOp_carry_i_3_n_0,plusOp_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/plusOp_carry__0 
       (.CI(\modsqr/plusOp_carry_n_0 ),
        .CO({\modsqr/plusOp_carry__0_n_0 ,\modsqr/plusOp_carry__0_n_1 ,\modsqr/plusOp_carry__0_n_2 ,\modsqr/plusOp_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/prodreg_reg_n_0_[7] ,\modsqr/prodreg_reg_n_0_[6] ,\modsqr/prodreg_reg_n_0_[5] ,\modsqr/prodreg_reg_n_0_[4] }),
        .O({\modsqr/plusOp_carry__0_n_4 ,\modsqr/plusOp_carry__0_n_5 ,\modsqr/plusOp_carry__0_n_6 ,\modsqr/plusOp_carry__0_n_7 }),
        .S({plusOp_carry__0_i_1_n_0,plusOp_carry__0_i_2_n_0,plusOp_carry__0_i_3_n_0,plusOp_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/plusOp_carry__1 
       (.CI(\modsqr/plusOp_carry__0_n_0 ),
        .CO({\modsqr/plusOp_carry__1_n_0 ,\modsqr/plusOp_carry__1_n_1 ,\modsqr/plusOp_carry__1_n_2 ,\modsqr/plusOp_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/prodreg_reg_n_0_[11] ,\modsqr/prodreg_reg_n_0_[10] ,\modsqr/prodreg_reg_n_0_[9] ,\modsqr/prodreg_reg_n_0_[8] }),
        .O({\modsqr/plusOp_carry__1_n_4 ,\modsqr/plusOp_carry__1_n_5 ,\modsqr/plusOp_carry__1_n_6 ,\modsqr/plusOp_carry__1_n_7 }),
        .S({plusOp_carry__1_i_1_n_0,plusOp_carry__1_i_2_n_0,plusOp_carry__1_i_3_n_0,plusOp_carry__1_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/plusOp_carry__2 
       (.CI(\modsqr/plusOp_carry__1_n_0 ),
        .CO({\modsqr/plusOp_carry__2_n_0 ,\modsqr/plusOp_carry__2_n_1 ,\modsqr/plusOp_carry__2_n_2 ,\modsqr/plusOp_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/prodreg_reg_n_0_[15] ,\modsqr/prodreg_reg_n_0_[14] ,\modsqr/prodreg_reg_n_0_[13] ,\modsqr/prodreg_reg_n_0_[12] }),
        .O({\modsqr/plusOp_carry__2_n_4 ,\modsqr/plusOp_carry__2_n_5 ,\modsqr/plusOp_carry__2_n_6 ,\modsqr/plusOp_carry__2_n_7 }),
        .S({plusOp_carry__2_i_1_n_0,plusOp_carry__2_i_2_n_0,plusOp_carry__2_i_3_n_0,plusOp_carry__2_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/plusOp_carry__3 
       (.CI(\modsqr/plusOp_carry__2_n_0 ),
        .CO({\modsqr/plusOp_carry__3_n_0 ,\modsqr/plusOp_carry__3_n_1 ,\modsqr/plusOp_carry__3_n_2 ,\modsqr/plusOp_carry__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/prodreg_reg_n_0_[19] ,\modsqr/prodreg_reg_n_0_[18] ,\modsqr/prodreg_reg_n_0_[17] ,\modsqr/prodreg_reg_n_0_[16] }),
        .O({\modsqr/plusOp_carry__3_n_4 ,\modsqr/plusOp_carry__3_n_5 ,\modsqr/plusOp_carry__3_n_6 ,\modsqr/plusOp_carry__3_n_7 }),
        .S({plusOp_carry__3_i_1_n_0,plusOp_carry__3_i_2_n_0,plusOp_carry__3_i_3_n_0,plusOp_carry__3_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/plusOp_carry__4 
       (.CI(\modsqr/plusOp_carry__3_n_0 ),
        .CO({\modsqr/plusOp_carry__4_n_0 ,\modsqr/plusOp_carry__4_n_1 ,\modsqr/plusOp_carry__4_n_2 ,\modsqr/plusOp_carry__4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/prodreg_reg_n_0_[23] ,\modsqr/prodreg_reg_n_0_[22] ,\modsqr/prodreg_reg_n_0_[21] ,\modsqr/prodreg_reg_n_0_[20] }),
        .O({\modsqr/plusOp_carry__4_n_4 ,\modsqr/plusOp_carry__4_n_5 ,\modsqr/plusOp_carry__4_n_6 ,\modsqr/plusOp_carry__4_n_7 }),
        .S({plusOp_carry__4_i_1_n_0,plusOp_carry__4_i_2_n_0,plusOp_carry__4_i_3_n_0,plusOp_carry__4_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/plusOp_carry__5 
       (.CI(\modsqr/plusOp_carry__4_n_0 ),
        .CO({\modsqr/plusOp_carry__5_n_0 ,\modsqr/plusOp_carry__5_n_1 ,\modsqr/plusOp_carry__5_n_2 ,\modsqr/plusOp_carry__5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/prodreg_reg_n_0_[27] ,\modsqr/prodreg_reg_n_0_[26] ,\modsqr/prodreg_reg_n_0_[25] ,\modsqr/prodreg_reg_n_0_[24] }),
        .O({\modsqr/plusOp_carry__5_n_4 ,\modsqr/plusOp_carry__5_n_5 ,\modsqr/plusOp_carry__5_n_6 ,\modsqr/plusOp_carry__5_n_7 }),
        .S({plusOp_carry__5_i_1_n_0,plusOp_carry__5_i_2_n_0,plusOp_carry__5_i_3_n_0,plusOp_carry__5_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/plusOp_carry__6 
       (.CI(\modsqr/plusOp_carry__5_n_0 ),
        .CO({\modsqr/plusOp_carry__6_n_0 ,\modsqr/plusOp_carry__6_n_1 ,\modsqr/plusOp_carry__6_n_2 ,\modsqr/plusOp_carry__6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\modsqr/prodreg_reg_n_0_[31] ,\modsqr/prodreg_reg_n_0_[30] ,\modsqr/prodreg_reg_n_0_[29] ,\modsqr/prodreg_reg_n_0_[28] }),
        .O({\modsqr/plusOp_carry__6_n_4 ,\modsqr/plusOp_carry__6_n_5 ,\modsqr/plusOp_carry__6_n_6 ,\modsqr/plusOp_carry__6_n_7 }),
        .S({plusOp_carry__6_i_1_n_0,plusOp_carry__6_i_2_n_0,plusOp_carry__6_i_3_n_0,plusOp_carry__6_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \modsqr/plusOp_carry__7 
       (.CI(\modsqr/plusOp_carry__6_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\modsqr/prodreg_reg_n_0_[32] }),
        .O({\modsqr/plusOp_carry__7_n_4 ,\modsqr/plusOp_carry__7_n_5 ,\modsqr/plusOp_carry__7_n_6 ,\modsqr/plusOp_carry__7_n_7 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,plusOp_carry__7_i_1_n_0,plusOp_carry__7_i_2_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[0] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[0]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_ ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[10] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[10]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[10] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[11] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[11]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[11] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[12] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[12]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[12] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[13] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[13]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[13] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[14] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[14]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[14] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[15] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[15]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[15] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[16] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[16]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[16] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[17] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[17]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[17] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[18] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[18]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[18] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[19] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[19]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[19] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[1] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[1]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[1] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[20] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[20]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[20] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[21] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[21]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[21] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[22] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[22]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[22] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[23] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[23]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[23] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[24] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[24]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[24] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[25] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[25]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[25] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[26] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[26]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[26] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[27] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[27]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[27] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[28] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[28]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[28] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[29] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[29]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[29] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[2] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[2]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[2] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[30] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[30]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[30] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[31] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[31]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[31] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[32] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[32]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[32] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[33] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[33]_i_3_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[33] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[3] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[3]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[3] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[4] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[4]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[4] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[5] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[5]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[5] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[6] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[6]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[6] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[7] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[7]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[7] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[8] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[8]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[8] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \modsqr/prodreg_reg[9] 
       (.C(clk),
        .CE(\modsqr/prodreg0 ),
        .D(\prodreg[9]_i_1_n_0 ),
        .Q(\modsqr/prodreg_reg_n_0_[9] ),
        .R(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[0]_i_1 
       (.I0(root[0]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[1] ),
        .O(\mpreg[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[0]_i_1__0 
       (.I0(sqrin_reg_n_0_),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[1] ),
        .O(mpreg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[10]_i_1 
       (.I0(root[10]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[11] ),
        .O(\mpreg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[10]_i_1__0 
       (.I0(\sqrin_reg_n_0_[10] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[11] ),
        .O(\mpreg[10]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[11]_i_1 
       (.I0(root[11]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[12] ),
        .O(\mpreg[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[11]_i_1__0 
       (.I0(\sqrin_reg_n_0_[11] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[12] ),
        .O(\mpreg[11]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[12]_i_1 
       (.I0(root[12]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[13] ),
        .O(\mpreg[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[12]_i_1__0 
       (.I0(\sqrin_reg_n_0_[12] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[13] ),
        .O(\mpreg[12]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[13]_i_1 
       (.I0(root[13]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[14] ),
        .O(\mpreg[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[13]_i_1__0 
       (.I0(\sqrin_reg_n_0_[13] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[14] ),
        .O(\mpreg[13]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[14]_i_1 
       (.I0(root[14]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[15] ),
        .O(\mpreg[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[14]_i_1__0 
       (.I0(\sqrin_reg_n_0_[14] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[15] ),
        .O(\mpreg[14]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[15]_i_1 
       (.I0(root[15]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[16] ),
        .O(\mpreg[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[15]_i_1__0 
       (.I0(\sqrin_reg_n_0_[15] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[16] ),
        .O(\mpreg[15]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[16]_i_1 
       (.I0(root[16]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[17] ),
        .O(\mpreg[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[16]_i_1__0 
       (.I0(\sqrin_reg_n_0_[16] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[17] ),
        .O(\mpreg[16]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[17]_i_1 
       (.I0(root[17]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[18] ),
        .O(\mpreg[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[17]_i_1__0 
       (.I0(\sqrin_reg_n_0_[17] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[18] ),
        .O(\mpreg[17]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[18]_i_1 
       (.I0(root[18]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[19] ),
        .O(\mpreg[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[18]_i_1__0 
       (.I0(\sqrin_reg_n_0_[18] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[19] ),
        .O(\mpreg[18]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[19]_i_1 
       (.I0(root[19]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[20] ),
        .O(\mpreg[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[19]_i_1__0 
       (.I0(\sqrin_reg_n_0_[19] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[20] ),
        .O(\mpreg[19]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[1]_i_1 
       (.I0(root[1]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[2] ),
        .O(\mpreg[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[1]_i_1__0 
       (.I0(\sqrin_reg_n_0_[1] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[2] ),
        .O(\mpreg[1]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[20]_i_1 
       (.I0(root[20]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[21] ),
        .O(\mpreg[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[20]_i_1__0 
       (.I0(\sqrin_reg_n_0_[20] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[21] ),
        .O(\mpreg[20]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[21]_i_1 
       (.I0(root[21]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[22] ),
        .O(\mpreg[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[21]_i_1__0 
       (.I0(\sqrin_reg_n_0_[21] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[22] ),
        .O(\mpreg[21]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[22]_i_1 
       (.I0(root[22]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[23] ),
        .O(\mpreg[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[22]_i_1__0 
       (.I0(\sqrin_reg_n_0_[22] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[23] ),
        .O(\mpreg[22]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[23]_i_1 
       (.I0(root[23]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[24] ),
        .O(\mpreg[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[23]_i_1__0 
       (.I0(\sqrin_reg_n_0_[23] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[24] ),
        .O(\mpreg[23]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[24]_i_1 
       (.I0(root[24]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[25] ),
        .O(\mpreg[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[24]_i_1__0 
       (.I0(\sqrin_reg_n_0_[24] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[25] ),
        .O(\mpreg[24]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[25]_i_1 
       (.I0(root[25]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[26] ),
        .O(\mpreg[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[25]_i_1__0 
       (.I0(\sqrin_reg_n_0_[25] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[26] ),
        .O(\mpreg[25]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[26]_i_1 
       (.I0(root[26]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[27] ),
        .O(\mpreg[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[26]_i_1__0 
       (.I0(\sqrin_reg_n_0_[26] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[27] ),
        .O(\mpreg[26]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[27]_i_1 
       (.I0(root[27]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[28] ),
        .O(\mpreg[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[27]_i_1__0 
       (.I0(\sqrin_reg_n_0_[27] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[28] ),
        .O(\mpreg[27]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[28]_i_1 
       (.I0(root[28]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[29] ),
        .O(\mpreg[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[28]_i_1__0 
       (.I0(\sqrin_reg_n_0_[28] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[29] ),
        .O(\mpreg[28]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[29]_i_1 
       (.I0(root[29]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[30] ),
        .O(\mpreg[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[29]_i_1__0 
       (.I0(\sqrin_reg_n_0_[29] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[30] ),
        .O(\mpreg[29]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[2]_i_1 
       (.I0(root[2]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[3] ),
        .O(\mpreg[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[2]_i_1__0 
       (.I0(\sqrin_reg_n_0_[2] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[3] ),
        .O(\mpreg[2]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[30]_i_1 
       (.I0(root[30]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[31] ),
        .O(\mpreg[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[30]_i_1__0 
       (.I0(\sqrin_reg_n_0_[30] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[31] ),
        .O(\mpreg[30]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \mpreg[31]_i_1 
       (.I0(\mpreg[31]_i_3_n_0 ),
        .I1(multrdy),
        .I2(multgo_reg_n_0),
        .I3(reset),
        .O(\modmultiply/mpreg0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \mpreg[31]_i_10 
       (.I0(\modmultiply/mpreg_reg_n_0_[31] ),
        .I1(\modmultiply/mpreg_reg_n_0_[28] ),
        .I2(\modmultiply/mpreg_reg_n_0_[30] ),
        .I3(\modmultiply/mpreg_reg_n_0_[29] ),
        .O(\mpreg[31]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \mpreg[31]_i_10__0 
       (.I0(\modsqr/mpreg_reg_n_0_[31] ),
        .I1(\modsqr/mpreg_reg_n_0_[28] ),
        .I2(\modsqr/mpreg_reg_n_0_[30] ),
        .I3(\modsqr/mpreg_reg_n_0_[29] ),
        .O(\mpreg[31]_i_10__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \mpreg[31]_i_11 
       (.I0(\modmultiply/mpreg_reg_n_0_[2] ),
        .I1(\modmultiply/mpreg_reg_n_0_[1] ),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .I3(\modmultiply/mpreg_reg_n_0_[3] ),
        .O(\mpreg[31]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \mpreg[31]_i_11__0 
       (.I0(\modsqr/mpreg_reg_n_0_[2] ),
        .I1(\modsqr/mpreg_reg_n_0_[1] ),
        .I2(\modsqr/mpreg_reg_n_0_ ),
        .I3(\modsqr/mpreg_reg_n_0_[3] ),
        .O(\mpreg[31]_i_11__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00CA)) 
    \mpreg[31]_i_1__0 
       (.I0(\mpreg[31]_i_3__0_n_0 ),
        .I1(multgo_reg_n_0),
        .I2(sqrrdy),
        .I3(reset),
        .O(\modsqr/mpreg0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \mpreg[31]_i_2 
       (.I0(sqrrdy),
        .I1(root[31]),
        .O(\mpreg[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \mpreg[31]_i_2__0 
       (.I0(multrdy),
        .I1(\sqrin_reg_n_0_[31] ),
        .O(\mpreg[31]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFEFF)) 
    \mpreg[31]_i_3 
       (.I0(\mpreg[31]_i_4_n_0 ),
        .I1(\mpreg[31]_i_5_n_0 ),
        .I2(\mpreg[31]_i_6_n_0 ),
        .I3(\mpreg[31]_i_7_n_0 ),
        .O(\mpreg[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFEFF)) 
    \mpreg[31]_i_3__0 
       (.I0(\mpreg[31]_i_4__0_n_0 ),
        .I1(\mpreg[31]_i_5__0_n_0 ),
        .I2(\mpreg[31]_i_6__0_n_0 ),
        .I3(\mpreg[31]_i_7__0_n_0 ),
        .O(\mpreg[31]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \mpreg[31]_i_4 
       (.I0(\modmultiply/mpreg_reg_n_0_[17] ),
        .I1(\modmultiply/mpreg_reg_n_0_[18] ),
        .I2(\modmultiply/mpreg_reg_n_0_[16] ),
        .I3(\modmultiply/mpreg_reg_n_0_[19] ),
        .I4(\mpreg[31]_i_8_n_0 ),
        .O(\mpreg[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \mpreg[31]_i_4__0 
       (.I0(\modsqr/mpreg_reg_n_0_[17] ),
        .I1(\modsqr/mpreg_reg_n_0_[18] ),
        .I2(\modsqr/mpreg_reg_n_0_[16] ),
        .I3(\modsqr/mpreg_reg_n_0_[19] ),
        .I4(\mpreg[31]_i_8__0_n_0 ),
        .O(\mpreg[31]_i_4__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \mpreg[31]_i_5 
       (.I0(\modmultiply/mpreg_reg_n_0_[9] ),
        .I1(\modmultiply/mpreg_reg_n_0_[10] ),
        .I2(\modmultiply/mpreg_reg_n_0_[8] ),
        .I3(\modmultiply/mpreg_reg_n_0_[11] ),
        .I4(\mpreg[31]_i_9_n_0 ),
        .O(\mpreg[31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \mpreg[31]_i_5__0 
       (.I0(\modsqr/mpreg_reg_n_0_[9] ),
        .I1(\modsqr/mpreg_reg_n_0_[10] ),
        .I2(\modsqr/mpreg_reg_n_0_[8] ),
        .I3(\modsqr/mpreg_reg_n_0_[11] ),
        .I4(\mpreg[31]_i_9__0_n_0 ),
        .O(\mpreg[31]_i_5__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \mpreg[31]_i_6 
       (.I0(\modmultiply/mpreg_reg_n_0_[5] ),
        .I1(\modmultiply/mpreg_reg_n_0_[6] ),
        .I2(\modmultiply/mpreg_reg_n_0_[4] ),
        .I3(\modmultiply/mpreg_reg_n_0_[7] ),
        .I4(\mpreg[31]_i_10_n_0 ),
        .O(\mpreg[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \mpreg[31]_i_6__0 
       (.I0(\modsqr/mpreg_reg_n_0_[5] ),
        .I1(\modsqr/mpreg_reg_n_0_[6] ),
        .I2(\modsqr/mpreg_reg_n_0_[4] ),
        .I3(\modsqr/mpreg_reg_n_0_[7] ),
        .I4(\mpreg[31]_i_10__0_n_0 ),
        .O(\mpreg[31]_i_6__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \mpreg[31]_i_7 
       (.I0(\modmultiply/mpreg_reg_n_0_[25] ),
        .I1(\modmultiply/mpreg_reg_n_0_[26] ),
        .I2(\modmultiply/mpreg_reg_n_0_[24] ),
        .I3(\modmultiply/mpreg_reg_n_0_[27] ),
        .I4(\mpreg[31]_i_11_n_0 ),
        .O(\mpreg[31]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \mpreg[31]_i_7__0 
       (.I0(\modsqr/mpreg_reg_n_0_[25] ),
        .I1(\modsqr/mpreg_reg_n_0_[26] ),
        .I2(\modsqr/mpreg_reg_n_0_[24] ),
        .I3(\modsqr/mpreg_reg_n_0_[27] ),
        .I4(\mpreg[31]_i_11__0_n_0 ),
        .O(\mpreg[31]_i_7__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \mpreg[31]_i_8 
       (.I0(\modmultiply/mpreg_reg_n_0_[15] ),
        .I1(\modmultiply/mpreg_reg_n_0_[12] ),
        .I2(\modmultiply/mpreg_reg_n_0_[14] ),
        .I3(\modmultiply/mpreg_reg_n_0_[13] ),
        .O(\mpreg[31]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \mpreg[31]_i_8__0 
       (.I0(\modsqr/mpreg_reg_n_0_[15] ),
        .I1(\modsqr/mpreg_reg_n_0_[12] ),
        .I2(\modsqr/mpreg_reg_n_0_[14] ),
        .I3(\modsqr/mpreg_reg_n_0_[13] ),
        .O(\mpreg[31]_i_8__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \mpreg[31]_i_9 
       (.I0(\modmultiply/mpreg_reg_n_0_[23] ),
        .I1(\modmultiply/mpreg_reg_n_0_[20] ),
        .I2(\modmultiply/mpreg_reg_n_0_[22] ),
        .I3(\modmultiply/mpreg_reg_n_0_[21] ),
        .O(\mpreg[31]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \mpreg[31]_i_9__0 
       (.I0(\modsqr/mpreg_reg_n_0_[23] ),
        .I1(\modsqr/mpreg_reg_n_0_[20] ),
        .I2(\modsqr/mpreg_reg_n_0_[22] ),
        .I3(\modsqr/mpreg_reg_n_0_[21] ),
        .O(\mpreg[31]_i_9__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[3]_i_1 
       (.I0(root[3]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[4] ),
        .O(\mpreg[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[3]_i_1__0 
       (.I0(\sqrin_reg_n_0_[3] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[4] ),
        .O(\mpreg[3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[4]_i_1 
       (.I0(root[4]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[5] ),
        .O(\mpreg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[4]_i_1__0 
       (.I0(\sqrin_reg_n_0_[4] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[5] ),
        .O(\mpreg[4]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[5]_i_1 
       (.I0(root[5]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[6] ),
        .O(\mpreg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[5]_i_1__0 
       (.I0(\sqrin_reg_n_0_[5] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[6] ),
        .O(\mpreg[5]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[6]_i_1 
       (.I0(root[6]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[7] ),
        .O(\mpreg[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[6]_i_1__0 
       (.I0(\sqrin_reg_n_0_[6] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[7] ),
        .O(\mpreg[6]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[7]_i_1 
       (.I0(root[7]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[8] ),
        .O(\mpreg[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[7]_i_1__0 
       (.I0(\sqrin_reg_n_0_[7] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[8] ),
        .O(\mpreg[7]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[8]_i_1 
       (.I0(root[8]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[9] ),
        .O(\mpreg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[8]_i_1__0 
       (.I0(\sqrin_reg_n_0_[8] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[9] ),
        .O(\mpreg[8]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[9]_i_1 
       (.I0(root[9]),
        .I1(sqrrdy),
        .I2(\modsqr/mpreg_reg_n_0_[10] ),
        .O(\mpreg[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \mpreg[9]_i_1__0 
       (.I0(\sqrin_reg_n_0_[9] ),
        .I1(multrdy),
        .I2(\modmultiply/mpreg_reg_n_0_[10] ),
        .O(\mpreg[9]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FF0D0D0D)) 
    multgo_i_1
       (.I0(\cypher[31]_i_3_n_0 ),
        .I1(multgo_i_2_n_0),
        .I2(multgo_i_3_n_0),
        .I3(ready),
        .I4(ds),
        .I5(multgo_reg_n_0),
        .O(multgo_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    multgo_i_2
       (.I0(\cypher[31]_i_11_n_0 ),
        .I1(\count_reg_n_0_[7] ),
        .I2(\count_reg_n_0_[4] ),
        .I3(\count_reg_n_0_[6] ),
        .I4(\count_reg_n_0_[5] ),
        .I5(\cypher[31]_i_4_n_0 ),
        .O(multgo_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    multgo_i_3
       (.I0(ready),
        .I1(sqrrdy),
        .I2(multrdy),
        .O(multgo_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    multgo_reg
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(reset),
        .D(multgo_i_1_n_0),
        .Q(multgo_reg_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__0_i_1
       (.I0(\modsqr/prodreg_reg_n_0_[7] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[7] ),
        .O(plusOp_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__0_i_1__0
       (.I0(prodreg[7]),
        .I1(mcreg[7]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__0_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__0_i_2
       (.I0(\modsqr/prodreg_reg_n_0_[6] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[6] ),
        .O(plusOp_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__0_i_2__0
       (.I0(prodreg[6]),
        .I1(mcreg[6]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__0_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__0_i_3
       (.I0(\modsqr/prodreg_reg_n_0_[5] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[5] ),
        .O(plusOp_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__0_i_3__0
       (.I0(prodreg[5]),
        .I1(mcreg[5]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__0_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__0_i_4
       (.I0(\modsqr/prodreg_reg_n_0_[4] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[4] ),
        .O(plusOp_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__0_i_4__0
       (.I0(prodreg[4]),
        .I1(mcreg[4]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__0_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__1_i_1
       (.I0(\modsqr/prodreg_reg_n_0_[11] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[11] ),
        .O(plusOp_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__1_i_1__0
       (.I0(prodreg[11]),
        .I1(mcreg[11]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__1_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__1_i_2
       (.I0(\modsqr/prodreg_reg_n_0_[10] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[10] ),
        .O(plusOp_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__1_i_2__0
       (.I0(prodreg[10]),
        .I1(mcreg[10]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__1_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__1_i_3
       (.I0(\modsqr/prodreg_reg_n_0_[9] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[9] ),
        .O(plusOp_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__1_i_3__0
       (.I0(prodreg[9]),
        .I1(mcreg[9]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__1_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__1_i_4
       (.I0(\modsqr/prodreg_reg_n_0_[8] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[8] ),
        .O(plusOp_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__1_i_4__0
       (.I0(prodreg[8]),
        .I1(mcreg[8]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__1_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__2_i_1
       (.I0(\modsqr/prodreg_reg_n_0_[15] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[15] ),
        .O(plusOp_carry__2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__2_i_1__0
       (.I0(prodreg[15]),
        .I1(mcreg[15]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__2_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__2_i_2
       (.I0(\modsqr/prodreg_reg_n_0_[14] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[14] ),
        .O(plusOp_carry__2_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__2_i_2__0
       (.I0(prodreg[14]),
        .I1(mcreg[14]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__2_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__2_i_3
       (.I0(\modsqr/prodreg_reg_n_0_[13] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[13] ),
        .O(plusOp_carry__2_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__2_i_3__0
       (.I0(prodreg[13]),
        .I1(mcreg[13]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__2_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__2_i_4
       (.I0(\modsqr/prodreg_reg_n_0_[12] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[12] ),
        .O(plusOp_carry__2_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__2_i_4__0
       (.I0(prodreg[12]),
        .I1(mcreg[12]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__2_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__3_i_1
       (.I0(\modsqr/prodreg_reg_n_0_[19] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[19] ),
        .O(plusOp_carry__3_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__3_i_1__0
       (.I0(prodreg[19]),
        .I1(mcreg[19]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__3_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__3_i_2
       (.I0(\modsqr/prodreg_reg_n_0_[18] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[18] ),
        .O(plusOp_carry__3_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__3_i_2__0
       (.I0(prodreg[18]),
        .I1(mcreg[18]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__3_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__3_i_3
       (.I0(\modsqr/prodreg_reg_n_0_[17] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[17] ),
        .O(plusOp_carry__3_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__3_i_3__0
       (.I0(prodreg[17]),
        .I1(mcreg[17]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__3_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__3_i_4
       (.I0(\modsqr/prodreg_reg_n_0_[16] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[16] ),
        .O(plusOp_carry__3_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__3_i_4__0
       (.I0(prodreg[16]),
        .I1(mcreg[16]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__3_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__4_i_1
       (.I0(\modsqr/prodreg_reg_n_0_[23] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[23] ),
        .O(plusOp_carry__4_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__4_i_1__0
       (.I0(prodreg[23]),
        .I1(mcreg[23]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__4_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__4_i_2
       (.I0(\modsqr/prodreg_reg_n_0_[22] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[22] ),
        .O(plusOp_carry__4_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__4_i_2__0
       (.I0(prodreg[22]),
        .I1(mcreg[22]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__4_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__4_i_3
       (.I0(\modsqr/prodreg_reg_n_0_[21] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[21] ),
        .O(plusOp_carry__4_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__4_i_3__0
       (.I0(prodreg[21]),
        .I1(mcreg[21]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__4_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__4_i_4
       (.I0(\modsqr/prodreg_reg_n_0_[20] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[20] ),
        .O(plusOp_carry__4_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__4_i_4__0
       (.I0(prodreg[20]),
        .I1(mcreg[20]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__4_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__5_i_1
       (.I0(\modsqr/prodreg_reg_n_0_[27] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[27] ),
        .O(plusOp_carry__5_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__5_i_1__0
       (.I0(prodreg[27]),
        .I1(mcreg[27]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__5_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__5_i_2
       (.I0(\modsqr/prodreg_reg_n_0_[26] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[26] ),
        .O(plusOp_carry__5_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__5_i_2__0
       (.I0(prodreg[26]),
        .I1(mcreg[26]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__5_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__5_i_3
       (.I0(\modsqr/prodreg_reg_n_0_[25] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[25] ),
        .O(plusOp_carry__5_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__5_i_3__0
       (.I0(prodreg[25]),
        .I1(mcreg[25]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__5_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__5_i_4
       (.I0(\modsqr/prodreg_reg_n_0_[24] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[24] ),
        .O(plusOp_carry__5_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__5_i_4__0
       (.I0(prodreg[24]),
        .I1(mcreg[24]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__5_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__6_i_1
       (.I0(\modsqr/prodreg_reg_n_0_[31] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[31] ),
        .O(plusOp_carry__6_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__6_i_1__0
       (.I0(prodreg[31]),
        .I1(mcreg[31]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__6_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__6_i_2
       (.I0(\modsqr/prodreg_reg_n_0_[30] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[30] ),
        .O(plusOp_carry__6_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__6_i_2__0
       (.I0(prodreg[30]),
        .I1(mcreg[30]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__6_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__6_i_3
       (.I0(\modsqr/prodreg_reg_n_0_[29] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[29] ),
        .O(plusOp_carry__6_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__6_i_3__0
       (.I0(prodreg[29]),
        .I1(mcreg[29]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__6_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__6_i_4
       (.I0(\modsqr/prodreg_reg_n_0_[28] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[28] ),
        .O(plusOp_carry__6_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__6_i_4__0
       (.I0(prodreg[28]),
        .I1(mcreg[28]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__6_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__7_i_1
       (.I0(\modsqr/prodreg_reg_n_0_[33] ),
        .I1(\modsqr/mcreg_reg_n_0_[33] ),
        .I2(\modsqr/mpreg_reg_n_0_ ),
        .O(plusOp_carry__7_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__7_i_1__0
       (.I0(prodreg[33]),
        .I1(mcreg[33]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry__7_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__7_i_2
       (.I0(\modsqr/prodreg_reg_n_0_[32] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[32] ),
        .O(plusOp_carry__7_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry__7_i_2__0
       (.I0(prodreg[32]),
        .I1(\modmultiply/mpreg_reg_n_0_ ),
        .I2(mcreg[32]),
        .O(plusOp_carry__7_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry_i_1
       (.I0(\modsqr/prodreg_reg_n_0_[3] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[3] ),
        .O(plusOp_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry_i_1__0
       (.I0(prodreg[3]),
        .I1(mcreg[3]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry_i_2
       (.I0(\modsqr/prodreg_reg_n_0_[2] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[2] ),
        .O(plusOp_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry_i_2__0
       (.I0(prodreg[2]),
        .I1(mcreg[2]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry_i_3
       (.I0(\modsqr/prodreg_reg_n_0_[1] ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_[1] ),
        .O(plusOp_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry_i_3__0
       (.I0(prodreg[1]),
        .I1(mcreg[1]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry_i_4
       (.I0(\modsqr/prodreg_reg_n_0_ ),
        .I1(\modsqr/mpreg_reg_n_0_ ),
        .I2(\modsqr/mcreg_reg_n_0_ ),
        .O(plusOp_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6A)) 
    plusOp_carry_i_4__0
       (.I0(prodreg[0]),
        .I1(mcreg[0]),
        .I2(\modmultiply/mpreg_reg_n_0_ ),
        .O(plusOp_carry_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[0]_i_1 
       (.I0(\modsqr/plusOp_carry_n_7 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry_n_7 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry_n_7 ),
        .O(\prodreg[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[10]_i_1 
       (.I0(\modsqr/plusOp_carry__1_n_5 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__1_n_5 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__1_n_5 ),
        .O(\prodreg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[11]_i_1 
       (.I0(\modsqr/plusOp_carry__1_n_4 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__1_n_4 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__1_n_4 ),
        .O(\prodreg[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[12]_i_1 
       (.I0(\modsqr/plusOp_carry__2_n_7 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__2_n_7 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__2_n_7 ),
        .O(\prodreg[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[13]_i_1 
       (.I0(\modsqr/plusOp_carry__2_n_6 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__2_n_6 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__2_n_6 ),
        .O(\prodreg[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[14]_i_1 
       (.I0(\modsqr/plusOp_carry__2_n_5 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__2_n_5 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__2_n_5 ),
        .O(\prodreg[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[15]_i_1 
       (.I0(\modsqr/plusOp_carry__2_n_4 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__2_n_4 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__2_n_4 ),
        .O(\prodreg[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[16]_i_1 
       (.I0(\modsqr/plusOp_carry__3_n_7 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__3_n_7 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__3_n_7 ),
        .O(\prodreg[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[17]_i_1 
       (.I0(\modsqr/plusOp_carry__3_n_6 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__3_n_6 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__3_n_6 ),
        .O(\prodreg[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[18]_i_1 
       (.I0(\modsqr/plusOp_carry__3_n_5 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__3_n_5 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__3_n_5 ),
        .O(\prodreg[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[19]_i_1 
       (.I0(\modsqr/plusOp_carry__3_n_4 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__3_n_4 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__3_n_4 ),
        .O(\prodreg[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[1]_i_1 
       (.I0(\modsqr/plusOp_carry_n_6 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry_n_6 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry_n_6 ),
        .O(\prodreg[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[20]_i_1 
       (.I0(\modsqr/plusOp_carry__4_n_7 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__4_n_7 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__4_n_7 ),
        .O(\prodreg[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[21]_i_1 
       (.I0(\modsqr/plusOp_carry__4_n_6 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__4_n_6 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__4_n_6 ),
        .O(\prodreg[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[22]_i_1 
       (.I0(\modsqr/plusOp_carry__4_n_5 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__4_n_5 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__4_n_5 ),
        .O(\prodreg[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[23]_i_1 
       (.I0(\modsqr/plusOp_carry__4_n_4 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__4_n_4 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__4_n_4 ),
        .O(\prodreg[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[24]_i_1 
       (.I0(\modsqr/plusOp_carry__5_n_7 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__5_n_7 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__5_n_7 ),
        .O(\prodreg[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[25]_i_1 
       (.I0(\modsqr/plusOp_carry__5_n_6 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__5_n_6 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__5_n_6 ),
        .O(\prodreg[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[26]_i_1 
       (.I0(\modsqr/plusOp_carry__5_n_5 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__5_n_5 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__5_n_5 ),
        .O(\prodreg[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[27]_i_1 
       (.I0(\modsqr/plusOp_carry__5_n_4 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__5_n_4 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__5_n_4 ),
        .O(\prodreg[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[28]_i_1 
       (.I0(\modsqr/plusOp_carry__6_n_7 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__6_n_7 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__6_n_7 ),
        .O(\prodreg[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[29]_i_1 
       (.I0(\modsqr/plusOp_carry__6_n_6 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__6_n_6 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__6_n_6 ),
        .O(\prodreg[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[2]_i_1 
       (.I0(\modsqr/plusOp_carry_n_5 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry_n_5 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry_n_5 ),
        .O(\prodreg[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[30]_i_1 
       (.I0(\modsqr/plusOp_carry__6_n_5 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__6_n_5 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__6_n_5 ),
        .O(\prodreg[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[31]_i_1 
       (.I0(\modsqr/plusOp_carry__6_n_4 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__6_n_4 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__6_n_4 ),
        .O(\prodreg[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[32]_i_1 
       (.I0(\modsqr/plusOp_carry__7_n_7 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__7_n_7 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__7_n_7 ),
        .O(\prodreg[32]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[32]_i_1__0 
       (.I0(prodreg1[32]),
        .I1(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modmultiply/minusOp_inferred__0_carry__7_n_7 ),
        .I3(minusOp0_in[33]),
        .I4(minusOp0_in[32]),
        .O(\prodreg[32]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \prodreg[33]_i_1 
       (.I0(reset),
        .I1(multgo_reg_n_0),
        .I2(multrdy),
        .O(\prodreg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \prodreg[33]_i_1__0 
       (.I0(reset),
        .I1(sqrrdy),
        .I2(multgo_reg_n_0),
        .O(\prodreg[33]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \prodreg[33]_i_2 
       (.I0(\mpreg[31]_i_3_n_0 ),
        .I1(reset),
        .I2(multrdy),
        .O(\modmultiply/prodreg0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \prodreg[33]_i_2__0 
       (.I0(\mpreg[31]_i_3__0_n_0 ),
        .I1(reset),
        .I2(sqrrdy),
        .O(\modsqr/prodreg0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \prodreg[33]_i_3 
       (.I0(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I1(\modsqr/plusOp_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .O(\prodreg[33]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \prodreg[33]_i_3__0 
       (.I0(\modmultiply/minusOp_inferred__0_carry__7_n_6 ),
        .I1(prodreg1[33]),
        .I2(minusOp0_in[33]),
        .O(\prodreg[33]_i_3__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[3]_i_1 
       (.I0(\modsqr/plusOp_carry_n_4 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry_n_4 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry_n_4 ),
        .O(\prodreg[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[4]_i_1 
       (.I0(\modsqr/plusOp_carry__0_n_7 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__0_n_7 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__0_n_7 ),
        .O(\prodreg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[5]_i_1 
       (.I0(\modsqr/plusOp_carry__0_n_6 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__0_n_6 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__0_n_6 ),
        .O(\prodreg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[6]_i_1 
       (.I0(\modsqr/plusOp_carry__0_n_5 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__0_n_5 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__0_n_5 ),
        .O(\prodreg[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[7]_i_1 
       (.I0(\modsqr/plusOp_carry__0_n_4 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__0_n_4 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__0_n_4 ),
        .O(\prodreg[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[8]_i_1 
       (.I0(\modsqr/plusOp_carry__1_n_7 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__1_n_7 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__1_n_7 ),
        .O(\prodreg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \prodreg[9]_i_1 
       (.I0(\modsqr/plusOp_carry__1_n_6 ),
        .I1(\modsqr/minusOp_inferred__0_carry__7_n_6 ),
        .I2(\modsqr/minusOp_inferred__0_carry__1_n_6 ),
        .I3(\modsqr/minusOp_inferred__1_carry__7_n_6 ),
        .I4(\modsqr/minusOp_inferred__1_carry__1_n_6 ),
        .O(\prodreg[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[0]_i_1 
       (.I0(indata[0]),
        .I1(ready),
        .I2(\prodreg[0]_i_1_n_0 ),
        .O(\root[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[10]_i_1 
       (.I0(indata[10]),
        .I1(ready),
        .I2(\prodreg[10]_i_1_n_0 ),
        .O(\root[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[11]_i_1 
       (.I0(indata[11]),
        .I1(ready),
        .I2(\prodreg[11]_i_1_n_0 ),
        .O(\root[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[12]_i_1 
       (.I0(indata[12]),
        .I1(ready),
        .I2(\prodreg[12]_i_1_n_0 ),
        .O(\root[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[13]_i_1 
       (.I0(indata[13]),
        .I1(ready),
        .I2(\prodreg[13]_i_1_n_0 ),
        .O(\root[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[14]_i_1 
       (.I0(indata[14]),
        .I1(ready),
        .I2(\prodreg[14]_i_1_n_0 ),
        .O(\root[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[15]_i_1 
       (.I0(indata[15]),
        .I1(ready),
        .I2(\prodreg[15]_i_1_n_0 ),
        .O(\root[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[16]_i_1 
       (.I0(indata[16]),
        .I1(ready),
        .I2(\prodreg[16]_i_1_n_0 ),
        .O(\root[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[17]_i_1 
       (.I0(indata[17]),
        .I1(ready),
        .I2(\prodreg[17]_i_1_n_0 ),
        .O(\root[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[18]_i_1 
       (.I0(indata[18]),
        .I1(ready),
        .I2(\prodreg[18]_i_1_n_0 ),
        .O(\root[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[19]_i_1 
       (.I0(indata[19]),
        .I1(ready),
        .I2(\prodreg[19]_i_1_n_0 ),
        .O(\root[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[1]_i_1 
       (.I0(indata[1]),
        .I1(ready),
        .I2(\prodreg[1]_i_1_n_0 ),
        .O(\root[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[20]_i_1 
       (.I0(indata[20]),
        .I1(ready),
        .I2(\prodreg[20]_i_1_n_0 ),
        .O(\root[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[21]_i_1 
       (.I0(indata[21]),
        .I1(ready),
        .I2(\prodreg[21]_i_1_n_0 ),
        .O(\root[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[22]_i_1 
       (.I0(indata[22]),
        .I1(ready),
        .I2(\prodreg[22]_i_1_n_0 ),
        .O(\root[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[23]_i_1 
       (.I0(indata[23]),
        .I1(ready),
        .I2(\prodreg[23]_i_1_n_0 ),
        .O(\root[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[24]_i_1 
       (.I0(indata[24]),
        .I1(ready),
        .I2(\prodreg[24]_i_1_n_0 ),
        .O(\root[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[25]_i_1 
       (.I0(indata[25]),
        .I1(ready),
        .I2(\prodreg[25]_i_1_n_0 ),
        .O(\root[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[26]_i_1 
       (.I0(indata[26]),
        .I1(ready),
        .I2(\prodreg[26]_i_1_n_0 ),
        .O(\root[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[27]_i_1 
       (.I0(indata[27]),
        .I1(ready),
        .I2(\prodreg[27]_i_1_n_0 ),
        .O(\root[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[28]_i_1 
       (.I0(indata[28]),
        .I1(ready),
        .I2(\prodreg[28]_i_1_n_0 ),
        .O(\root[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[29]_i_1 
       (.I0(indata[29]),
        .I1(ready),
        .I2(\prodreg[29]_i_1_n_0 ),
        .O(\root[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[2]_i_1 
       (.I0(indata[2]),
        .I1(ready),
        .I2(\prodreg[2]_i_1_n_0 ),
        .O(\root[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[30]_i_1 
       (.I0(indata[30]),
        .I1(ready),
        .I2(\prodreg[30]_i_1_n_0 ),
        .O(\root[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \root[31]_i_1 
       (.I0(ds),
        .I1(ready),
        .O(sqrin));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[31]_i_2 
       (.I0(indata[31]),
        .I1(ready),
        .I2(\prodreg[31]_i_1_n_0 ),
        .O(\root[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[3]_i_1 
       (.I0(indata[3]),
        .I1(ready),
        .I2(\prodreg[3]_i_1_n_0 ),
        .O(\root[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[4]_i_1 
       (.I0(indata[4]),
        .I1(ready),
        .I2(\prodreg[4]_i_1_n_0 ),
        .O(\root[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[5]_i_1 
       (.I0(indata[5]),
        .I1(ready),
        .I2(\prodreg[5]_i_1_n_0 ),
        .O(\root[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[6]_i_1 
       (.I0(indata[6]),
        .I1(ready),
        .I2(\prodreg[6]_i_1_n_0 ),
        .O(\root[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[7]_i_1 
       (.I0(indata[7]),
        .I1(ready),
        .I2(\prodreg[7]_i_1_n_0 ),
        .O(\root[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[8]_i_1 
       (.I0(indata[8]),
        .I1(ready),
        .I2(\prodreg[8]_i_1_n_0 ),
        .O(\root[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \root[9]_i_1 
       (.I0(indata[9]),
        .I1(ready),
        .I2(\prodreg[9]_i_1_n_0 ),
        .O(\root[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[0] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[0]_i_1_n_0 ),
        .Q(root[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[10] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[10]_i_1_n_0 ),
        .Q(root[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[11] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[11]_i_1_n_0 ),
        .Q(root[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[12] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[12]_i_1_n_0 ),
        .Q(root[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[13] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[13]_i_1_n_0 ),
        .Q(root[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[14] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[14]_i_1_n_0 ),
        .Q(root[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[15] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[15]_i_1_n_0 ),
        .Q(root[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[16] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[16]_i_1_n_0 ),
        .Q(root[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[17] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[17]_i_1_n_0 ),
        .Q(root[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[18] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[18]_i_1_n_0 ),
        .Q(root[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[19] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[19]_i_1_n_0 ),
        .Q(root[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[1] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[1]_i_1_n_0 ),
        .Q(root[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[20] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[20]_i_1_n_0 ),
        .Q(root[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[21] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[21]_i_1_n_0 ),
        .Q(root[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[22] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[22]_i_1_n_0 ),
        .Q(root[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[23] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[23]_i_1_n_0 ),
        .Q(root[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[24] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[24]_i_1_n_0 ),
        .Q(root[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[25] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[25]_i_1_n_0 ),
        .Q(root[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[26] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[26]_i_1_n_0 ),
        .Q(root[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[27] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[27]_i_1_n_0 ),
        .Q(root[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[28] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[28]_i_1_n_0 ),
        .Q(root[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[29] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[29]_i_1_n_0 ),
        .Q(root[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[2] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[2]_i_1_n_0 ),
        .Q(root[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[30] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[30]_i_1_n_0 ),
        .Q(root[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[31] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[31]_i_2_n_0 ),
        .Q(root[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[3] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[3]_i_1_n_0 ),
        .Q(root[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[4] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[4]_i_1_n_0 ),
        .Q(root[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[5] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[5]_i_1_n_0 ),
        .Q(root[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[6] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[6]_i_1_n_0 ),
        .Q(root[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[7] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[7]_i_1_n_0 ),
        .Q(root[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[8] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[8]_i_1_n_0 ),
        .Q(root[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \root_reg[9] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\root[9]_i_1_n_0 ),
        .Q(root[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    \sqrin[0]_i_1 
       (.I0(\prodreg[0]_i_1_n_0 ),
        .I1(count_reg_n_0_),
        .I2(ready),
        .O(\sqrin[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[10]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[10]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[11]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[11]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[12]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[12]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[13]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[13]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[14]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[14]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[15]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[15]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[16]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[16]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[17]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[17]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[18]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[18]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[19]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[19]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[1]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[1]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[20]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[20]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[21]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[21]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[22]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[22]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[23]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[23]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[24]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[24]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[25]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[25]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[26]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[26]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[27]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[27]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[28]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[28]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[29]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[29]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[2]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[2]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[30]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[30]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[31]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[31]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[3]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[3]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[4]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[4]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[5]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[5]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[6]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[6]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[7]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[7]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[8]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[8]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sqrin[9]_i_1 
       (.I0(count_reg_n_0_),
        .I1(\prodreg[9]_i_1_n_0 ),
        .I2(ready),
        .O(\sqrin[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[0] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[0]_i_1_n_0 ),
        .Q(sqrin_reg_n_0_));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[10] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[10]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[11] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[11]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[12] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[12]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[12] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[13] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[13]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[13] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[14] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[14]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[14] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[15] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[15]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[15] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[16] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[16]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[16] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[17] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[17]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[17] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[18] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[18]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[18] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[19] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[19]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[19] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[1] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[1]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[20] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[20]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[20] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[21] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[21]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[21] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[22] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[22]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[22] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[23] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[23]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[23] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[24] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[24]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[24] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[25] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[25]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[25] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[26] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[26]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[26] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[27] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[27]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[27] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[28] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[28]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[28] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[29] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[29]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[29] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[2] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[2]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[30] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[30]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[30] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[31] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[31]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[31] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[3] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[3]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[4] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[4]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[5] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[5]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[6] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[6]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[7] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[7]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[8] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[8]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sqrin_reg[9] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\sqrin[9]_i_1_n_0 ),
        .Q(\sqrin_reg_n_0_[9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT4 #(
    .INIT(16'hBFB0)) 
    \tempin[0]_i_1 
       (.I0(indata[0]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[0]_i_1_n_0 ),
        .O(\tempin[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[10]_i_1 
       (.I0(indata[10]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[10]_i_1_n_0 ),
        .O(\tempin[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[11]_i_1 
       (.I0(indata[11]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[11]_i_1_n_0 ),
        .O(\tempin[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[12]_i_1 
       (.I0(indata[12]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[12]_i_1_n_0 ),
        .O(\tempin[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[13]_i_1 
       (.I0(indata[13]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[13]_i_1_n_0 ),
        .O(\tempin[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[14]_i_1 
       (.I0(indata[14]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[14]_i_1_n_0 ),
        .O(\tempin[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[15]_i_1 
       (.I0(indata[15]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[15]_i_1_n_0 ),
        .O(\tempin[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[16]_i_1 
       (.I0(indata[16]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[16]_i_1_n_0 ),
        .O(\tempin[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[17]_i_1 
       (.I0(indata[17]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[17]_i_1_n_0 ),
        .O(\tempin[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[18]_i_1 
       (.I0(indata[18]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[18]_i_1_n_0 ),
        .O(\tempin[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[19]_i_1 
       (.I0(indata[19]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[19]_i_1_n_0 ),
        .O(\tempin[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[1]_i_1 
       (.I0(indata[1]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[1]_i_1_n_0 ),
        .O(\tempin[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[20]_i_1 
       (.I0(indata[20]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[20]_i_1_n_0 ),
        .O(\tempin[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[21]_i_1 
       (.I0(indata[21]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[21]_i_1_n_0 ),
        .O(\tempin[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[22]_i_1 
       (.I0(indata[22]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[22]_i_1_n_0 ),
        .O(\tempin[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[23]_i_1 
       (.I0(indata[23]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[23]_i_1_n_0 ),
        .O(\tempin[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[24]_i_1 
       (.I0(indata[24]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[24]_i_1_n_0 ),
        .O(\tempin[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[25]_i_1 
       (.I0(indata[25]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[25]_i_1_n_0 ),
        .O(\tempin[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[26]_i_1 
       (.I0(indata[26]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[26]_i_1_n_0 ),
        .O(\tempin[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[27]_i_1 
       (.I0(indata[27]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[27]_i_1_n_0 ),
        .O(\tempin[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[28]_i_1 
       (.I0(indata[28]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[28]_i_1_n_0 ),
        .O(\tempin[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[29]_i_1 
       (.I0(indata[29]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[29]_i_1_n_0 ),
        .O(\tempin[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[2]_i_1 
       (.I0(indata[2]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[2]_i_1_n_0 ),
        .O(\tempin[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[30]_i_1 
       (.I0(indata[30]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[30]_i_1_n_0 ),
        .O(\tempin[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[31]_i_1 
       (.I0(indata[31]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[31]_i_2_n_0 ),
        .O(\tempin[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[3]_i_1 
       (.I0(indata[3]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[3]_i_1_n_0 ),
        .O(\tempin[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[4]_i_1 
       (.I0(indata[4]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[4]_i_1_n_0 ),
        .O(\tempin[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[5]_i_1 
       (.I0(indata[5]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[5]_i_1_n_0 ),
        .O(\tempin[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[6]_i_1 
       (.I0(indata[6]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[6]_i_1_n_0 ),
        .O(\tempin[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[7]_i_1 
       (.I0(indata[7]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[7]_i_1_n_0 ),
        .O(\tempin[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[8]_i_1 
       (.I0(indata[8]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[8]_i_1_n_0 ),
        .O(\tempin[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT4 #(
    .INIT(16'h8F80)) 
    \tempin[9]_i_1 
       (.I0(indata[9]),
        .I1(inExp[0]),
        .I2(ready),
        .I3(\cypher[9]_i_1_n_0 ),
        .O(\tempin[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[0] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[0]_i_1_n_0 ),
        .Q(tempin[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[10] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[10]_i_1_n_0 ),
        .Q(tempin[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[11] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[11]_i_1_n_0 ),
        .Q(tempin[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[12] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[12]_i_1_n_0 ),
        .Q(tempin[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[13] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[13]_i_1_n_0 ),
        .Q(tempin[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[14] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[14]_i_1_n_0 ),
        .Q(tempin[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[15] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[15]_i_1_n_0 ),
        .Q(tempin[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[16] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[16]_i_1_n_0 ),
        .Q(tempin[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[17] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[17]_i_1_n_0 ),
        .Q(tempin[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[18] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[18]_i_1_n_0 ),
        .Q(tempin[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[19] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[19]_i_1_n_0 ),
        .Q(tempin[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[1] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[1]_i_1_n_0 ),
        .Q(tempin[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[20] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[20]_i_1_n_0 ),
        .Q(tempin[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[21] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[21]_i_1_n_0 ),
        .Q(tempin[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[22] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[22]_i_1_n_0 ),
        .Q(tempin[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[23] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[23]_i_1_n_0 ),
        .Q(tempin[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[24] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[24]_i_1_n_0 ),
        .Q(tempin[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[25] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[25]_i_1_n_0 ),
        .Q(tempin[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[26] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[26]_i_1_n_0 ),
        .Q(tempin[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[27] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[27]_i_1_n_0 ),
        .Q(tempin[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[28] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[28]_i_1_n_0 ),
        .Q(tempin[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[29] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[29]_i_1_n_0 ),
        .Q(tempin[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[2] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[2]_i_1_n_0 ),
        .Q(tempin[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[30] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[30]_i_1_n_0 ),
        .Q(tempin[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[31] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[31]_i_1_n_0 ),
        .Q(tempin[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[3] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[3]_i_1_n_0 ),
        .Q(tempin[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[4] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[4]_i_1_n_0 ),
        .Q(tempin[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[5] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[5]_i_1_n_0 ),
        .Q(tempin[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[6] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[6]_i_1_n_0 ),
        .Q(tempin[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[7] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[7]_i_1_n_0 ),
        .Q(tempin[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[8] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[8]_i_1_n_0 ),
        .Q(tempin[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \tempin_reg[9] 
       (.C(clk),
        .CE(sqrin),
        .CLR(reset),
        .D(\tempin[9]_i_1_n_0 ),
        .Q(tempin[9]));
endmodule
