module des3_perf
   (desOut,
    desIn,
    key1,
    key2,
    key3,
    decrypt,
    backdoor,
    clk);
  output backdoor;
  output [63:0]desOut;
  input [63:0]desIn;
  input [55:0]key1;
  input [55:0]key2;
  input [55:0]key3;
  input decrypt;
  input clk;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire decrypt;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]desIn;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]desOut;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]key1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]key2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]key3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]key_a;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire key_b_r_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][10]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][11]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][12]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][13]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][14]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][15]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][16]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][17]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][18]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][19]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][1]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][20]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][21]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][22]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][23]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][24]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][25]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][26]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][27]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][28]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][29]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][2]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][30]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][31]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][32]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][33]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][34]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][35]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][36]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][37]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][38]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][39]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][3]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][40]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][41]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][42]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][43]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][44]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][45]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][46]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][47]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][48]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][49]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][4]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][50]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][51]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][52]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][53]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][54]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][55]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][5]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][6]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][7]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][8]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg[16][9]_srl16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire key_b_r_reg_n_0_;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_b_r_reg_n_0_[0][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]key_c;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire key_c_r_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][10]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][11]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][12]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][13]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][14]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][15]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][16]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][17]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][18]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][19]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][1]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][20]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][21]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][22]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][23]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][24]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][25]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][26]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][27]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][28]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][29]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][2]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][30]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][31]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][32]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][33]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][34]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][35]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][36]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][37]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][38]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][39]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][3]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][40]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][41]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][42]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][43]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][44]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][45]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][46]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][47]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][48]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][49]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][4]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][50]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][51]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][52]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][53]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][54]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][55]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][5]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][6]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][7]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][8]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[31][9]_srl32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][0]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][10]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][11]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][12]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][13]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][14]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][15]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][16]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][17]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][18]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][19]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][1]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][20]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][21]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][22]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][23]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][24]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][25]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][26]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][27]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][28]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][29]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][2]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][30]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][31]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][32]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][33]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][34]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][35]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][36]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][37]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][38]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][39]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][3]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][40]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][41]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][42]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][43]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][44]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][45]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][46]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][47]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][48]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][49]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][4]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][50]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][51]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][52]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][53]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][54]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][55]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][5]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][6]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][7]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][8]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \key_c_r_reg[33][9]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]stage1_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]stage2_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:64]\u0/FP ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:64]\u0/IP ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L14 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/L9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R00 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/R10_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R30 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R40 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R50 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/R9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u0/R90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u0/key_r ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out14 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out15 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u0/out9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u0/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u1/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u10/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u11/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u12/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u13/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u14/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u15/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u2/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u3/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u4/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u5/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u6/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u7/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u8/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u0/u9/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r0_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u0/uk/K_r1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u0/uk/K_r10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u0/uk/K_r11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u0/uk/K_r12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u0/uk/K_r13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r14_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u0/uk/K_r2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u0/uk/K_r3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r4_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u0/uk/K_r5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r6_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/K_r7_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u0/uk/K_r8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u0/uk/K_r9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_10_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_11_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_12_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_13_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_14_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_15_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_16_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_17_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_18_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_19_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_20_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_21_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_22_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_23_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_24_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_25_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_26_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_27_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_28_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_29_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_2_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_30_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_31_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_32_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_33_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_34_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_35_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_36_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_37_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_38_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_39_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_3_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_40_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_41_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_42_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_43_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_44_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_45_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_47_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_48_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_49_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_4_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_50_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_51_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_52_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_53_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_5_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_6_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_7_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_8_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u0/uk/p_9_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:64]\u1/FP ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:64]\u1/IP ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L14 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/L9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R00 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/R10_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R30 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R40 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R50 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/R9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u1/R90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u1/key_r ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out14 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out15 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u1/out9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u0/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u1/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u10/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u11/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u12/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u13/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u14/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u15/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u2/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u3/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u4/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u5/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u6/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u7/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u8/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u1/u9/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r0_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u1/uk/K_r1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u1/uk/K_r10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u1/uk/K_r11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u1/uk/K_r12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u1/uk/K_r13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r14_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u1/uk/K_r2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u1/uk/K_r3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r4_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u1/uk/K_r5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r6_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/K_r7_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u1/uk/K_r8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u1/uk/K_r9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_10_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_11_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_12_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_13_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_14_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_15_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_16_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_17_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_18_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_19_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_20_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_21_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_22_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_23_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_24_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_25_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_26_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_27_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_28_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_29_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_2_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_30_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_31_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_32_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_33_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_34_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_35_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_36_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_37_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_38_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_39_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_3_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_40_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_41_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_42_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_43_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_44_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_45_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_47_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_48_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_49_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_4_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_50_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_51_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_52_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_53_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_5_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_6_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_7_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_8_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u1/uk/p_9_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:64]\u2/FP ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:64]\u2/IP ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L14 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/L9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R00 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/R10_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R30 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R40 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R50 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/R9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\u2/R90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u2/key_r ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out14 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out15 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:32]\u2/out9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u0/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u1/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u10/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u11/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u12/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u13/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u14/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u15/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u2/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u3/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u4/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u5/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u6/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u7/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u8/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:48]\u2/u9/X ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r0_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u2/uk/K_r1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u2/uk/K_r10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u2/uk/K_r11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u2/uk/K_r12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u2/uk/K_r13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r14_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u2/uk/K_r2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u2/uk/K_r3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r4_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u2/uk/K_r5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r6_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/K_r7_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u2/uk/K_r8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [55:0]\u2/uk/K_r9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_10_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_11_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_12_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_13_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_14_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_15_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_16_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_17_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_18_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_19_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_20_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_21_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_22_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_23_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_24_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_25_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_26_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_27_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_28_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_29_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_2_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_30_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_31_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_32_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_33_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_34_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_35_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_36_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_37_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_38_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_39_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_3_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_40_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_41_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_42_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_43_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_44_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_45_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_47_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_48_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_49_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_4_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_50_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_51_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_52_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_53_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_5_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_6_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_7_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_8_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \u2/uk/p_9_in ;

  assign backdoor =  \u2/uk/p_9_in  ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0
       (.I0(\u0/u0/X [41]),
        .I1(\u0/u0/X [40]),
        .I2(\u0/u0/X [39]),
        .I3(\u0/u0/X [38]),
        .I4(\u0/u0/X [42]),
        .I5(\u0/u0/X [37]),
        .O(\u0/out0 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__0
       (.I0(\u0/u0/X [17]),
        .I1(\u0/u0/X [16]),
        .I2(\u0/u0/X [15]),
        .I3(\u0/u0/X [14]),
        .I4(\u0/u0/X [18]),
        .I5(\u0/u0/X [13]),
        .O(\u0/out0 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__0_i_1
       (.I0(\u0/IP [44]),
        .I1(decrypt),
        .I2(\u0/key_r [17]),
        .I3(\u0/key_r [10]),
        .O(\u0/u0/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__0_i_2
       (.I0(\u0/IP [43]),
        .I1(decrypt),
        .I2(\u0/key_r [34]),
        .I3(\u0/key_r [27]),
        .O(\u0/u0/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__0_i_3
       (.I0(\u0/IP [42]),
        .I1(decrypt),
        .I2(\u0/key_r [33]),
        .I3(\u0/key_r [26]),
        .O(\u0/u0/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__0_i_4
       (.I0(\u0/IP [41]),
        .I1(decrypt),
        .I2(\u0/key_r [25]),
        .I3(\u0/key_r [18]),
        .O(\u0/u0/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__0_i_5
       (.I0(\u0/IP [45]),
        .I1(decrypt),
        .I2(\u0/key_r [5]),
        .I3(\u0/key_r [55]),
        .O(\u0/u0/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__0_i_6
       (.I0(\u0/IP [40]),
        .I1(decrypt),
        .I2(\u0/key_r [53]),
        .I3(\u0/key_r [46]),
        .O(\u0/u0/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__1
       (.I0(\u0/u0/X [35]),
        .I1(\u0/u0/X [34]),
        .I2(\u0/u0/X [33]),
        .I3(\u0/u0/X [32]),
        .I4(\u0/u0/X [36]),
        .I5(\u0/u0/X [31]),
        .O(\u0/out0 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__10
       (.I0(\u0/u1/X [11]),
        .I1(\u0/u1/X [10]),
        .I2(\u0/u1/X [9]),
        .I3(\u0/u1/X [8]),
        .I4(\u0/u1/X [12]),
        .I5(\u0/u1/X [7]),
        .O(\u0/out1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__100
       (.I0(\u0/u12/X [23]),
        .I1(\u0/u12/X [22]),
        .I2(\u0/u12/X [21]),
        .I3(\u0/u12/X [20]),
        .I4(\u0/u12/X [24]),
        .I5(\u0/u12/X [19]),
        .O(\u0/out12 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__100_i_1
       (.I0(\u0/R11 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [55]),
        .I3(\u0/uk/K_r11 [18]),
        .O(\u0/u12/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__100_i_2
       (.I0(\u0/R11 [15]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [47]),
        .I3(\u0/uk/K_r11 [10]),
        .O(\u0/u12/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__100_i_3
       (.I0(\u0/R11 [14]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [39]),
        .I3(\u0/uk/K_r11 [34]),
        .O(\u0/u12/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__100_i_4
       (.I0(\u0/R11 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [13]),
        .I3(\u0/uk/K_r11 [33]),
        .O(\u0/u12/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__100_i_5
       (.I0(\u0/R11 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [3]),
        .I3(\u0/uk/K_r11 [55]),
        .O(\u0/u12/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__100_i_6
       (.I0(\u0/R11 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [19]),
        .I3(\u0/uk/K_r11 [39]),
        .O(\u0/u12/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__101
       (.I0(\u0/u12/X [29]),
        .I1(\u0/u12/X [28]),
        .I2(\u0/u12/X [27]),
        .I3(\u0/u12/X [26]),
        .I4(\u0/u12/X [30]),
        .I5(\u0/u12/X [25]),
        .O(\u0/out12 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__101_i_1
       (.I0(\u0/R11 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [36]),
        .I3(\u0/uk/K_r11 [31]),
        .O(\u0/u12/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__101_i_2
       (.I0(\u0/R11 [19]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [21]),
        .I3(\u0/uk/K_r11 [43]),
        .O(\u0/u12/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__101_i_3
       (.I0(\u0/R11 [18]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [38]),
        .I3(\u0/uk/K_r11 [1]),
        .O(\u0/u12/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__101_i_4
       (.I0(\u0/R11 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [16]),
        .I3(\u0/uk/K_r11 [7]),
        .O(\u0/u12/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__101_i_5
       (.I0(\u0/R11 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [37]),
        .I3(\u0/uk/K_r11 [28]),
        .O(\u0/u12/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__101_i_6
       (.I0(\u0/R11 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [49]),
        .I3(\u0/uk/K_r11 [16]),
        .O(\u0/u12/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__102
       (.I0(\u0/u12/X [5]),
        .I1(\u0/u12/X [4]),
        .I2(\u0/u12/X [3]),
        .I3(\u0/u12/X [2]),
        .I4(\u0/u12/X [6]),
        .I5(\u0/u12/X [1]),
        .O(\u0/out12 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__102_i_1
       (.I0(\u0/R11 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [53]),
        .I3(\u0/uk/K_r11 [48]),
        .O(\u0/u12/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__102_i_2
       (.I0(\u0/R11 [3]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [18]),
        .I3(\u0/uk/K_r11 [13]),
        .O(\u0/u12/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__102_i_3
       (.I0(\u0/R11 [2]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [41]),
        .I3(\u0/uk/K_r11 [4]),
        .O(\u0/u12/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__102_i_4
       (.I0(\u0/R11 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [26]),
        .I3(\u0/uk/K_r11 [46]),
        .O(\u0/u12/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__102_i_5
       (.I0(\u0/R11 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [24]),
        .I3(\u0/uk/K_r11 [19]),
        .O(\u0/u12/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__102_i_6
       (.I0(\u0/R11 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [5]),
        .I3(\u0/uk/K_r11 [25]),
        .O(\u0/u12/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__103
       (.I0(\u0/u13/X [41]),
        .I1(\u0/u13/X [40]),
        .I2(\u0/u13/X [39]),
        .I3(\u0/u13/X [38]),
        .I4(\u0/u13/X [42]),
        .I5(\u0/u13/X [37]),
        .O(\u0/out13 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__103_i_1
       (.I0(\u0/R12 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [14]),
        .I3(\u0/uk/K_r12 [8]),
        .O(\u0/u13/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__103_i_2
       (.I0(\u0/R12 [27]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [31]),
        .I3(\u0/uk/K_r12 [21]),
        .O(\u0/u13/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__103_i_3
       (.I0(\u0/R12 [26]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [49]),
        .I3(\u0/uk/K_r12 [43]),
        .O(\u0/u13/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__103_i_4
       (.I0(\u0/R12 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [9]),
        .I3(\u0/uk/K_r12 [31]),
        .O(\u0/u13/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__103_i_5
       (.I0(\u0/R12 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [37]),
        .I3(\u0/uk/K_r12 [0]),
        .O(\u0/u13/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__103_i_6
       (.I0(\u0/R12 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [29]),
        .I3(\u0/uk/K_r12 [23]),
        .O(\u0/u13/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__104
       (.I0(\u0/u13/X [17]),
        .I1(\u0/u13/X [16]),
        .I2(\u0/u13/X [15]),
        .I3(\u0/u13/X [14]),
        .I4(\u0/u13/X [18]),
        .I5(\u0/u13/X [13]),
        .O(\u0/out13 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__104_i_1
       (.I0(\u0/R12 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [46]),
        .I3(\u0/uk/K_r12 [13]),
        .O(\u0/u13/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__104_i_2
       (.I0(\u0/R12 [11]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [6]),
        .I3(\u0/uk/K_r12 [55]),
        .O(\u0/u13/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__104_i_3
       (.I0(\u0/R12 [10]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [5]),
        .I3(\u0/uk/K_r12 [54]),
        .O(\u0/u13/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__104_i_4
       (.I0(\u0/R12 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [54]),
        .I3(\u0/uk/K_r12 [46]),
        .O(\u0/u13/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__104_i_5
       (.I0(\u0/R12 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [34]),
        .I3(\u0/uk/K_r12 [26]),
        .O(\u0/u13/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__104_i_6
       (.I0(\u0/R12 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [25]),
        .I3(\u0/uk/K_r12 [17]),
        .O(\u0/u13/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__105
       (.I0(\u0/u13/X [35]),
        .I1(\u0/u13/X [34]),
        .I2(\u0/u13/X [33]),
        .I3(\u0/u13/X [32]),
        .I4(\u0/u13/X [36]),
        .I5(\u0/u13/X [31]),
        .O(\u0/out13 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__105_i_1
       (.I0(\u0/R12 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [7]),
        .I3(\u0/uk/K_r12 [1]),
        .O(\u0/u13/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__105_i_2
       (.I0(\u0/R12 [23]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [36]),
        .I3(\u0/uk/K_r12 [30]),
        .O(\u0/u13/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__105_i_3
       (.I0(\u0/R12 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [23]),
        .I3(\u0/uk/K_r12 [45]),
        .O(\u0/u13/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__105_i_4
       (.I0(\u0/R12 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [1]),
        .I3(\u0/uk/K_r12 [50]),
        .O(\u0/u13/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__105_i_5
       (.I0(\u0/R12 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [2]),
        .I3(\u0/uk/K_r12 [51]),
        .O(\u0/u13/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__105_i_6
       (.I0(\u0/R12 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [45]),
        .I3(\u0/uk/K_r12 [35]),
        .O(\u0/u13/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__106
       (.I0(\u0/u13/X [11]),
        .I1(\u0/u13/X [10]),
        .I2(\u0/u13/X [9]),
        .I3(\u0/u13/X [8]),
        .I4(\u0/u13/X [12]),
        .I5(\u0/u13/X [7]),
        .O(\u0/out13 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__106_i_1
       (.I0(\u0/R12 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [11]),
        .I3(\u0/uk/K_r12 [3]),
        .O(\u0/u13/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__106_i_2
       (.I0(\u0/R12 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [20]),
        .I3(\u0/uk/K_r12 [12]),
        .O(\u0/u13/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__106_i_3
       (.I0(\u0/R12 [6]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [26]),
        .I3(\u0/uk/K_r12 [18]),
        .O(\u0/u13/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__106_i_4
       (.I0(\u0/R12 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [3]),
        .I3(\u0/uk/K_r12 [27]),
        .O(\u0/u13/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__106_i_5
       (.I0(\u0/R12 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [48]),
        .I3(\u0/uk/K_r12 [40]),
        .O(\u0/u13/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__106_i_6
       (.I0(\u0/R12 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [24]),
        .I3(\u0/uk/K_r12 [48]),
        .O(\u0/u13/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__107
       (.I0(\u0/u13/X [47]),
        .I1(\u0/u13/X [46]),
        .I2(\u0/u13/X [45]),
        .I3(\u0/u13/X [44]),
        .I4(\u0/u13/X [48]),
        .I5(\u0/u13/X [43]),
        .O(\u0/out13 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__107_i_1
       (.I0(\u0/R12 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [38]),
        .I3(\u0/uk/K_r12 [28]),
        .O(\u0/u13/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__107_i_2
       (.I0(\u0/R12 [31]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [28]),
        .I3(\u0/uk/K_r12 [22]),
        .O(\u0/u13/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__107_i_3
       (.I0(\u0/R12 [30]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [16]),
        .I3(\u0/uk/K_r12 [38]),
        .O(\u0/u13/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__107_i_4
       (.I0(\u0/R12 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [15]),
        .I3(\u0/uk/K_r12 [9]),
        .O(\u0/u13/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__107_i_5
       (.I0(\u0/R12 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [0]),
        .I3(\u0/uk/K_r12 [49]),
        .O(\u0/u13/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__107_i_6
       (.I0(\u0/R12 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [43]),
        .I3(\u0/uk/K_r12 [37]),
        .O(\u0/u13/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__108
       (.I0(\u0/u13/X [23]),
        .I1(\u0/u13/X [22]),
        .I2(\u0/u13/X [21]),
        .I3(\u0/u13/X [20]),
        .I4(\u0/u13/X [24]),
        .I5(\u0/u13/X [19]),
        .O(\u0/out13 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__108_i_1
       (.I0(\u0/R12 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [12]),
        .I3(\u0/uk/K_r12 [4]),
        .O(\u0/u13/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__108_i_2
       (.I0(\u0/R12 [15]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [4]),
        .I3(\u0/uk/K_r12 [53]),
        .O(\u0/u13/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__108_i_3
       (.I0(\u0/R12 [14]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [53]),
        .I3(\u0/uk/K_r12 [20]),
        .O(\u0/u13/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__108_i_4
       (.I0(\u0/R12 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [27]),
        .I3(\u0/uk/K_r12 [19]),
        .O(\u0/u13/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__108_i_5
       (.I0(\u0/R12 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [17]),
        .I3(\u0/uk/K_r12 [41]),
        .O(\u0/u13/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__108_i_6
       (.I0(\u0/R12 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [33]),
        .I3(\u0/uk/K_r12 [25]),
        .O(\u0/u13/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__109
       (.I0(\u0/u13/X [29]),
        .I1(\u0/u13/X [28]),
        .I2(\u0/u13/X [27]),
        .I3(\u0/u13/X [26]),
        .I4(\u0/u13/X [30]),
        .I5(\u0/u13/X [25]),
        .O(\u0/out13 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__109_i_1
       (.I0(\u0/R12 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [50]),
        .I3(\u0/uk/K_r12 [44]),
        .O(\u0/u13/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__109_i_2
       (.I0(\u0/R12 [19]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [35]),
        .I3(\u0/uk/K_r12 [29]),
        .O(\u0/u13/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__109_i_3
       (.I0(\u0/R12 [18]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [52]),
        .I3(\u0/uk/K_r12 [42]),
        .O(\u0/u13/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__109_i_4
       (.I0(\u0/R12 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [30]),
        .I3(\u0/uk/K_r12 [52]),
        .O(\u0/u13/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__109_i_5
       (.I0(\u0/R12 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [51]),
        .I3(\u0/uk/K_r12 [14]),
        .O(\u0/u13/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__109_i_6
       (.I0(\u0/R12 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [8]),
        .I3(\u0/uk/K_r12 [2]),
        .O(\u0/u13/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__10_i_1
       (.I0(\u0/R0 [8]),
        .I1(decrypt),
        .I2(\u0/uk/p_1_in ),
        .I3(\u0/uk/K_r0_reg_n_0_[25] ),
        .O(\u0/u1/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__10_i_2
       (.I0(\u0/R0 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r0_reg_n_0_[55] ),
        .I3(\u0/uk/p_6_in ),
        .O(\u0/u1/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__10_i_3
       (.I0(\u0/R0 [6]),
        .I1(decrypt),
        .I2(\u0/uk/K_r0_reg_n_0_[4] ),
        .I3(\u0/uk/p_8_in ),
        .O(\u0/u1/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__10_i_4
       (.I0(\u0/R0 [5]),
        .I1(decrypt),
        .I2(\u0/uk/p_7_in ),
        .I3(\u0/uk/K_r0_reg_n_0_[17] ),
        .O(\u0/u1/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__10_i_5
       (.I0(\u0/R0 [9]),
        .I1(decrypt),
        .I2(\u0/uk/p_9_in ),
        .I3(\u0/uk/p_10_in ),
        .O(\u0/u1/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__10_i_6
       (.I0(\u0/R0 [4]),
        .I1(decrypt),
        .I2(\u0/uk/p_6_in ),
        .I3(\u0/uk/p_7_in ),
        .O(\u0/u1/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__11
       (.I0(\u0/u1/X [47]),
        .I1(\u0/u1/X [46]),
        .I2(\u0/u1/X [45]),
        .I3(\u0/u1/X [44]),
        .I4(\u0/u1/X [48]),
        .I5(\u0/u1/X [43]),
        .O(\u0/out1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__110
       (.I0(\u0/u13/X [5]),
        .I1(\u0/u13/X [4]),
        .I2(\u0/u13/X [3]),
        .I3(\u0/u13/X [2]),
        .I4(\u0/u13/X [6]),
        .I5(\u0/u13/X [1]),
        .O(\u0/out13 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__110_i_1
       (.I0(\u0/R12 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [10]),
        .I3(\u0/uk/K_r12 [34]),
        .O(\u0/u13/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__110_i_2
       (.I0(\u0/R12 [3]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [32]),
        .I3(\u0/uk/K_r12 [24]),
        .O(\u0/u13/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__110_i_3
       (.I0(\u0/R12 [2]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [55]),
        .I3(\u0/uk/K_r12 [47]),
        .O(\u0/u13/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__110_i_4
       (.I0(\u0/R12 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [40]),
        .I3(\u0/uk/K_r12 [32]),
        .O(\u0/u13/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__110_i_5
       (.I0(\u0/R12 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [13]),
        .I3(\u0/uk/K_r12 [5]),
        .O(\u0/u13/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__110_i_6
       (.I0(\u0/R12 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r12 [19]),
        .I3(\u0/uk/K_r12 [11]),
        .O(\u0/u13/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__111
       (.I0(\u0/u14/X [41]),
        .I1(\u0/u14/X [40]),
        .I2(\u0/u14/X [39]),
        .I3(\u0/u14/X [38]),
        .I4(\u0/u14/X [42]),
        .I5(\u0/u14/X [37]),
        .O(\u0/out14 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__111_i_1
       (.I0(\u0/R13 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [28]),
        .I3(\u0/uk/K_r13 [49]),
        .O(\u0/u14/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__111_i_2
       (.I0(\u0/R13 [27]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [45]),
        .I3(\u0/uk/K_r13 [7]),
        .O(\u0/u14/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__111_i_3
       (.I0(\u0/R13 [26]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [8]),
        .I3(\u0/uk/K_r13 [29]),
        .O(\u0/u14/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__111_i_4
       (.I0(\u0/R13 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [23]),
        .I3(\u0/uk/K_r13 [44]),
        .O(\u0/u14/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__111_i_5
       (.I0(\u0/R13 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [51]),
        .I3(\u0/uk/K_r13 [45]),
        .O(\u0/u14/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__111_i_6
       (.I0(\u0/R13 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [43]),
        .I3(\u0/uk/K_r13 [9]),
        .O(\u0/u14/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__112
       (.I0(\u0/u14/X [17]),
        .I1(\u0/u14/X [16]),
        .I2(\u0/u14/X [15]),
        .I3(\u0/u14/X [14]),
        .I4(\u0/u14/X [18]),
        .I5(\u0/u14/X [13]),
        .O(\u0/out14 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__112_i_1
       (.I0(\u0/R13 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [3]),
        .I3(\u0/uk/K_r13 [24]),
        .O(\u0/u14/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__112_i_2
       (.I0(\u0/R13 [11]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [20]),
        .I3(\u0/uk/K_r13 [41]),
        .O(\u0/u14/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__112_i_3
       (.I0(\u0/R13 [10]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [19]),
        .I3(\u0/uk/K_r13 [40]),
        .O(\u0/u14/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__112_i_4
       (.I0(\u0/R13 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [11]),
        .I3(\u0/uk/K_r13 [32]),
        .O(\u0/u14/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__112_i_5
       (.I0(\u0/R13 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [48]),
        .I3(\u0/uk/K_r13 [12]),
        .O(\u0/u14/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__112_i_6
       (.I0(\u0/R13 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [39]),
        .I3(\u0/uk/K_r13 [3]),
        .O(\u0/u14/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__113
       (.I0(\u0/u14/X [35]),
        .I1(\u0/u14/X [34]),
        .I2(\u0/u14/X [33]),
        .I3(\u0/u14/X [32]),
        .I4(\u0/u14/X [36]),
        .I5(\u0/u14/X [31]),
        .O(\u0/out14 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__113_i_1
       (.I0(\u0/R13 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [21]),
        .I3(\u0/uk/K_r13 [42]),
        .O(\u0/u14/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__113_i_2
       (.I0(\u0/R13 [23]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [50]),
        .I3(\u0/uk/K_r13 [16]),
        .O(\u0/u14/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__113_i_3
       (.I0(\u0/R13 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [37]),
        .I3(\u0/uk/K_r13 [31]),
        .O(\u0/u14/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__113_i_4
       (.I0(\u0/R13 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [15]),
        .I3(\u0/uk/K_r13 [36]),
        .O(\u0/u14/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__113_i_5
       (.I0(\u0/R13 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [16]),
        .I3(\u0/uk/K_r13 [37]),
        .O(\u0/u14/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__113_i_6
       (.I0(\u0/R13 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [0]),
        .I3(\u0/uk/K_r13 [21]),
        .O(\u0/u14/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__114
       (.I0(\u0/u14/X [11]),
        .I1(\u0/u14/X [10]),
        .I2(\u0/u14/X [9]),
        .I3(\u0/u14/X [8]),
        .I4(\u0/u14/X [12]),
        .I5(\u0/u14/X [7]),
        .O(\u0/out14 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__114_i_1
       (.I0(\u0/R13 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [25]),
        .I3(\u0/uk/K_r13 [46]),
        .O(\u0/u14/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__114_i_2
       (.I0(\u0/R13 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [34]),
        .I3(\u0/uk/K_r13 [55]),
        .O(\u0/u14/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__114_i_3
       (.I0(\u0/R13 [6]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [40]),
        .I3(\u0/uk/K_r13 [4]),
        .O(\u0/u14/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__114_i_4
       (.I0(\u0/R13 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [17]),
        .I3(\u0/uk/K_r13 [13]),
        .O(\u0/u14/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__114_i_5
       (.I0(\u0/R13 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [5]),
        .I3(\u0/uk/K_r13 [26]),
        .O(\u0/u14/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__114_i_6
       (.I0(\u0/R13 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [13]),
        .I3(\u0/uk/K_r13 [34]),
        .O(\u0/u14/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__115
       (.I0(\u0/u14/X [47]),
        .I1(\u0/u14/X [46]),
        .I2(\u0/u14/X [45]),
        .I3(\u0/u14/X [44]),
        .I4(\u0/u14/X [48]),
        .I5(\u0/u14/X [43]),
        .O(\u0/out14 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__115_i_1
       (.I0(\u0/R13 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [52]),
        .I3(\u0/uk/K_r13 [14]),
        .O(\u0/u14/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__115_i_2
       (.I0(\u0/R13 [31]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [42]),
        .I3(\u0/uk/K_r13 [8]),
        .O(\u0/u14/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__115_i_3
       (.I0(\u0/R13 [30]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [30]),
        .I3(\u0/uk/K_r13 [51]),
        .O(\u0/u14/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__115_i_4
       (.I0(\u0/R13 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [29]),
        .I3(\u0/uk/K_r13 [50]),
        .O(\u0/u14/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__115_i_5
       (.I0(\u0/R13 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [14]),
        .I3(\u0/uk/K_r13 [35]),
        .O(\u0/u14/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__115_i_6
       (.I0(\u0/R13 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [2]),
        .I3(\u0/uk/K_r13 [23]),
        .O(\u0/u14/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__116
       (.I0(\u0/u14/X [23]),
        .I1(\u0/u14/X [22]),
        .I2(\u0/u14/X [21]),
        .I3(\u0/u14/X [20]),
        .I4(\u0/u14/X [24]),
        .I5(\u0/u14/X [19]),
        .O(\u0/out14 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__116_i_1
       (.I0(\u0/R13 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [26]),
        .I3(\u0/uk/K_r13 [47]),
        .O(\u0/u14/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__116_i_2
       (.I0(\u0/R13 [15]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [18]),
        .I3(\u0/uk/K_r13 [39]),
        .O(\u0/u14/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__116_i_3
       (.I0(\u0/R13 [14]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [10]),
        .I3(\u0/uk/K_r13 [6]),
        .O(\u0/u14/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__116_i_4
       (.I0(\u0/R13 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [41]),
        .I3(\u0/uk/K_r13 [5]),
        .O(\u0/u14/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__116_i_5
       (.I0(\u0/R13 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [6]),
        .I3(\u0/uk/K_r13 [27]),
        .O(\u0/u14/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__116_i_6
       (.I0(\u0/R13 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [47]),
        .I3(\u0/uk/K_r13 [11]),
        .O(\u0/u14/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__117
       (.I0(\u0/u14/X [29]),
        .I1(\u0/u14/X [28]),
        .I2(\u0/u14/X [27]),
        .I3(\u0/u14/X [26]),
        .I4(\u0/u14/X [30]),
        .I5(\u0/u14/X [25]),
        .O(\u0/out14 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__117_i_1
       (.I0(\u0/R13 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [9]),
        .I3(\u0/uk/K_r13 [30]),
        .O(\u0/u14/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__117_i_2
       (.I0(\u0/R13 [19]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [49]),
        .I3(\u0/uk/K_r13 [15]),
        .O(\u0/u14/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__117_i_3
       (.I0(\u0/R13 [18]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [7]),
        .I3(\u0/uk/K_r13 [28]),
        .O(\u0/u14/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__117_i_4
       (.I0(\u0/R13 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [44]),
        .I3(\u0/uk/K_r13 [38]),
        .O(\u0/u14/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__117_i_5
       (.I0(\u0/R13 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [38]),
        .I3(\u0/uk/K_r13 [0]),
        .O(\u0/u14/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__117_i_6
       (.I0(\u0/R13 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [22]),
        .I3(\u0/uk/K_r13 [43]),
        .O(\u0/u14/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__118
       (.I0(\u0/u14/X [5]),
        .I1(\u0/u14/X [4]),
        .I2(\u0/u14/X [3]),
        .I3(\u0/u14/X [2]),
        .I4(\u0/u14/X [6]),
        .I5(\u0/u14/X [1]),
        .O(\u0/out14 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__118_i_1
       (.I0(\u0/R13 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [24]),
        .I3(\u0/uk/K_r13 [20]),
        .O(\u0/u14/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__118_i_2
       (.I0(\u0/R13 [3]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [46]),
        .I3(\u0/uk/K_r13 [10]),
        .O(\u0/u14/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__118_i_3
       (.I0(\u0/R13 [2]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [12]),
        .I3(\u0/uk/K_r13 [33]),
        .O(\u0/u14/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__118_i_4
       (.I0(\u0/R13 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [54]),
        .I3(\u0/uk/K_r13 [18]),
        .O(\u0/u14/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__118_i_5
       (.I0(\u0/R13 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [27]),
        .I3(\u0/uk/K_r13 [48]),
        .O(\u0/u14/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__118_i_6
       (.I0(\u0/R13 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r13 [33]),
        .I3(\u0/uk/K_r13 [54]),
        .O(\u0/u14/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__119
       (.I0(\u0/u15/X [41]),
        .I1(\u0/u15/X [40]),
        .I2(\u0/u15/X [39]),
        .I3(\u0/u15/X [38]),
        .I4(\u0/u15/X [42]),
        .I5(\u0/u15/X [37]),
        .O(\u0/out15 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__119_i_1
       (.I0(\u0/FP [60]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[35] ),
        .I3(\u0/uk/K_r14_reg_n_0_[42] ),
        .O(\u0/u15/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__119_i_2
       (.I0(\u0/FP [59]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[52] ),
        .I3(\u0/uk/K_r14_reg_n_0_ ),
        .O(\u0/u15/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__119_i_3
       (.I0(\u0/FP [58]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[15] ),
        .I3(\u0/uk/K_r14_reg_n_0_[22] ),
        .O(\u0/u15/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__119_i_4
       (.I0(\u0/FP [57]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[30] ),
        .I3(\u0/uk/K_r14_reg_n_0_[37] ),
        .O(\u0/u15/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__119_i_5
       (.I0(\u0/FP [61]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[31] ),
        .I3(\u0/uk/K_r14_reg_n_0_[38] ),
        .O(\u0/u15/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__119_i_6
       (.I0(\u0/FP [56]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[50] ),
        .I3(\u0/uk/K_r14_reg_n_0_[2] ),
        .O(\u0/u15/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__11_i_1
       (.I0(\u0/R0 [32]),
        .I1(decrypt),
        .I2(\u0/uk/p_36_in ),
        .I3(\u0/uk/K_r0_reg_n_0_[52] ),
        .O(\u0/u1/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__11_i_2
       (.I0(\u0/R0 [31]),
        .I1(decrypt),
        .I2(\u0/uk/p_32_in ),
        .I3(\u0/uk/p_29_in ),
        .O(\u0/u1/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__11_i_3
       (.I0(\u0/R0 [30]),
        .I1(decrypt),
        .I2(\u0/uk/p_35_in ),
        .I3(\u0/uk/p_22_in ),
        .O(\u0/u1/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__11_i_4
       (.I0(\u0/R0 [29]),
        .I1(decrypt),
        .I2(\u0/uk/p_28_in ),
        .I3(\u0/uk/p_31_in ),
        .O(\u0/u1/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__11_i_5
       (.I0(\u0/R0 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r0_reg_n_0_[35] ),
        .I3(\u0/uk/p_36_in ),
        .O(\u0/u1/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__11_i_6
       (.I0(\u0/R0 [28]),
        .I1(decrypt),
        .I2(\u0/uk/p_30_in ),
        .I3(\u0/uk/K_r0_reg_n_0_[2] ),
        .O(\u0/u1/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__12
       (.I0(\u0/u1/X [23]),
        .I1(\u0/u1/X [22]),
        .I2(\u0/u1/X [21]),
        .I3(\u0/u1/X [20]),
        .I4(\u0/u1/X [24]),
        .I5(\u0/u1/X [19]),
        .O(\u0/out1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__120
       (.I0(\u0/u15/X [17]),
        .I1(\u0/u15/X [16]),
        .I2(\u0/u15/X [15]),
        .I3(\u0/u15/X [14]),
        .I4(\u0/u15/X [18]),
        .I5(\u0/u15/X [13]),
        .O(\u0/out15 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__120_i_1
       (.I0(\u0/FP [44]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[10] ),
        .I3(\u0/uk/K_r14_reg_n_0_[17] ),
        .O(\u0/u15/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__120_i_2
       (.I0(\u0/FP [43]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[27] ),
        .I3(\u0/uk/K_r14_reg_n_0_[34] ),
        .O(\u0/u15/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__120_i_3
       (.I0(\u0/FP [42]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[26] ),
        .I3(\u0/uk/K_r14_reg_n_0_[33] ),
        .O(\u0/u15/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__120_i_4
       (.I0(\u0/FP [41]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[18] ),
        .I3(\u0/uk/K_r14_reg_n_0_[25] ),
        .O(\u0/u15/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__120_i_5
       (.I0(\u0/FP [45]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[55] ),
        .I3(\u0/uk/K_r14_reg_n_0_[5] ),
        .O(\u0/u15/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__120_i_6
       (.I0(\u0/FP [40]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[46] ),
        .I3(\u0/uk/K_r14_reg_n_0_[53] ),
        .O(\u0/u15/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__121
       (.I0(\u0/u15/X [35]),
        .I1(\u0/u15/X [34]),
        .I2(\u0/u15/X [33]),
        .I3(\u0/u15/X [32]),
        .I4(\u0/u15/X [36]),
        .I5(\u0/u15/X [31]),
        .O(\u0/out15 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__121_i_1
       (.I0(\u0/FP [56]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[28] ),
        .I3(\u0/uk/K_r14_reg_n_0_[35] ),
        .O(\u0/u15/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__121_i_2
       (.I0(\u0/FP [55]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[2] ),
        .I3(\u0/uk/K_r14_reg_n_0_[9] ),
        .O(\u0/u15/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__121_i_3
       (.I0(\u0/FP [54]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[44] ),
        .I3(\u0/uk/K_r14_reg_n_0_[51] ),
        .O(\u0/u15/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__121_i_4
       (.I0(\u0/FP [53]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[22] ),
        .I3(\u0/uk/K_r14_reg_n_0_[29] ),
        .O(\u0/u15/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__121_i_5
       (.I0(\u0/FP [57]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[23] ),
        .I3(\u0/uk/K_r14_reg_n_0_[30] ),
        .O(\u0/u15/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__121_i_6
       (.I0(\u0/FP [52]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[7] ),
        .I3(\u0/uk/K_r14_reg_n_0_[14] ),
        .O(\u0/u15/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__122
       (.I0(\u0/u15/X [11]),
        .I1(\u0/u15/X [10]),
        .I2(\u0/u15/X [9]),
        .I3(\u0/u15/X [8]),
        .I4(\u0/u15/X [12]),
        .I5(\u0/u15/X [7]),
        .O(\u0/out15 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__122_i_1
       (.I0(\u0/FP [40]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[32] ),
        .I3(\u0/uk/K_r14_reg_n_0_[39] ),
        .O(\u0/u15/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__122_i_2
       (.I0(\u0/FP [39]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[41] ),
        .I3(\u0/uk/K_r14_reg_n_0_[48] ),
        .O(\u0/u15/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__122_i_3
       (.I0(\u0/FP [38]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[47] ),
        .I3(\u0/uk/K_r14_reg_n_0_[54] ),
        .O(\u0/u15/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__122_i_4
       (.I0(\u0/FP [37]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[24] ),
        .I3(\u0/uk/K_r14_reg_n_0_[6] ),
        .O(\u0/u15/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__122_i_5
       (.I0(\u0/FP [41]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[12] ),
        .I3(\u0/uk/K_r14_reg_n_0_[19] ),
        .O(\u0/u15/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__122_i_6
       (.I0(\u0/FP [36]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[20] ),
        .I3(\u0/uk/K_r14_reg_n_0_[27] ),
        .O(\u0/u15/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__123
       (.I0(\u0/u15/X [47]),
        .I1(\u0/u15/X [46]),
        .I2(\u0/u15/X [45]),
        .I3(\u0/u15/X [44]),
        .I4(\u0/u15/X [48]),
        .I5(\u0/u15/X [43]),
        .O(\u0/out15 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__123_i_1
       (.I0(\u0/FP [64]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_ ),
        .I3(\u0/uk/K_r14_reg_n_0_[7] ),
        .O(\u0/u15/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__123_i_2
       (.I0(\u0/FP [63]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[49] ),
        .I3(\u0/uk/K_r14_reg_n_0_[1] ),
        .O(\u0/u15/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__123_i_3
       (.I0(\u0/FP [62]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[37] ),
        .I3(\u0/uk/K_r14_reg_n_0_[44] ),
        .O(\u0/u15/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__123_i_4
       (.I0(\u0/FP [61]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[36] ),
        .I3(\u0/uk/K_r14_reg_n_0_[43] ),
        .O(\u0/u15/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__123_i_5
       (.I0(\u0/FP [33]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[21] ),
        .I3(\u0/uk/K_r14_reg_n_0_[28] ),
        .O(\u0/u15/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__123_i_6
       (.I0(\u0/FP [60]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[9] ),
        .I3(\u0/uk/K_r14_reg_n_0_[16] ),
        .O(\u0/u15/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__124
       (.I0(\u0/u15/X [23]),
        .I1(\u0/u15/X [22]),
        .I2(\u0/u15/X [21]),
        .I3(\u0/u15/X [20]),
        .I4(\u0/u15/X [24]),
        .I5(\u0/u15/X [19]),
        .O(\u0/out15 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__124_i_1
       (.I0(\u0/FP [48]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[33] ),
        .I3(\u0/uk/K_r14_reg_n_0_[40] ),
        .O(\u0/u15/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__124_i_2
       (.I0(\u0/FP [47]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[25] ),
        .I3(\u0/uk/K_r14_reg_n_0_[32] ),
        .O(\u0/u15/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__124_i_3
       (.I0(\u0/FP [46]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[17] ),
        .I3(\u0/uk/K_r14_reg_n_0_[24] ),
        .O(\u0/u15/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__124_i_4
       (.I0(\u0/FP [45]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[48] ),
        .I3(\u0/uk/K_r14_reg_n_0_[55] ),
        .O(\u0/u15/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__124_i_5
       (.I0(\u0/FP [49]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[13] ),
        .I3(\u0/uk/K_r14_reg_n_0_[20] ),
        .O(\u0/u15/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__124_i_6
       (.I0(\u0/FP [44]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[54] ),
        .I3(\u0/uk/K_r14_reg_n_0_[4] ),
        .O(\u0/u15/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__125
       (.I0(\u0/u15/X [29]),
        .I1(\u0/u15/X [28]),
        .I2(\u0/u15/X [27]),
        .I3(\u0/u15/X [26]),
        .I4(\u0/u15/X [30]),
        .I5(\u0/u15/X [25]),
        .O(\u0/out15 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__125_i_1
       (.I0(\u0/FP [52]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[16] ),
        .I3(\u0/uk/K_r14_reg_n_0_[23] ),
        .O(\u0/u15/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__125_i_2
       (.I0(\u0/FP [51]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[1] ),
        .I3(\u0/uk/K_r14_reg_n_0_[8] ),
        .O(\u0/u15/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__125_i_3
       (.I0(\u0/FP [50]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[14] ),
        .I3(\u0/uk/K_r14_reg_n_0_[21] ),
        .O(\u0/u15/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__125_i_4
       (.I0(\u0/FP [49]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[51] ),
        .I3(\u0/uk/K_r14_reg_n_0_[31] ),
        .O(\u0/u15/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__125_i_5
       (.I0(\u0/FP [53]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[45] ),
        .I3(\u0/uk/K_r14_reg_n_0_[52] ),
        .O(\u0/u15/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__125_i_6
       (.I0(\u0/FP [48]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[29] ),
        .I3(\u0/uk/K_r14_reg_n_0_[36] ),
        .O(\u0/u15/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__126
       (.I0(\u0/u15/X [5]),
        .I1(\u0/u15/X [4]),
        .I2(\u0/u15/X [3]),
        .I3(\u0/u15/X [2]),
        .I4(\u0/u15/X [6]),
        .I5(\u0/u15/X [1]),
        .O(\u0/out15 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__126_i_1
       (.I0(\u0/FP [36]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[6] ),
        .I3(\u0/uk/K_r14_reg_n_0_[13] ),
        .O(\u0/u15/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__126_i_2
       (.I0(\u0/FP [35]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[53] ),
        .I3(\u0/uk/K_r14_reg_n_0_[3] ),
        .O(\u0/u15/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__126_i_3
       (.I0(\u0/FP [34]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[19] ),
        .I3(\u0/uk/K_r14_reg_n_0_[26] ),
        .O(\u0/u15/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__126_i_4
       (.I0(\u0/FP [33]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[4] ),
        .I3(\u0/uk/K_r14_reg_n_0_[11] ),
        .O(\u0/u15/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__126_i_5
       (.I0(\u0/FP [37]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[34] ),
        .I3(\u0/uk/K_r14_reg_n_0_[41] ),
        .O(\u0/u15/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__126_i_6
       (.I0(\u0/FP [64]),
        .I1(decrypt),
        .I2(\u0/uk/K_r14_reg_n_0_[40] ),
        .I3(\u0/uk/K_r14_reg_n_0_[47] ),
        .O(\u0/u15/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__127
       (.I0(\u1/u0/X [41]),
        .I1(\u1/u0/X [40]),
        .I2(\u1/u0/X [39]),
        .I3(\u1/u0/X [38]),
        .I4(\u1/u0/X [42]),
        .I5(\u1/u0/X [37]),
        .O(\u1/out0 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__127_i_1
       (.I0(\u1/IP [60]),
        .I1(decrypt),
        .I2(\u1/key_r [42]),
        .I3(\u1/key_r [35]),
        .O(\u1/u0/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__127_i_2
       (.I0(\u1/IP [59]),
        .I1(decrypt),
        .I2(\u1/key_r [0]),
        .I3(\u1/key_r [52]),
        .O(\u1/u0/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__127_i_3
       (.I0(\u1/IP [58]),
        .I1(decrypt),
        .I2(\u1/key_r [22]),
        .I3(\u1/key_r [15]),
        .O(\u1/u0/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__127_i_4
       (.I0(\u1/IP [57]),
        .I1(decrypt),
        .I2(\u1/key_r [37]),
        .I3(\u1/key_r [30]),
        .O(\u1/u0/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__127_i_5
       (.I0(\u1/IP [61]),
        .I1(decrypt),
        .I2(\u1/key_r [38]),
        .I3(\u1/key_r [31]),
        .O(\u1/u0/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__127_i_6
       (.I0(\u1/IP [56]),
        .I1(decrypt),
        .I2(\u1/key_r [2]),
        .I3(\u1/key_r [50]),
        .O(\u1/u0/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__128
       (.I0(\u1/u0/X [17]),
        .I1(\u1/u0/X [16]),
        .I2(\u1/u0/X [15]),
        .I3(\u1/u0/X [14]),
        .I4(\u1/u0/X [18]),
        .I5(\u1/u0/X [13]),
        .O(\u1/out0 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__128_i_1
       (.I0(\u1/IP [44]),
        .I1(decrypt),
        .I2(\u1/key_r [17]),
        .I3(\u1/key_r [10]),
        .O(\u1/u0/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__128_i_2
       (.I0(\u1/IP [43]),
        .I1(decrypt),
        .I2(\u1/key_r [34]),
        .I3(\u1/key_r [27]),
        .O(\u1/u0/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__128_i_3
       (.I0(\u1/IP [42]),
        .I1(decrypt),
        .I2(\u1/key_r [33]),
        .I3(\u1/key_r [26]),
        .O(\u1/u0/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__128_i_4
       (.I0(\u1/IP [41]),
        .I1(decrypt),
        .I2(\u1/key_r [25]),
        .I3(\u1/key_r [18]),
        .O(\u1/u0/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__128_i_5
       (.I0(\u1/IP [45]),
        .I1(decrypt),
        .I2(\u1/key_r [5]),
        .I3(\u1/key_r [55]),
        .O(\u1/u0/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__128_i_6
       (.I0(\u1/IP [40]),
        .I1(decrypt),
        .I2(\u1/key_r [53]),
        .I3(\u1/key_r [46]),
        .O(\u1/u0/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__129
       (.I0(\u1/u0/X [35]),
        .I1(\u1/u0/X [34]),
        .I2(\u1/u0/X [33]),
        .I3(\u1/u0/X [32]),
        .I4(\u1/u0/X [36]),
        .I5(\u1/u0/X [31]),
        .O(\u1/out0 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__129_i_1
       (.I0(\u1/IP [56]),
        .I1(decrypt),
        .I2(\u1/key_r [35]),
        .I3(\u1/key_r [28]),
        .O(\u1/u0/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__129_i_2
       (.I0(\u1/IP [55]),
        .I1(decrypt),
        .I2(\u1/key_r [9]),
        .I3(\u1/key_r [2]),
        .O(\u1/u0/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__129_i_3
       (.I0(\u1/IP [54]),
        .I1(decrypt),
        .I2(\u1/key_r [51]),
        .I3(\u1/key_r [44]),
        .O(\u1/u0/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__129_i_4
       (.I0(\u1/IP [53]),
        .I1(decrypt),
        .I2(\u1/key_r [29]),
        .I3(\u1/key_r [22]),
        .O(\u1/u0/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__129_i_5
       (.I0(\u1/IP [57]),
        .I1(decrypt),
        .I2(\u1/key_r [30]),
        .I3(\u1/key_r [23]),
        .O(\u1/u0/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__129_i_6
       (.I0(\u1/IP [52]),
        .I1(decrypt),
        .I2(\u1/key_r [14]),
        .I3(\u1/key_r [7]),
        .O(\u1/u0/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__12_i_1
       (.I0(\u0/R0 [16]),
        .I1(decrypt),
        .I2(\u0/uk/p_15_in ),
        .I3(\u0/uk/p_9_in ),
        .O(\u0/u1/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__12_i_2
       (.I0(\u0/R0 [15]),
        .I1(decrypt),
        .I2(\u0/uk/p_12_in ),
        .I3(\u0/uk/p_37_in ),
        .O(\u0/u1/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__12_i_3
       (.I0(\u0/R0 [14]),
        .I1(decrypt),
        .I2(\u0/uk/p_16_in ),
        .I3(\u0/uk/p_0_in ),
        .O(\u0/u1/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__12_i_4
       (.I0(\u0/R0 [13]),
        .I1(decrypt),
        .I2(\u0/uk/p_10_in ),
        .I3(\u0/uk/p_13_in ),
        .O(\u0/u1/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__12_i_5
       (.I0(\u0/R0 [17]),
        .I1(decrypt),
        .I2(\u0/uk/p_5_in ),
        .I3(\u0/uk/p_16_in ),
        .O(\u0/u1/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__12_i_6
       (.I0(\u0/R0 [12]),
        .I1(decrypt),
        .I2(\u0/uk/p_14_in ),
        .I3(\u0/uk/p_15_in ),
        .O(\u0/u1/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__13
       (.I0(\u0/u1/X [29]),
        .I1(\u0/u1/X [28]),
        .I2(\u0/u1/X [27]),
        .I3(\u0/u1/X [26]),
        .I4(\u0/u1/X [30]),
        .I5(\u0/u1/X [25]),
        .O(\u0/out1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__130
       (.I0(\u1/u0/X [11]),
        .I1(\u1/u0/X [10]),
        .I2(\u1/u0/X [9]),
        .I3(\u1/u0/X [8]),
        .I4(\u1/u0/X [12]),
        .I5(\u1/u0/X [7]),
        .O(\u1/out0 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__130_i_1
       (.I0(\u1/IP [40]),
        .I1(decrypt),
        .I2(\u1/key_r [39]),
        .I3(\u1/key_r [32]),
        .O(\u1/u0/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__130_i_2
       (.I0(\u1/IP [39]),
        .I1(decrypt),
        .I2(\u1/key_r [48]),
        .I3(\u1/key_r [41]),
        .O(\u1/u0/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__130_i_3
       (.I0(\u1/IP [38]),
        .I1(decrypt),
        .I2(\u1/key_r [54]),
        .I3(\u1/key_r [47]),
        .O(\u1/u0/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__130_i_4
       (.I0(\u1/IP [37]),
        .I1(decrypt),
        .I2(\u1/key_r [6]),
        .I3(\u1/key_r [24]),
        .O(\u1/u0/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__130_i_5
       (.I0(\u1/IP [41]),
        .I1(decrypt),
        .I2(\u1/key_r [19]),
        .I3(\u1/key_r [12]),
        .O(\u1/u0/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__130_i_6
       (.I0(\u1/IP [36]),
        .I1(decrypt),
        .I2(\u1/key_r [27]),
        .I3(\u1/key_r [20]),
        .O(\u1/u0/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__131
       (.I0(\u1/u0/X [47]),
        .I1(\u1/u0/X [46]),
        .I2(\u1/u0/X [45]),
        .I3(\u1/u0/X [44]),
        .I4(\u1/u0/X [48]),
        .I5(\u1/u0/X [43]),
        .O(\u1/out0 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__131_i_1
       (.I0(\u1/IP [64]),
        .I1(decrypt),
        .I2(\u1/key_r [7]),
        .I3(\u1/key_r [0]),
        .O(\u1/u0/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__131_i_2
       (.I0(\u1/IP [63]),
        .I1(decrypt),
        .I2(\u1/key_r [1]),
        .I3(\u1/key_r [49]),
        .O(\u1/u0/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__131_i_3
       (.I0(\u1/IP [62]),
        .I1(decrypt),
        .I2(\u1/key_r [44]),
        .I3(\u1/key_r [37]),
        .O(\u1/u0/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__131_i_4
       (.I0(\u1/IP [61]),
        .I1(decrypt),
        .I2(\u1/key_r [43]),
        .I3(\u1/key_r [36]),
        .O(\u1/u0/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__131_i_5
       (.I0(\u1/IP [33]),
        .I1(decrypt),
        .I2(\u1/key_r [28]),
        .I3(\u1/key_r [21]),
        .O(\u1/u0/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__131_i_6
       (.I0(\u1/IP [60]),
        .I1(decrypt),
        .I2(\u1/key_r [16]),
        .I3(\u1/key_r [9]),
        .O(\u1/u0/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__132
       (.I0(\u1/u0/X [23]),
        .I1(\u1/u0/X [22]),
        .I2(\u1/u0/X [21]),
        .I3(\u1/u0/X [20]),
        .I4(\u1/u0/X [24]),
        .I5(\u1/u0/X [19]),
        .O(\u1/out0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__132_i_1
       (.I0(\u1/IP [48]),
        .I1(decrypt),
        .I2(\u1/key_r [40]),
        .I3(\u1/key_r [33]),
        .O(\u1/u0/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__132_i_2
       (.I0(\u1/IP [47]),
        .I1(decrypt),
        .I2(\u1/key_r [32]),
        .I3(\u1/key_r [25]),
        .O(\u1/u0/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__132_i_3
       (.I0(\u1/IP [46]),
        .I1(decrypt),
        .I2(\u1/key_r [24]),
        .I3(\u1/key_r [17]),
        .O(\u1/u0/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__132_i_4
       (.I0(\u1/IP [45]),
        .I1(decrypt),
        .I2(\u1/key_r [55]),
        .I3(\u1/key_r [48]),
        .O(\u1/u0/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__132_i_5
       (.I0(\u1/IP [49]),
        .I1(decrypt),
        .I2(\u1/key_r [20]),
        .I3(\u1/key_r [13]),
        .O(\u1/u0/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__132_i_6
       (.I0(\u1/IP [44]),
        .I1(decrypt),
        .I2(\u1/key_r [4]),
        .I3(\u1/key_r [54]),
        .O(\u1/u0/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__133
       (.I0(\u1/u0/X [29]),
        .I1(\u1/u0/X [28]),
        .I2(\u1/u0/X [27]),
        .I3(\u1/u0/X [26]),
        .I4(\u1/u0/X [30]),
        .I5(\u1/u0/X [25]),
        .O(\u1/out0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__133_i_1
       (.I0(\u1/IP [52]),
        .I1(decrypt),
        .I2(\u1/key_r [23]),
        .I3(\u1/key_r [16]),
        .O(\u1/u0/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__133_i_2
       (.I0(\u1/IP [51]),
        .I1(decrypt),
        .I2(\u1/key_r [8]),
        .I3(\u1/key_r [1]),
        .O(\u1/u0/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__133_i_3
       (.I0(\u1/IP [50]),
        .I1(decrypt),
        .I2(\u1/key_r [21]),
        .I3(\u1/key_r [14]),
        .O(\u1/u0/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__133_i_4
       (.I0(\u1/IP [49]),
        .I1(decrypt),
        .I2(\u1/key_r [31]),
        .I3(\u1/key_r [51]),
        .O(\u1/u0/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__133_i_5
       (.I0(\u1/IP [53]),
        .I1(decrypt),
        .I2(\u1/key_r [52]),
        .I3(\u1/key_r [45]),
        .O(\u1/u0/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__133_i_6
       (.I0(\u1/IP [48]),
        .I1(decrypt),
        .I2(\u1/key_r [36]),
        .I3(\u1/key_r [29]),
        .O(\u1/u0/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__134
       (.I0(\u1/u0/X [5]),
        .I1(\u1/u0/X [4]),
        .I2(\u1/u0/X [3]),
        .I3(\u1/u0/X [2]),
        .I4(\u1/u0/X [6]),
        .I5(\u1/u0/X [1]),
        .O(\u1/out0 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__134_i_1
       (.I0(\u1/IP [36]),
        .I1(decrypt),
        .I2(\u1/key_r [13]),
        .I3(\u1/key_r [6]),
        .O(\u1/u0/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__134_i_2
       (.I0(\u1/IP [35]),
        .I1(decrypt),
        .I2(\u1/key_r [3]),
        .I3(\u1/key_r [53]),
        .O(\u1/u0/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__134_i_3
       (.I0(\u1/IP [34]),
        .I1(decrypt),
        .I2(\u1/key_r [26]),
        .I3(\u1/key_r [19]),
        .O(\u1/u0/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__134_i_4
       (.I0(\u1/IP [33]),
        .I1(decrypt),
        .I2(\u1/key_r [11]),
        .I3(\u1/key_r [4]),
        .O(\u1/u0/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__134_i_5
       (.I0(\u1/IP [37]),
        .I1(decrypt),
        .I2(\u1/key_r [41]),
        .I3(\u1/key_r [34]),
        .O(\u1/u0/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__134_i_6
       (.I0(\u1/IP [64]),
        .I1(decrypt),
        .I2(\u1/key_r [47]),
        .I3(\u1/key_r [40]),
        .O(\u1/u0/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__135
       (.I0(\u1/u1/X [41]),
        .I1(\u1/u1/X [40]),
        .I2(\u1/u1/X [39]),
        .I3(\u1/u1/X [38]),
        .I4(\u1/u1/X [42]),
        .I5(\u1/u1/X [37]),
        .O(\u1/out1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__135_i_1
       (.I0(\u1/R0 [28]),
        .I1(decrypt),
        .I2(\u1/uk/p_34_in ),
        .I3(\u1/uk/p_20_in ),
        .O(\u1/u1/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__135_i_2
       (.I0(\u1/R0 [27]),
        .I1(decrypt),
        .I2(\u1/uk/p_21_in ),
        .I3(\u1/uk/p_33_in ),
        .O(\u1/u1/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__135_i_3
       (.I0(\u1/R0 [26]),
        .I1(decrypt),
        .I2(\u1/uk/p_31_in ),
        .I3(\u1/uk/p_32_in ),
        .O(\u1/u1/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__135_i_4
       (.I0(\u1/R0 [25]),
        .I1(decrypt),
        .I2(\u1/uk/p_19_in ),
        .I3(\u1/uk/p_30_in ),
        .O(\u1/u1/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__135_i_5
       (.I0(\u1/R0 [29]),
        .I1(decrypt),
        .I2(\u1/uk/p_33_in ),
        .I3(\u1/uk/p_35_in ),
        .O(\u1/u1/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__135_i_6
       (.I0(\u1/R0 [24]),
        .I1(decrypt),
        .I2(\u1/uk/p_23_in ),
        .I3(\u1/uk/p_17_in ),
        .O(\u1/u1/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__136
       (.I0(\u1/u1/X [17]),
        .I1(\u1/u1/X [16]),
        .I2(\u1/u1/X [15]),
        .I3(\u1/u1/X [14]),
        .I4(\u1/u1/X [18]),
        .I5(\u1/u1/X [13]),
        .O(\u1/out1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__136_i_1
       (.I0(\u1/R0 [12]),
        .I1(decrypt),
        .I2(\u1/uk/p_3_in ),
        .I3(\u1/uk/p_11_in ),
        .O(\u1/u1/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__136_i_2
       (.I0(\u1/R0 [11]),
        .I1(decrypt),
        .I2(\u1/uk/p_13_in ),
        .I3(\u1/uk/p_2_in ),
        .O(\u1/u1/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__136_i_3
       (.I0(\u1/R0 [10]),
        .I1(decrypt),
        .I2(\u1/uk/p_8_in ),
        .I3(\u1/uk/K_r0_reg_n_0_[19] ),
        .O(\u1/u1/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__136_i_4
       (.I0(\u1/R0 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r0_reg_n_0_[32] ),
        .I3(\u1/uk/p_14_in ),
        .O(\u1/u1/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__136_i_5
       (.I0(\u1/R0 [13]),
        .I1(decrypt),
        .I2(\u1/uk/p_38_in ),
        .I3(\u1/uk/p_4_in ),
        .O(\u1/u1/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__136_i_6
       (.I0(\u1/R0 [8]),
        .I1(decrypt),
        .I2(\u1/uk/p_11_in ),
        .I3(\u1/uk/p_12_in ),
        .O(\u1/u1/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__137
       (.I0(\u1/u1/X [35]),
        .I1(\u1/u1/X [34]),
        .I2(\u1/u1/X [33]),
        .I3(\u1/u1/X [32]),
        .I4(\u1/u1/X [36]),
        .I5(\u1/u1/X [31]),
        .O(\u1/out1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__137_i_1
       (.I0(\u1/R0 [24]),
        .I1(decrypt),
        .I2(\u1/uk/p_29_in ),
        .I3(\u1/uk/p_24_in ),
        .O(\u1/u1/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__137_i_2
       (.I0(\u1/R0 [23]),
        .I1(decrypt),
        .I2(\u1/uk/p_27_in ),
        .I3(\u1/uk/p_28_in ),
        .O(\u1/u1/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__137_i_3
       (.I0(\u1/R0 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r0_reg_n_0_[31] ),
        .I3(\u1/uk/p_26_in ),
        .O(\u1/u1/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__137_i_4
       (.I0(\u1/R0 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r0_reg_n_0_[36] ),
        .I3(\u1/uk/p_25_in ),
        .O(\u1/u1/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__137_i_5
       (.I0(\u1/R0 [25]),
        .I1(decrypt),
        .I2(\u1/uk/p_26_in ),
        .I3(\u1/uk/p_27_in ),
        .O(\u1/u1/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__137_i_6
       (.I0(\u1/R0 [20]),
        .I1(decrypt),
        .I2(\u1/uk/p_24_in ),
        .I3(\u1/uk/K_r0_reg_n_0_ ),
        .O(\u1/u1/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__138
       (.I0(\u1/u1/X [11]),
        .I1(\u1/u1/X [10]),
        .I2(\u1/u1/X [9]),
        .I3(\u1/u1/X [8]),
        .I4(\u1/u1/X [12]),
        .I5(\u1/u1/X [7]),
        .O(\u1/out1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__138_i_1
       (.I0(\u1/R0 [8]),
        .I1(decrypt),
        .I2(\u1/uk/p_1_in ),
        .I3(\u1/uk/K_r0_reg_n_0_[25] ),
        .O(\u1/u1/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__138_i_2
       (.I0(\u1/R0 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r0_reg_n_0_[55] ),
        .I3(\u1/uk/p_6_in ),
        .O(\u1/u1/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__138_i_3
       (.I0(\u1/R0 [6]),
        .I1(decrypt),
        .I2(\u1/uk/K_r0_reg_n_0_[4] ),
        .I3(\u1/uk/p_8_in ),
        .O(\u1/u1/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__138_i_4
       (.I0(\u1/R0 [5]),
        .I1(decrypt),
        .I2(\u1/uk/p_7_in ),
        .I3(\u1/uk/K_r0_reg_n_0_[17] ),
        .O(\u1/u1/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__138_i_5
       (.I0(\u1/R0 [9]),
        .I1(decrypt),
        .I2(\u1/uk/p_9_in ),
        .I3(\u1/uk/p_10_in ),
        .O(\u1/u1/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__138_i_6
       (.I0(\u1/R0 [4]),
        .I1(decrypt),
        .I2(\u1/uk/p_6_in ),
        .I3(\u1/uk/p_7_in ),
        .O(\u1/u1/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__139
       (.I0(\u1/u1/X [47]),
        .I1(\u1/u1/X [46]),
        .I2(\u1/u1/X [45]),
        .I3(\u1/u1/X [44]),
        .I4(\u1/u1/X [48]),
        .I5(\u1/u1/X [43]),
        .O(\u1/out1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__139_i_1
       (.I0(\u1/R0 [32]),
        .I1(decrypt),
        .I2(\u1/uk/p_36_in ),
        .I3(\u1/uk/K_r0_reg_n_0_[52] ),
        .O(\u1/u1/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__139_i_2
       (.I0(\u1/R0 [31]),
        .I1(decrypt),
        .I2(\u1/uk/p_32_in ),
        .I3(\u1/uk/p_29_in ),
        .O(\u1/u1/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__139_i_3
       (.I0(\u1/R0 [30]),
        .I1(decrypt),
        .I2(\u1/uk/p_35_in ),
        .I3(\u1/uk/p_22_in ),
        .O(\u1/u1/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__139_i_4
       (.I0(\u1/R0 [29]),
        .I1(decrypt),
        .I2(\u1/uk/p_28_in ),
        .I3(\u1/uk/p_31_in ),
        .O(\u1/u1/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__139_i_5
       (.I0(\u1/R0 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r0_reg_n_0_[35] ),
        .I3(\u1/uk/p_36_in ),
        .O(\u1/u1/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__139_i_6
       (.I0(\u1/R0 [28]),
        .I1(decrypt),
        .I2(\u1/uk/p_30_in ),
        .I3(\u1/uk/K_r0_reg_n_0_[2] ),
        .O(\u1/u1/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__13_i_1
       (.I0(\u0/R0 [20]),
        .I1(decrypt),
        .I2(\u0/uk/p_22_in ),
        .I3(\u0/uk/p_23_in ),
        .O(\u0/u1/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__13_i_2
       (.I0(\u0/R0 [19]),
        .I1(decrypt),
        .I2(\u0/uk/p_25_in ),
        .I3(\u0/uk/p_34_in ),
        .O(\u0/u1/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__13_i_3
       (.I0(\u0/R0 [18]),
        .I1(decrypt),
        .I2(\u0/uk/p_20_in ),
        .I3(\u0/uk/p_21_in ),
        .O(\u0/u1/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__13_i_4
       (.I0(\u0/R0 [17]),
        .I1(decrypt),
        .I2(\u0/uk/p_18_in ),
        .I3(\u0/uk/p_19_in ),
        .O(\u0/u1/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__13_i_5
       (.I0(\u0/R0 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r0_reg_n_0_ ),
        .I3(\u0/uk/p_18_in ),
        .O(\u0/u1/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__13_i_6
       (.I0(\u0/R0 [16]),
        .I1(decrypt),
        .I2(\u0/uk/p_17_in ),
        .I3(\u0/uk/K_r0_reg_n_0_[22] ),
        .O(\u0/u1/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__14
       (.I0(\u0/u1/X [5]),
        .I1(\u0/u1/X [4]),
        .I2(\u0/u1/X [3]),
        .I3(\u0/u1/X [2]),
        .I4(\u0/u1/X [6]),
        .I5(\u0/u1/X [1]),
        .O(\u0/out1 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__140
       (.I0(\u1/u1/X [23]),
        .I1(\u1/u1/X [22]),
        .I2(\u1/u1/X [21]),
        .I3(\u1/u1/X [20]),
        .I4(\u1/u1/X [24]),
        .I5(\u1/u1/X [19]),
        .O(\u1/out1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__140_i_1
       (.I0(\u1/R0 [16]),
        .I1(decrypt),
        .I2(\u1/uk/p_15_in ),
        .I3(\u1/uk/p_9_in ),
        .O(\u1/u1/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__140_i_2
       (.I0(\u1/R0 [15]),
        .I1(decrypt),
        .I2(\u1/uk/p_12_in ),
        .I3(\u1/uk/p_37_in ),
        .O(\u1/u1/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__140_i_3
       (.I0(\u1/R0 [14]),
        .I1(decrypt),
        .I2(\u1/uk/p_16_in ),
        .I3(\u1/uk/p_0_in ),
        .O(\u1/u1/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__140_i_4
       (.I0(\u1/R0 [13]),
        .I1(decrypt),
        .I2(\u1/uk/p_10_in ),
        .I3(\u1/uk/p_13_in ),
        .O(\u1/u1/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__140_i_5
       (.I0(\u1/R0 [17]),
        .I1(decrypt),
        .I2(\u1/uk/p_5_in ),
        .I3(\u1/uk/p_16_in ),
        .O(\u1/u1/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__140_i_6
       (.I0(\u1/R0 [12]),
        .I1(decrypt),
        .I2(\u1/uk/p_14_in ),
        .I3(\u1/uk/p_15_in ),
        .O(\u1/u1/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__141
       (.I0(\u1/u1/X [29]),
        .I1(\u1/u1/X [28]),
        .I2(\u1/u1/X [27]),
        .I3(\u1/u1/X [26]),
        .I4(\u1/u1/X [30]),
        .I5(\u1/u1/X [25]),
        .O(\u1/out1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__141_i_1
       (.I0(\u1/R0 [20]),
        .I1(decrypt),
        .I2(\u1/uk/p_22_in ),
        .I3(\u1/uk/p_23_in ),
        .O(\u1/u1/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__141_i_2
       (.I0(\u1/R0 [19]),
        .I1(decrypt),
        .I2(\u1/uk/p_25_in ),
        .I3(\u1/uk/p_34_in ),
        .O(\u1/u1/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__141_i_3
       (.I0(\u1/R0 [18]),
        .I1(decrypt),
        .I2(\u1/uk/p_20_in ),
        .I3(\u1/uk/p_21_in ),
        .O(\u1/u1/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__141_i_4
       (.I0(\u1/R0 [17]),
        .I1(decrypt),
        .I2(\u1/uk/p_18_in ),
        .I3(\u1/uk/p_19_in ),
        .O(\u1/u1/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__141_i_5
       (.I0(\u1/R0 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r0_reg_n_0_ ),
        .I3(\u1/uk/p_18_in ),
        .O(\u1/u1/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__141_i_6
       (.I0(\u1/R0 [16]),
        .I1(decrypt),
        .I2(\u1/uk/p_17_in ),
        .I3(\u1/uk/K_r0_reg_n_0_[22] ),
        .O(\u1/u1/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__142
       (.I0(\u1/u1/X [5]),
        .I1(\u1/u1/X [4]),
        .I2(\u1/u1/X [3]),
        .I3(\u1/u1/X [2]),
        .I4(\u1/u1/X [6]),
        .I5(\u1/u1/X [1]),
        .O(\u1/out1 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__142_i_1
       (.I0(\u1/R0 [4]),
        .I1(decrypt),
        .I2(\u1/uk/p_2_in ),
        .I3(\u1/uk/p_3_in ),
        .O(\u1/u1/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__142_i_2
       (.I0(\u1/R0 [3]),
        .I1(decrypt),
        .I2(\u1/uk/p_0_in ),
        .I3(\u1/uk/p_1_in ),
        .O(\u1/u1/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__142_i_3
       (.I0(\u1/R0 [2]),
        .I1(decrypt),
        .I2(\u1/uk/p_39_in ),
        .I3(\u1/uk/p_38_in ),
        .O(\u1/u1/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__142_i_4
       (.I0(\u1/R0 [1]),
        .I1(decrypt),
        .I2(\u1/uk/p_37_in ),
        .I3(\u1/uk/p_40_in ),
        .O(\u1/u1/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__142_i_5
       (.I0(\u1/R0 [5]),
        .I1(decrypt),
        .I2(\u1/uk/p_4_in ),
        .I3(\u1/uk/p_5_in ),
        .O(\u1/u1/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__142_i_6
       (.I0(\u1/R0 [32]),
        .I1(decrypt),
        .I2(\u1/uk/p_40_in ),
        .I3(\u1/uk/p_39_in ),
        .O(\u1/u1/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__143
       (.I0(\u1/u2/X [41]),
        .I1(\u1/u2/X [40]),
        .I2(\u1/u2/X [39]),
        .I3(\u1/u2/X [38]),
        .I4(\u1/u2/X [42]),
        .I5(\u1/u2/X [37]),
        .O(\u1/out2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__143_i_1
       (.I0(\u1/R1 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [8]),
        .I3(\u1/uk/K_r1 [14]),
        .O(\u1/u2/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__143_i_2
       (.I0(\u1/R1 [27]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [21]),
        .I3(\u1/uk/K_r1 [31]),
        .O(\u1/u2/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__143_i_3
       (.I0(\u1/R1 [26]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [43]),
        .I3(\u1/uk/K_r1 [49]),
        .O(\u1/u2/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__143_i_4
       (.I0(\u1/R1 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [31]),
        .I3(\u1/uk/K_r1 [9]),
        .O(\u1/u2/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__143_i_5
       (.I0(\u1/R1 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [0]),
        .I3(\u1/uk/K_r1 [37]),
        .O(\u1/u2/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__143_i_6
       (.I0(\u1/R1 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [23]),
        .I3(\u1/uk/K_r1 [29]),
        .O(\u1/u2/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__144
       (.I0(\u1/u2/X [17]),
        .I1(\u1/u2/X [16]),
        .I2(\u1/u2/X [15]),
        .I3(\u1/u2/X [14]),
        .I4(\u1/u2/X [18]),
        .I5(\u1/u2/X [13]),
        .O(\u1/out2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__144_i_1
       (.I0(\u1/R1 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [13]),
        .I3(\u1/uk/K_r1 [46]),
        .O(\u1/u2/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__144_i_2
       (.I0(\u1/R1 [11]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [55]),
        .I3(\u1/uk/K_r1 [6]),
        .O(\u1/u2/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__144_i_3
       (.I0(\u1/R1 [10]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [54]),
        .I3(\u1/uk/K_r1 [5]),
        .O(\u1/u2/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__144_i_4
       (.I0(\u1/R1 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [46]),
        .I3(\u1/uk/K_r1 [54]),
        .O(\u1/u2/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__144_i_5
       (.I0(\u1/R1 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [26]),
        .I3(\u1/uk/K_r1 [34]),
        .O(\u1/u2/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__144_i_6
       (.I0(\u1/R1 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [17]),
        .I3(\u1/uk/K_r1 [25]),
        .O(\u1/u2/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__145
       (.I0(\u1/u2/X [35]),
        .I1(\u1/u2/X [34]),
        .I2(\u1/u2/X [33]),
        .I3(\u1/u2/X [32]),
        .I4(\u1/u2/X [36]),
        .I5(\u1/u2/X [31]),
        .O(\u1/out2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__145_i_1
       (.I0(\u1/R1 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [1]),
        .I3(\u1/uk/K_r1 [7]),
        .O(\u1/u2/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__145_i_2
       (.I0(\u1/R1 [23]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [30]),
        .I3(\u1/uk/K_r1 [36]),
        .O(\u1/u2/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__145_i_3
       (.I0(\u1/R1 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [45]),
        .I3(\u1/uk/K_r1 [23]),
        .O(\u1/u2/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__145_i_4
       (.I0(\u1/R1 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [50]),
        .I3(\u1/uk/K_r1 [1]),
        .O(\u1/u2/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__145_i_5
       (.I0(\u1/R1 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [51]),
        .I3(\u1/uk/K_r1 [2]),
        .O(\u1/u2/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__145_i_6
       (.I0(\u1/R1 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [35]),
        .I3(\u1/uk/K_r1 [45]),
        .O(\u1/u2/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__146
       (.I0(\u1/u2/X [11]),
        .I1(\u1/u2/X [10]),
        .I2(\u1/u2/X [9]),
        .I3(\u1/u2/X [8]),
        .I4(\u1/u2/X [12]),
        .I5(\u1/u2/X [7]),
        .O(\u1/out2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__146_i_1
       (.I0(\u1/R1 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [3]),
        .I3(\u1/uk/K_r1 [11]),
        .O(\u1/u2/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__146_i_2
       (.I0(\u1/R1 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [12]),
        .I3(\u1/uk/K_r1 [20]),
        .O(\u1/u2/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__146_i_3
       (.I0(\u1/R1 [6]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [18]),
        .I3(\u1/uk/K_r1 [26]),
        .O(\u1/u2/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__146_i_4
       (.I0(\u1/R1 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [27]),
        .I3(\u1/uk/K_r1 [3]),
        .O(\u1/u2/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__146_i_5
       (.I0(\u1/R1 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [40]),
        .I3(\u1/uk/K_r1 [48]),
        .O(\u1/u2/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__146_i_6
       (.I0(\u1/R1 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [48]),
        .I3(\u1/uk/K_r1 [24]),
        .O(\u1/u2/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__147
       (.I0(\u1/u2/X [47]),
        .I1(\u1/u2/X [46]),
        .I2(\u1/u2/X [45]),
        .I3(\u1/u2/X [44]),
        .I4(\u1/u2/X [48]),
        .I5(\u1/u2/X [43]),
        .O(\u1/out2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__147_i_1
       (.I0(\u1/R1 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [28]),
        .I3(\u1/uk/K_r1 [38]),
        .O(\u1/u2/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__147_i_2
       (.I0(\u1/R1 [31]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [22]),
        .I3(\u1/uk/K_r1 [28]),
        .O(\u1/u2/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__147_i_3
       (.I0(\u1/R1 [30]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [38]),
        .I3(\u1/uk/K_r1 [16]),
        .O(\u1/u2/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__147_i_4
       (.I0(\u1/R1 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [9]),
        .I3(\u1/uk/K_r1 [15]),
        .O(\u1/u2/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__147_i_5
       (.I0(\u1/R1 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [49]),
        .I3(\u1/uk/K_r1 [0]),
        .O(\u1/u2/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__147_i_6
       (.I0(\u1/R1 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [37]),
        .I3(\u1/uk/K_r1 [43]),
        .O(\u1/u2/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__148
       (.I0(\u1/u2/X [23]),
        .I1(\u1/u2/X [22]),
        .I2(\u1/u2/X [21]),
        .I3(\u1/u2/X [20]),
        .I4(\u1/u2/X [24]),
        .I5(\u1/u2/X [19]),
        .O(\u1/out2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__148_i_1
       (.I0(\u1/R1 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [4]),
        .I3(\u1/uk/K_r1 [12]),
        .O(\u1/u2/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__148_i_2
       (.I0(\u1/R1 [15]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [53]),
        .I3(\u1/uk/K_r1 [4]),
        .O(\u1/u2/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__148_i_3
       (.I0(\u1/R1 [14]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [20]),
        .I3(\u1/uk/K_r1 [53]),
        .O(\u1/u2/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__148_i_4
       (.I0(\u1/R1 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [19]),
        .I3(\u1/uk/K_r1 [27]),
        .O(\u1/u2/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__148_i_5
       (.I0(\u1/R1 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [41]),
        .I3(\u1/uk/K_r1 [17]),
        .O(\u1/u2/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__148_i_6
       (.I0(\u1/R1 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [25]),
        .I3(\u1/uk/K_r1 [33]),
        .O(\u1/u2/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__149
       (.I0(\u1/u2/X [29]),
        .I1(\u1/u2/X [28]),
        .I2(\u1/u2/X [27]),
        .I3(\u1/u2/X [26]),
        .I4(\u1/u2/X [30]),
        .I5(\u1/u2/X [25]),
        .O(\u1/out2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__149_i_1
       (.I0(\u1/R1 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [44]),
        .I3(\u1/uk/K_r1 [50]),
        .O(\u1/u2/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__149_i_2
       (.I0(\u1/R1 [19]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [29]),
        .I3(\u1/uk/K_r1 [35]),
        .O(\u1/u2/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__149_i_3
       (.I0(\u1/R1 [18]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [42]),
        .I3(\u1/uk/K_r1 [52]),
        .O(\u1/u2/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__149_i_4
       (.I0(\u1/R1 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [52]),
        .I3(\u1/uk/K_r1 [30]),
        .O(\u1/u2/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__149_i_5
       (.I0(\u1/R1 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [14]),
        .I3(\u1/uk/K_r1 [51]),
        .O(\u1/u2/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__149_i_6
       (.I0(\u1/R1 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [2]),
        .I3(\u1/uk/K_r1 [8]),
        .O(\u1/u2/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__14_i_1
       (.I0(\u0/R0 [4]),
        .I1(decrypt),
        .I2(\u0/uk/p_2_in ),
        .I3(\u0/uk/p_3_in ),
        .O(\u0/u1/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__14_i_2
       (.I0(\u0/R0 [3]),
        .I1(decrypt),
        .I2(\u0/uk/p_0_in ),
        .I3(\u0/uk/p_1_in ),
        .O(\u0/u1/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__14_i_3
       (.I0(\u0/R0 [2]),
        .I1(decrypt),
        .I2(\u0/uk/p_39_in ),
        .I3(\u0/uk/p_38_in ),
        .O(\u0/u1/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__14_i_4
       (.I0(\u0/R0 [1]),
        .I1(decrypt),
        .I2(\u0/uk/p_37_in ),
        .I3(\u0/uk/p_40_in ),
        .O(\u0/u1/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__14_i_5
       (.I0(\u0/R0 [5]),
        .I1(decrypt),
        .I2(\u0/uk/p_4_in ),
        .I3(\u0/uk/p_5_in ),
        .O(\u0/u1/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__14_i_6
       (.I0(\u0/R0 [32]),
        .I1(decrypt),
        .I2(\u0/uk/p_40_in ),
        .I3(\u0/uk/p_39_in ),
        .O(\u0/u1/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__15
       (.I0(\u0/u2/X [41]),
        .I1(\u0/u2/X [40]),
        .I2(\u0/u2/X [39]),
        .I3(\u0/u2/X [38]),
        .I4(\u0/u2/X [42]),
        .I5(\u0/u2/X [37]),
        .O(\u0/out2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__150
       (.I0(\u1/u2/X [5]),
        .I1(\u1/u2/X [4]),
        .I2(\u1/u2/X [3]),
        .I3(\u1/u2/X [2]),
        .I4(\u1/u2/X [6]),
        .I5(\u1/u2/X [1]),
        .O(\u1/out2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__150_i_1
       (.I0(\u1/R1 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [34]),
        .I3(\u1/uk/K_r1 [10]),
        .O(\u1/u2/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__150_i_2
       (.I0(\u1/R1 [3]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [24]),
        .I3(\u1/uk/K_r1 [32]),
        .O(\u1/u2/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__150_i_3
       (.I0(\u1/R1 [2]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [47]),
        .I3(\u1/uk/K_r1 [55]),
        .O(\u1/u2/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__150_i_4
       (.I0(\u1/R1 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [32]),
        .I3(\u1/uk/K_r1 [40]),
        .O(\u1/u2/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__150_i_5
       (.I0(\u1/R1 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [5]),
        .I3(\u1/uk/K_r1 [13]),
        .O(\u1/u2/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__150_i_6
       (.I0(\u1/R1 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r1 [11]),
        .I3(\u1/uk/K_r1 [19]),
        .O(\u1/u2/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__151
       (.I0(\u1/u3/X [41]),
        .I1(\u1/u3/X [40]),
        .I2(\u1/u3/X [39]),
        .I3(\u1/u3/X [38]),
        .I4(\u1/u3/X [42]),
        .I5(\u1/u3/X [37]),
        .O(\u1/out3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__151_i_1
       (.I0(\u1/R2 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [22]),
        .I3(\u1/uk/K_r2 [0]),
        .O(\u1/u3/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__151_i_2
       (.I0(\u1/R2 [27]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [35]),
        .I3(\u1/uk/K_r2 [44]),
        .O(\u1/u3/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__151_i_3
       (.I0(\u1/R2 [26]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [2]),
        .I3(\u1/uk/K_r2 [35]),
        .O(\u1/u3/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__151_i_4
       (.I0(\u1/R2 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [45]),
        .I3(\u1/uk/K_r2 [50]),
        .O(\u1/u3/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__151_i_5
       (.I0(\u1/R2 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [14]),
        .I3(\u1/uk/K_r2 [23]),
        .O(\u1/u3/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__151_i_6
       (.I0(\u1/R2 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [37]),
        .I3(\u1/uk/K_r2 [15]),
        .O(\u1/u3/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__152
       (.I0(\u1/u3/X [17]),
        .I1(\u1/u3/X [16]),
        .I2(\u1/u3/X [15]),
        .I3(\u1/u3/X [14]),
        .I4(\u1/u3/X [18]),
        .I5(\u1/u3/X [13]),
        .O(\u1/out3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__152_i_1
       (.I0(\u1/R2 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [27]),
        .I3(\u1/uk/K_r2 [32]),
        .O(\u1/u3/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__152_i_2
       (.I0(\u1/R2 [11]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [12]),
        .I3(\u1/uk/K_r2 [17]),
        .O(\u1/u3/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__152_i_3
       (.I0(\u1/R2 [10]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [11]),
        .I3(\u1/uk/K_r2 [48]),
        .O(\u1/u3/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__152_i_4
       (.I0(\u1/R2 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [3]),
        .I3(\u1/uk/K_r2 [40]),
        .O(\u1/u3/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__152_i_5
       (.I0(\u1/R2 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [40]),
        .I3(\u1/uk/K_r2 [20]),
        .O(\u1/u3/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__152_i_6
       (.I0(\u1/R2 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [6]),
        .I3(\u1/uk/K_r2 [11]),
        .O(\u1/u3/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__153
       (.I0(\u1/u3/X [35]),
        .I1(\u1/u3/X [34]),
        .I2(\u1/u3/X [33]),
        .I3(\u1/u3/X [32]),
        .I4(\u1/u3/X [36]),
        .I5(\u1/u3/X [31]),
        .O(\u1/out3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__153_i_1
       (.I0(\u1/R2 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [15]),
        .I3(\u1/uk/K_r2 [52]),
        .O(\u1/u3/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__153_i_2
       (.I0(\u1/R2 [23]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [44]),
        .I3(\u1/uk/K_r2 [22]),
        .O(\u1/u3/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__153_i_3
       (.I0(\u1/R2 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [0]),
        .I3(\u1/uk/K_r2 [9]),
        .O(\u1/u3/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__153_i_4
       (.I0(\u1/R2 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [9]),
        .I3(\u1/uk/K_r2 [42]),
        .O(\u1/u3/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__153_i_5
       (.I0(\u1/R2 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [38]),
        .I3(\u1/uk/K_r2 [43]),
        .O(\u1/u3/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__153_i_6
       (.I0(\u1/R2 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [49]),
        .I3(\u1/uk/K_r2 [31]),
        .O(\u1/u3/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__154
       (.I0(\u1/u3/X [11]),
        .I1(\u1/u3/X [10]),
        .I2(\u1/u3/X [9]),
        .I3(\u1/u3/X [8]),
        .I4(\u1/u3/X [12]),
        .I5(\u1/u3/X [7]),
        .O(\u1/out3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__154_i_1
       (.I0(\u1/R2 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [17]),
        .I3(\u1/uk/K_r2 [54]),
        .O(\u1/u3/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__154_i_2
       (.I0(\u1/R2 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [26]),
        .I3(\u1/uk/K_r2 [6]),
        .O(\u1/u3/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__154_i_3
       (.I0(\u1/R2 [6]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [32]),
        .I3(\u1/uk/K_r2 [12]),
        .O(\u1/u3/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__154_i_4
       (.I0(\u1/R2 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [41]),
        .I3(\u1/uk/K_r2 [46]),
        .O(\u1/u3/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__154_i_5
       (.I0(\u1/R2 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [54]),
        .I3(\u1/uk/K_r2 [34]),
        .O(\u1/u3/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__154_i_6
       (.I0(\u1/R2 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [5]),
        .I3(\u1/uk/K_r2 [10]),
        .O(\u1/u3/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__155
       (.I0(\u1/u3/X [47]),
        .I1(\u1/u3/X [46]),
        .I2(\u1/u3/X [45]),
        .I3(\u1/u3/X [44]),
        .I4(\u1/u3/X [48]),
        .I5(\u1/u3/X [43]),
        .O(\u1/out3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__155_i_1
       (.I0(\u1/R2 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [42]),
        .I3(\u1/uk/K_r2 [51]),
        .O(\u1/u3/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__155_i_2
       (.I0(\u1/R2 [31]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [36]),
        .I3(\u1/uk/K_r2 [14]),
        .O(\u1/u3/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__155_i_3
       (.I0(\u1/R2 [30]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [52]),
        .I3(\u1/uk/K_r2 [2]),
        .O(\u1/u3/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__155_i_4
       (.I0(\u1/R2 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [23]),
        .I3(\u1/uk/K_r2 [1]),
        .O(\u1/u3/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__155_i_5
       (.I0(\u1/R2 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [8]),
        .I3(\u1/uk/K_r2 [45]),
        .O(\u1/u3/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__155_i_6
       (.I0(\u1/R2 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [51]),
        .I3(\u1/uk/K_r2 [29]),
        .O(\u1/u3/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__156
       (.I0(\u1/u3/X [23]),
        .I1(\u1/u3/X [22]),
        .I2(\u1/u3/X [21]),
        .I3(\u1/u3/X [20]),
        .I4(\u1/u3/X [24]),
        .I5(\u1/u3/X [19]),
        .O(\u1/out3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__156_i_1
       (.I0(\u1/R2 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [18]),
        .I3(\u1/uk/K_r2 [55]),
        .O(\u1/u3/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__156_i_2
       (.I0(\u1/R2 [15]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [10]),
        .I3(\u1/uk/K_r2 [47]),
        .O(\u1/u3/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__156_i_3
       (.I0(\u1/R2 [14]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [34]),
        .I3(\u1/uk/K_r2 [39]),
        .O(\u1/u3/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__156_i_4
       (.I0(\u1/R2 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [33]),
        .I3(\u1/uk/K_r2 [13]),
        .O(\u1/u3/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__156_i_5
       (.I0(\u1/R2 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [55]),
        .I3(\u1/uk/K_r2 [3]),
        .O(\u1/u3/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__156_i_6
       (.I0(\u1/R2 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [39]),
        .I3(\u1/uk/K_r2 [19]),
        .O(\u1/u3/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__157
       (.I0(\u1/u3/X [29]),
        .I1(\u1/u3/X [28]),
        .I2(\u1/u3/X [27]),
        .I3(\u1/u3/X [26]),
        .I4(\u1/u3/X [30]),
        .I5(\u1/u3/X [25]),
        .O(\u1/out3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__157_i_1
       (.I0(\u1/R2 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [31]),
        .I3(\u1/uk/K_r2 [36]),
        .O(\u1/u3/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__157_i_2
       (.I0(\u1/R2 [19]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [43]),
        .I3(\u1/uk/K_r2 [21]),
        .O(\u1/u3/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__157_i_3
       (.I0(\u1/R2 [18]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [1]),
        .I3(\u1/uk/K_r2 [38]),
        .O(\u1/u3/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__157_i_4
       (.I0(\u1/R2 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [7]),
        .I3(\u1/uk/K_r2 [16]),
        .O(\u1/u3/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__157_i_5
       (.I0(\u1/R2 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [28]),
        .I3(\u1/uk/K_r2 [37]),
        .O(\u1/u3/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__157_i_6
       (.I0(\u1/R2 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [16]),
        .I3(\u1/uk/K_r2 [49]),
        .O(\u1/u3/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__158
       (.I0(\u1/u3/X [5]),
        .I1(\u1/u3/X [4]),
        .I2(\u1/u3/X [3]),
        .I3(\u1/u3/X [2]),
        .I4(\u1/u3/X [6]),
        .I5(\u1/u3/X [1]),
        .O(\u1/out3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__158_i_1
       (.I0(\u1/R2 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [48]),
        .I3(\u1/uk/K_r2 [53]),
        .O(\u1/u3/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__158_i_2
       (.I0(\u1/R2 [3]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [13]),
        .I3(\u1/uk/K_r2 [18]),
        .O(\u1/u3/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__158_i_3
       (.I0(\u1/R2 [2]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [4]),
        .I3(\u1/uk/K_r2 [41]),
        .O(\u1/u3/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__158_i_4
       (.I0(\u1/R2 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [46]),
        .I3(\u1/uk/K_r2 [26]),
        .O(\u1/u3/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__158_i_5
       (.I0(\u1/R2 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [19]),
        .I3(\u1/uk/K_r2 [24]),
        .O(\u1/u3/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__158_i_6
       (.I0(\u1/R2 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r2 [25]),
        .I3(\u1/uk/K_r2 [5]),
        .O(\u1/u3/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__159
       (.I0(\u1/u4/X [41]),
        .I1(\u1/u4/X [40]),
        .I2(\u1/u4/X [39]),
        .I3(\u1/u4/X [38]),
        .I4(\u1/u4/X [42]),
        .I5(\u1/u4/X [37]),
        .O(\u1/out4 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__159_i_1
       (.I0(\u1/R3 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [36]),
        .I3(\u1/uk/K_r3 [45]),
        .O(\u1/u4/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__159_i_2
       (.I0(\u1/R3 [27]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [49]),
        .I3(\u1/uk/K_r3 [30]),
        .O(\u1/u4/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__159_i_3
       (.I0(\u1/R3 [26]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [16]),
        .I3(\u1/uk/K_r3 [21]),
        .O(\u1/u4/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__159_i_4
       (.I0(\u1/R3 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [0]),
        .I3(\u1/uk/K_r3 [36]),
        .O(\u1/u4/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__159_i_5
       (.I0(\u1/R3 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [28]),
        .I3(\u1/uk/K_r3 [9]),
        .O(\u1/u4/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__159_i_6
       (.I0(\u1/R3 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [51]),
        .I3(\u1/uk/K_r3 [1]),
        .O(\u1/u4/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__15_i_1
       (.I0(\u0/R1 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [8]),
        .I3(\u0/uk/K_r1 [14]),
        .O(\u0/u2/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__15_i_2
       (.I0(\u0/R1 [27]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [21]),
        .I3(\u0/uk/K_r1 [31]),
        .O(\u0/u2/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__15_i_3
       (.I0(\u0/R1 [26]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [43]),
        .I3(\u0/uk/K_r1 [49]),
        .O(\u0/u2/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__15_i_4
       (.I0(\u0/R1 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [31]),
        .I3(\u0/uk/K_r1 [9]),
        .O(\u0/u2/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__15_i_5
       (.I0(\u0/R1 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [0]),
        .I3(\u0/uk/K_r1 [37]),
        .O(\u0/u2/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__15_i_6
       (.I0(\u0/R1 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [23]),
        .I3(\u0/uk/K_r1 [29]),
        .O(\u0/u2/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__16
       (.I0(\u0/u2/X [17]),
        .I1(\u0/u2/X [16]),
        .I2(\u0/u2/X [15]),
        .I3(\u0/u2/X [14]),
        .I4(\u0/u2/X [18]),
        .I5(\u0/u2/X [13]),
        .O(\u0/out2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__160
       (.I0(\u1/u4/X [17]),
        .I1(\u1/u4/X [16]),
        .I2(\u1/u4/X [15]),
        .I3(\u1/u4/X [14]),
        .I4(\u1/u4/X [18]),
        .I5(\u1/u4/X [13]),
        .O(\u1/out4 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__160_i_1
       (.I0(\u1/R3 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [41]),
        .I3(\u1/uk/K_r3 [18]),
        .O(\u1/u4/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__160_i_2
       (.I0(\u1/R3 [11]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [26]),
        .I3(\u1/uk/K_r3 [3]),
        .O(\u1/u4/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__160_i_3
       (.I0(\u1/R3 [10]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [25]),
        .I3(\u1/uk/K_r3 [34]),
        .O(\u1/u4/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__160_i_4
       (.I0(\u1/R3 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [17]),
        .I3(\u1/uk/K_r3 [26]),
        .O(\u1/u4/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__160_i_5
       (.I0(\u1/R3 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [54]),
        .I3(\u1/uk/K_r3 [6]),
        .O(\u1/u4/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__160_i_6
       (.I0(\u1/R3 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [20]),
        .I3(\u1/uk/K_r3 [54]),
        .O(\u1/u4/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__161
       (.I0(\u1/u4/X [35]),
        .I1(\u1/u4/X [34]),
        .I2(\u1/u4/X [33]),
        .I3(\u1/u4/X [32]),
        .I4(\u1/u4/X [36]),
        .I5(\u1/u4/X [31]),
        .O(\u1/out4 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__161_i_1
       (.I0(\u1/R3 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [29]),
        .I3(\u1/uk/K_r3 [38]),
        .O(\u1/u4/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__161_i_2
       (.I0(\u1/R3 [23]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [31]),
        .I3(\u1/uk/K_r3 [8]),
        .O(\u1/u4/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__161_i_3
       (.I0(\u1/R3 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [14]),
        .I3(\u1/uk/K_r3 [50]),
        .O(\u1/u4/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__161_i_4
       (.I0(\u1/R3 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [23]),
        .I3(\u1/uk/K_r3 [28]),
        .O(\u1/u4/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__161_i_5
       (.I0(\u1/R3 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [52]),
        .I3(\u1/uk/K_r3 [29]),
        .O(\u1/u4/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__161_i_6
       (.I0(\u1/R3 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [8]),
        .I3(\u1/uk/K_r3 [44]),
        .O(\u1/u4/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__162
       (.I0(\u1/u4/X [11]),
        .I1(\u1/u4/X [10]),
        .I2(\u1/u4/X [9]),
        .I3(\u1/u4/X [8]),
        .I4(\u1/u4/X [12]),
        .I5(\u1/u4/X [7]),
        .O(\u1/out4 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__162_i_1
       (.I0(\u1/R3 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [6]),
        .I3(\u1/uk/K_r3 [40]),
        .O(\u1/u4/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__162_i_2
       (.I0(\u1/R3 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [40]),
        .I3(\u1/uk/K_r3 [17]),
        .O(\u1/u4/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__162_i_3
       (.I0(\u1/R3 [6]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [46]),
        .I3(\u1/uk/K_r3 [55]),
        .O(\u1/u4/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__162_i_4
       (.I0(\u1/R3 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [55]),
        .I3(\u1/uk/K_r3 [32]),
        .O(\u1/u4/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__162_i_5
       (.I0(\u1/R3 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [11]),
        .I3(\u1/uk/K_r3 [20]),
        .O(\u1/u4/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__162_i_6
       (.I0(\u1/R3 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [19]),
        .I3(\u1/uk/K_r3 [53]),
        .O(\u1/u4/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__163
       (.I0(\u1/u4/X [47]),
        .I1(\u1/u4/X [46]),
        .I2(\u1/u4/X [45]),
        .I3(\u1/u4/X [44]),
        .I4(\u1/u4/X [48]),
        .I5(\u1/u4/X [43]),
        .O(\u1/out4 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__163_i_1
       (.I0(\u1/R3 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [1]),
        .I3(\u1/uk/K_r3 [37]),
        .O(\u1/u4/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__163_i_2
       (.I0(\u1/R3 [31]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [50]),
        .I3(\u1/uk/K_r3 [0]),
        .O(\u1/u4/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__163_i_3
       (.I0(\u1/R3 [30]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [7]),
        .I3(\u1/uk/K_r3 [43]),
        .O(\u1/u4/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__163_i_4
       (.I0(\u1/R3 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [37]),
        .I3(\u1/uk/K_r3 [42]),
        .O(\u1/u4/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__163_i_5
       (.I0(\u1/R3 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [22]),
        .I3(\u1/uk/K_r3 [31]),
        .O(\u1/u4/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__163_i_6
       (.I0(\u1/R3 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [38]),
        .I3(\u1/uk/K_r3 [15]),
        .O(\u1/u4/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__164
       (.I0(\u1/u4/X [23]),
        .I1(\u1/u4/X [22]),
        .I2(\u1/u4/X [21]),
        .I3(\u1/u4/X [20]),
        .I4(\u1/u4/X [24]),
        .I5(\u1/u4/X [19]),
        .O(\u1/out4 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__164_i_1
       (.I0(\u1/R3 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [32]),
        .I3(\u1/uk/K_r3 [41]),
        .O(\u1/u4/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__164_i_2
       (.I0(\u1/R3 [15]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [24]),
        .I3(\u1/uk/K_r3 [33]),
        .O(\u1/u4/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__164_i_3
       (.I0(\u1/R3 [14]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [48]),
        .I3(\u1/uk/K_r3 [25]),
        .O(\u1/u4/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__164_i_4
       (.I0(\u1/R3 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [47]),
        .I3(\u1/uk/K_r3 [24]),
        .O(\u1/u4/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__164_i_5
       (.I0(\u1/R3 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [12]),
        .I3(\u1/uk/K_r3 [46]),
        .O(\u1/u4/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__164_i_6
       (.I0(\u1/R3 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [53]),
        .I3(\u1/uk/K_r3 [5]),
        .O(\u1/u4/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__165
       (.I0(\u1/u4/X [29]),
        .I1(\u1/u4/X [28]),
        .I2(\u1/u4/X [27]),
        .I3(\u1/u4/X [26]),
        .I4(\u1/u4/X [30]),
        .I5(\u1/u4/X [25]),
        .O(\u1/out4 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__165_i_1
       (.I0(\u1/R3 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [45]),
        .I3(\u1/uk/K_r3 [22]),
        .O(\u1/u4/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__165_i_2
       (.I0(\u1/R3 [19]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [2]),
        .I3(\u1/uk/K_r3 [7]),
        .O(\u1/u4/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__165_i_3
       (.I0(\u1/R3 [18]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [15]),
        .I3(\u1/uk/K_r3 [51]),
        .O(\u1/u4/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__165_i_4
       (.I0(\u1/R3 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [21]),
        .I3(\u1/uk/K_r3 [2]),
        .O(\u1/u4/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__165_i_5
       (.I0(\u1/R3 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [42]),
        .I3(\u1/uk/K_r3 [23]),
        .O(\u1/u4/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__165_i_6
       (.I0(\u1/R3 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [30]),
        .I3(\u1/uk/K_r3 [35]),
        .O(\u1/u4/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__166
       (.I0(\u1/u4/X [5]),
        .I1(\u1/u4/X [4]),
        .I2(\u1/u4/X [3]),
        .I3(\u1/u4/X [2]),
        .I4(\u1/u4/X [6]),
        .I5(\u1/u4/X [1]),
        .O(\u1/out4 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__166_i_1
       (.I0(\u1/R3 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [5]),
        .I3(\u1/uk/K_r3 [39]),
        .O(\u1/u4/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__166_i_2
       (.I0(\u1/R3 [3]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [27]),
        .I3(\u1/uk/K_r3 [4]),
        .O(\u1/u4/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__166_i_3
       (.I0(\u1/R3 [2]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [18]),
        .I3(\u1/uk/K_r3 [27]),
        .O(\u1/u4/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__166_i_4
       (.I0(\u1/R3 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [3]),
        .I3(\u1/uk/K_r3 [12]),
        .O(\u1/u4/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__166_i_5
       (.I0(\u1/R3 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [33]),
        .I3(\u1/uk/K_r3 [10]),
        .O(\u1/u4/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__166_i_6
       (.I0(\u1/R3 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r3 [39]),
        .I3(\u1/uk/K_r3 [48]),
        .O(\u1/u4/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__167
       (.I0(\u1/u5/X [41]),
        .I1(\u1/u5/X [40]),
        .I2(\u1/u5/X [39]),
        .I3(\u1/u5/X [38]),
        .I4(\u1/u5/X [42]),
        .I5(\u1/u5/X [37]),
        .O(\u1/out5 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__167_i_1
       (.I0(\u1/R4 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[50] ),
        .I3(\u1/uk/K_r4_reg_n_0_[31] ),
        .O(\u1/u5/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__167_i_2
       (.I0(\u1/R4 [27]),
        .I1(decrypt),
        .I2(\u1/uk/p_42_in ),
        .I3(\u1/uk/K_r4_reg_n_0_[16] ),
        .O(\u1/u5/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__167_i_3
       (.I0(\u1/R4 [26]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[30] ),
        .I3(\u1/uk/K_r4_reg_n_0_[7] ),
        .O(\u1/u5/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__167_i_4
       (.I0(\u1/R4 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[14] ),
        .I3(\u1/uk/K_r4_reg_n_0_[22] ),
        .O(\u1/u5/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__167_i_5
       (.I0(\u1/R4 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[42] ),
        .I3(\u1/uk/K_r4_reg_n_0_[50] ),
        .O(\u1/u5/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__167_i_6
       (.I0(\u1/R4 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[38] ),
        .I3(\u1/uk/K_r4_reg_n_0_[42] ),
        .O(\u1/u5/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__168
       (.I0(\u1/u5/X [17]),
        .I1(\u1/u5/X [16]),
        .I2(\u1/u5/X [15]),
        .I3(\u1/u5/X [14]),
        .I4(\u1/u5/X [18]),
        .I5(\u1/u5/X [13]),
        .O(\u1/out5 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__168_i_1
       (.I0(\u1/R4 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[55] ),
        .I3(\u1/uk/K_r4_reg_n_0_[4] ),
        .O(\u1/u5/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__168_i_2
       (.I0(\u1/R4 [11]),
        .I1(decrypt),
        .I2(\u1/uk/p_49_in ),
        .I3(\u1/uk/p_47_in ),
        .O(\u1/u5/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__168_i_3
       (.I0(\u1/R4 [10]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[39] ),
        .I3(\u1/uk/K_r4_reg_n_0_[20] ),
        .O(\u1/u5/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__168_i_4
       (.I0(\u1/R4 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[6] ),
        .I3(\u1/uk/K_r4_reg_n_0_[12] ),
        .O(\u1/u5/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__168_i_5
       (.I0(\u1/R4 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[11] ),
        .I3(\u1/uk/K_r4_reg_n_0_[17] ),
        .O(\u1/u5/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__168_i_6
       (.I0(\u1/R4 [8]),
        .I1(decrypt),
        .I2(\u1/uk/p_50_in ),
        .I3(\u1/uk/p_49_in ),
        .O(\u1/u5/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__169
       (.I0(\u1/u5/X [35]),
        .I1(\u1/u5/X [34]),
        .I2(\u1/u5/X [33]),
        .I3(\u1/u5/X [32]),
        .I4(\u1/u5/X [36]),
        .I5(\u1/u5/X [31]),
        .O(\u1/out5 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__169_i_1
       (.I0(\u1/R4 [24]),
        .I1(decrypt),
        .I2(\u1/uk/p_44_in ),
        .I3(\u1/uk/K_r4_reg_n_0_[51] ),
        .O(\u1/u5/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__169_i_2
       (.I0(\u1/R4 [23]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[45] ),
        .I3(\u1/uk/K_r4_reg_n_0_[49] ),
        .O(\u1/u5/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__169_i_3
       (.I0(\u1/R4 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[28] ),
        .I3(\u1/uk/K_r4_reg_n_0_[36] ),
        .O(\u1/u5/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__169_i_4
       (.I0(\u1/R4 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[37] ),
        .I3(\u1/uk/K_r4_reg_n_0_[14] ),
        .O(\u1/u5/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__169_i_5
       (.I0(\u1/R4 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[7] ),
        .I3(\u1/uk/K_r4_reg_n_0_[15] ),
        .O(\u1/u5/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__169_i_6
       (.I0(\u1/R4 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[22] ),
        .I3(\u1/uk/K_r4_reg_n_0_[30] ),
        .O(\u1/u5/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__16_i_1
       (.I0(\u0/R1 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [13]),
        .I3(\u0/uk/K_r1 [46]),
        .O(\u0/u2/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__16_i_2
       (.I0(\u0/R1 [11]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [55]),
        .I3(\u0/uk/K_r1 [6]),
        .O(\u0/u2/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__16_i_3
       (.I0(\u0/R1 [10]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [54]),
        .I3(\u0/uk/K_r1 [5]),
        .O(\u0/u2/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__16_i_4
       (.I0(\u0/R1 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [46]),
        .I3(\u0/uk/K_r1 [54]),
        .O(\u0/u2/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__16_i_5
       (.I0(\u0/R1 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [26]),
        .I3(\u0/uk/K_r1 [34]),
        .O(\u0/u2/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__16_i_6
       (.I0(\u0/R1 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [17]),
        .I3(\u0/uk/K_r1 [25]),
        .O(\u0/u2/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__17
       (.I0(\u0/u2/X [35]),
        .I1(\u0/u2/X [34]),
        .I2(\u0/u2/X [33]),
        .I3(\u0/u2/X [32]),
        .I4(\u0/u2/X [36]),
        .I5(\u0/u2/X [31]),
        .O(\u0/out2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__170
       (.I0(\u1/u5/X [11]),
        .I1(\u1/u5/X [10]),
        .I2(\u1/u5/X [9]),
        .I3(\u1/u5/X [8]),
        .I4(\u1/u5/X [12]),
        .I5(\u1/u5/X [7]),
        .O(\u1/out5 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__170_i_1
       (.I0(\u1/R4 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[20] ),
        .I3(\u1/uk/K_r4_reg_n_0_[26] ),
        .O(\u1/u5/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__170_i_2
       (.I0(\u1/R4 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[54] ),
        .I3(\u1/uk/K_r4_reg_n_0_[3] ),
        .O(\u1/u5/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__170_i_3
       (.I0(\u1/R4 [6]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[3] ),
        .I3(\u1/uk/K_r4_reg_n_0_[41] ),
        .O(\u1/u5/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__170_i_4
       (.I0(\u1/R4 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[12] ),
        .I3(\u1/uk/K_r4_reg_n_0_[18] ),
        .O(\u1/u5/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__170_i_5
       (.I0(\u1/R4 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[25] ),
        .I3(\u1/uk/K_r4_reg_n_0_[6] ),
        .O(\u1/u5/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__170_i_6
       (.I0(\u1/R4 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[33] ),
        .I3(\u1/uk/K_r4_reg_n_0_[39] ),
        .O(\u1/u5/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__171
       (.I0(\u1/u5/X [47]),
        .I1(\u1/u5/X [46]),
        .I2(\u1/u5/X [45]),
        .I3(\u1/u5/X [44]),
        .I4(\u1/u5/X [48]),
        .I5(\u1/u5/X [43]),
        .O(\u1/out5 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__171_i_1
       (.I0(\u1/R4 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[15] ),
        .I3(\u1/uk/K_r4_reg_n_0_[23] ),
        .O(\u1/u5/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__171_i_2
       (.I0(\u1/R4 [31]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[9] ),
        .I3(\u1/uk/K_r4_reg_n_0_[45] ),
        .O(\u1/u5/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__171_i_3
       (.I0(\u1/R4 [30]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[21] ),
        .I3(\u1/uk/K_r4_reg_n_0_[29] ),
        .O(\u1/u5/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__171_i_4
       (.I0(\u1/R4 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[51] ),
        .I3(\u1/uk/K_r4_reg_n_0_[28] ),
        .O(\u1/u5/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__171_i_5
       (.I0(\u1/R4 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[36] ),
        .I3(\u1/uk/K_r4_reg_n_0_[44] ),
        .O(\u1/u5/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__171_i_6
       (.I0(\u1/R4 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[52] ),
        .I3(\u1/uk/K_r4_reg_n_0_[1] ),
        .O(\u1/u5/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__172
       (.I0(\u1/u5/X [23]),
        .I1(\u1/u5/X [22]),
        .I2(\u1/u5/X [21]),
        .I3(\u1/u5/X [20]),
        .I4(\u1/u5/X [24]),
        .I5(\u1/u5/X [19]),
        .O(\u1/out5 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__172_i_1
       (.I0(\u1/R4 [16]),
        .I1(decrypt),
        .I2(\u1/uk/p_47_in ),
        .I3(\u1/uk/K_r4_reg_n_0_[27] ),
        .O(\u1/u5/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__172_i_2
       (.I0(\u1/R4 [15]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[13] ),
        .I3(\u1/uk/K_r4_reg_n_0_[19] ),
        .O(\u1/u5/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__172_i_3
       (.I0(\u1/R4 [14]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[5] ),
        .I3(\u1/uk/K_r4_reg_n_0_[11] ),
        .O(\u1/u5/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__172_i_4
       (.I0(\u1/R4 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[4] ),
        .I3(\u1/uk/K_r4_reg_n_0_[10] ),
        .O(\u1/u5/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__172_i_5
       (.I0(\u1/R4 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[26] ),
        .I3(\u1/uk/K_r4_reg_n_0_[32] ),
        .O(\u1/u5/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__172_i_6
       (.I0(\u1/R4 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[10] ),
        .I3(\u1/uk/K_r4_reg_n_0_[48] ),
        .O(\u1/u5/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__173
       (.I0(\u1/u5/X [29]),
        .I1(\u1/u5/X [28]),
        .I2(\u1/u5/X [27]),
        .I3(\u1/u5/X [26]),
        .I4(\u1/u5/X [30]),
        .I5(\u1/u5/X [25]),
        .O(\u1/out5 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__173_i_1
       (.I0(\u1/R4 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_ ),
        .I3(\u1/uk/p_42_in ),
        .O(\u1/u5/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__173_i_2
       (.I0(\u1/R4 [19]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[16] ),
        .I3(\u1/uk/K_r4_reg_n_0_[52] ),
        .O(\u1/u5/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__173_i_3
       (.I0(\u1/R4 [18]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[29] ),
        .I3(\u1/uk/K_r4_reg_n_0_[37] ),
        .O(\u1/u5/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__173_i_4
       (.I0(\u1/R4 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[35] ),
        .I3(\u1/uk/p_44_in ),
        .O(\u1/u5/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__173_i_5
       (.I0(\u1/R4 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[1] ),
        .I3(\u1/uk/K_r4_reg_n_0_[9] ),
        .O(\u1/u5/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__173_i_6
       (.I0(\u1/R4 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[44] ),
        .I3(\u1/uk/K_r4_reg_n_0_[21] ),
        .O(\u1/u5/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__174
       (.I0(\u1/u5/X [5]),
        .I1(\u1/u5/X [4]),
        .I2(\u1/u5/X [3]),
        .I3(\u1/u5/X [2]),
        .I4(\u1/u5/X [6]),
        .I5(\u1/u5/X [1]),
        .O(\u1/out5 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__174_i_1
       (.I0(\u1/R4 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[19] ),
        .I3(\u1/uk/K_r4_reg_n_0_[25] ),
        .O(\u1/u5/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__174_i_2
       (.I0(\u1/R4 [3]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[41] ),
        .I3(\u1/uk/K_r4_reg_n_0_[47] ),
        .O(\u1/u5/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__174_i_3
       (.I0(\u1/R4 [2]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[32] ),
        .I3(\u1/uk/K_r4_reg_n_0_[13] ),
        .O(\u1/u5/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__174_i_4
       (.I0(\u1/R4 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[17] ),
        .I3(\u1/uk/K_r4_reg_n_0_[55] ),
        .O(\u1/u5/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__174_i_5
       (.I0(\u1/R4 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r4_reg_n_0_[47] ),
        .I3(\u1/uk/p_51_in ),
        .O(\u1/u5/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__174_i_6
       (.I0(\u1/R4 [32]),
        .I1(decrypt),
        .I2(\u1/uk/p_51_in ),
        .I3(\u1/uk/p_50_in ),
        .O(\u1/u5/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__175
       (.I0(\u1/u6/X [41]),
        .I1(\u1/u6/X [40]),
        .I2(\u1/u6/X [39]),
        .I3(\u1/u6/X [38]),
        .I4(\u1/u6/X [42]),
        .I5(\u1/u6/X [37]),
        .O(\u1/out6 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__175_i_1
       (.I0(\u1/R5 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [9]),
        .I3(\u1/uk/K_r5 [44]),
        .O(\u1/u6/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__175_i_2
       (.I0(\u1/R5 [27]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [22]),
        .I3(\u1/uk/K_r5 [2]),
        .O(\u1/u6/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__175_i_3
       (.I0(\u1/R5 [26]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [44]),
        .I3(\u1/uk/K_r5 [52]),
        .O(\u1/u6/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__175_i_4
       (.I0(\u1/R5 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [28]),
        .I3(\u1/uk/K_r5 [8]),
        .O(\u1/u6/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__175_i_5
       (.I0(\u1/R5 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [1]),
        .I3(\u1/uk/K_r5 [36]),
        .O(\u1/u6/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__175_i_6
       (.I0(\u1/R5 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [52]),
        .I3(\u1/uk/K_r5 [28]),
        .O(\u1/u6/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__176
       (.I0(\u1/u6/X [17]),
        .I1(\u1/u6/X [16]),
        .I2(\u1/u6/X [15]),
        .I3(\u1/u6/X [14]),
        .I4(\u1/u6/X [18]),
        .I5(\u1/u6/X [13]),
        .O(\u1/out6 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__176_i_1
       (.I0(\u1/R5 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [12]),
        .I3(\u1/uk/K_r5 [47]),
        .O(\u1/u6/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__176_i_2
       (.I0(\u1/R5 [11]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [54]),
        .I3(\u1/uk/K_r5 [32]),
        .O(\u1/u6/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__176_i_3
       (.I0(\u1/R5 [10]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [53]),
        .I3(\u1/uk/K_r5 [6]),
        .O(\u1/u6/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__176_i_4
       (.I0(\u1/R5 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [20]),
        .I3(\u1/uk/K_r5 [55]),
        .O(\u1/u6/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__176_i_5
       (.I0(\u1/R5 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [25]),
        .I3(\u1/uk/K_r5 [3]),
        .O(\u1/u6/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__176_i_6
       (.I0(\u1/R5 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [48]),
        .I3(\u1/uk/K_r5 [26]),
        .O(\u1/u6/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__177
       (.I0(\u1/u6/X [35]),
        .I1(\u1/u6/X [34]),
        .I2(\u1/u6/X [33]),
        .I3(\u1/u6/X [32]),
        .I4(\u1/u6/X [36]),
        .I5(\u1/u6/X [31]),
        .O(\u1/out6 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__177_i_1
       (.I0(\u1/R5 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [2]),
        .I3(\u1/uk/K_r5 [37]),
        .O(\u1/u6/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__177_i_2
       (.I0(\u1/R5 [23]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [0]),
        .I3(\u1/uk/K_r5 [35]),
        .O(\u1/u6/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__177_i_3
       (.I0(\u1/R5 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [42]),
        .I3(\u1/uk/K_r5 [22]),
        .O(\u1/u6/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__177_i_4
       (.I0(\u1/R5 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [51]),
        .I3(\u1/uk/K_r5 [0]),
        .O(\u1/u6/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__177_i_5
       (.I0(\u1/R5 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [21]),
        .I3(\u1/uk/K_r5 [1]),
        .O(\u1/u6/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__177_i_6
       (.I0(\u1/R5 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [36]),
        .I3(\u1/uk/K_r5 [16]),
        .O(\u1/u6/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__178
       (.I0(\u1/u6/X [11]),
        .I1(\u1/u6/X [10]),
        .I2(\u1/u6/X [9]),
        .I3(\u1/u6/X [8]),
        .I4(\u1/u6/X [12]),
        .I5(\u1/u6/X [7]),
        .O(\u1/out6 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__178_i_1
       (.I0(\u1/R5 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [34]),
        .I3(\u1/uk/K_r5 [12]),
        .O(\u1/u6/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__178_i_2
       (.I0(\u1/R5 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [11]),
        .I3(\u1/uk/K_r5 [46]),
        .O(\u1/u6/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__178_i_3
       (.I0(\u1/R5 [6]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [17]),
        .I3(\u1/uk/K_r5 [27]),
        .O(\u1/u6/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__178_i_4
       (.I0(\u1/R5 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [26]),
        .I3(\u1/uk/K_r5 [4]),
        .O(\u1/u6/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__178_i_5
       (.I0(\u1/R5 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [39]),
        .I3(\u1/uk/K_r5 [17]),
        .O(\u1/u6/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__178_i_6
       (.I0(\u1/R5 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [47]),
        .I3(\u1/uk/K_r5 [25]),
        .O(\u1/u6/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__179
       (.I0(\u1/u6/X [47]),
        .I1(\u1/u6/X [46]),
        .I2(\u1/u6/X [45]),
        .I3(\u1/u6/X [44]),
        .I4(\u1/u6/X [48]),
        .I5(\u1/u6/X [43]),
        .O(\u1/out6 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__179_i_1
       (.I0(\u1/R5 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [29]),
        .I3(\u1/uk/K_r5 [9]),
        .O(\u1/u6/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__179_i_2
       (.I0(\u1/R5 [31]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [23]),
        .I3(\u1/uk/K_r5 [31]),
        .O(\u1/u6/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__179_i_3
       (.I0(\u1/R5 [30]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [35]),
        .I3(\u1/uk/K_r5 [15]),
        .O(\u1/u6/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__179_i_4
       (.I0(\u1/R5 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [38]),
        .I3(\u1/uk/K_r5 [14]),
        .O(\u1/u6/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__179_i_5
       (.I0(\u1/R5 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [50]),
        .I3(\u1/uk/K_r5 [30]),
        .O(\u1/u6/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__179_i_6
       (.I0(\u1/R5 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [7]),
        .I3(\u1/uk/K_r5 [42]),
        .O(\u1/u6/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__17_i_1
       (.I0(\u0/R1 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [1]),
        .I3(\u0/uk/K_r1 [7]),
        .O(\u0/u2/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__17_i_2
       (.I0(\u0/R1 [23]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [30]),
        .I3(\u0/uk/K_r1 [36]),
        .O(\u0/u2/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__17_i_3
       (.I0(\u0/R1 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [45]),
        .I3(\u0/uk/K_r1 [23]),
        .O(\u0/u2/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__17_i_4
       (.I0(\u0/R1 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [50]),
        .I3(\u0/uk/K_r1 [1]),
        .O(\u0/u2/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__17_i_5
       (.I0(\u0/R1 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [51]),
        .I3(\u0/uk/K_r1 [2]),
        .O(\u0/u2/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__17_i_6
       (.I0(\u0/R1 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [35]),
        .I3(\u0/uk/K_r1 [45]),
        .O(\u0/u2/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__18
       (.I0(\u0/u2/X [11]),
        .I1(\u0/u2/X [10]),
        .I2(\u0/u2/X [9]),
        .I3(\u0/u2/X [8]),
        .I4(\u0/u2/X [12]),
        .I5(\u0/u2/X [7]),
        .O(\u0/out2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__180
       (.I0(\u1/u6/X [23]),
        .I1(\u1/u6/X [22]),
        .I2(\u1/u6/X [21]),
        .I3(\u1/u6/X [20]),
        .I4(\u1/u6/X [24]),
        .I5(\u1/u6/X [19]),
        .O(\u1/out6 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__180_i_1
       (.I0(\u1/R5 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [3]),
        .I3(\u1/uk/K_r5 [13]),
        .O(\u1/u6/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__180_i_2
       (.I0(\u1/R5 [15]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [27]),
        .I3(\u1/uk/K_r5 [5]),
        .O(\u1/u6/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__180_i_3
       (.I0(\u1/R5 [14]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [19]),
        .I3(\u1/uk/K_r5 [54]),
        .O(\u1/u6/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__180_i_4
       (.I0(\u1/R5 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [18]),
        .I3(\u1/uk/K_r5 [53]),
        .O(\u1/u6/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__180_i_5
       (.I0(\u1/R5 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [40]),
        .I3(\u1/uk/K_r5 [18]),
        .O(\u1/u6/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__180_i_6
       (.I0(\u1/R5 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [24]),
        .I3(\u1/uk/K_r5 [34]),
        .O(\u1/u6/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__181
       (.I0(\u1/u6/X [29]),
        .I1(\u1/u6/X [28]),
        .I2(\u1/u6/X [27]),
        .I3(\u1/u6/X [26]),
        .I4(\u1/u6/X [30]),
        .I5(\u1/u6/X [25]),
        .O(\u1/out6 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__181_i_1
       (.I0(\u1/R5 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [14]),
        .I3(\u1/uk/K_r5 [49]),
        .O(\u1/u6/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__181_i_2
       (.I0(\u1/R5 [19]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [30]),
        .I3(\u1/uk/K_r5 [38]),
        .O(\u1/u6/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__181_i_3
       (.I0(\u1/R5 [18]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [43]),
        .I3(\u1/uk/K_r5 [23]),
        .O(\u1/u6/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__181_i_4
       (.I0(\u1/R5 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [49]),
        .I3(\u1/uk/K_r5 [29]),
        .O(\u1/u6/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__181_i_5
       (.I0(\u1/R5 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [15]),
        .I3(\u1/uk/K_r5 [50]),
        .O(\u1/u6/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__181_i_6
       (.I0(\u1/R5 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [31]),
        .I3(\u1/uk/K_r5 [7]),
        .O(\u1/u6/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__182
       (.I0(\u1/u6/X [5]),
        .I1(\u1/u6/X [4]),
        .I2(\u1/u6/X [3]),
        .I3(\u1/u6/X [2]),
        .I4(\u1/u6/X [6]),
        .I5(\u1/u6/X [1]),
        .O(\u1/out6 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__182_i_1
       (.I0(\u1/R5 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [33]),
        .I3(\u1/uk/K_r5 [11]),
        .O(\u1/u6/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__182_i_2
       (.I0(\u1/R5 [3]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [55]),
        .I3(\u1/uk/K_r5 [33]),
        .O(\u1/u6/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__182_i_3
       (.I0(\u1/R5 [2]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [46]),
        .I3(\u1/uk/K_r5 [24]),
        .O(\u1/u6/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__182_i_4
       (.I0(\u1/R5 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [6]),
        .I3(\u1/uk/K_r5 [41]),
        .O(\u1/u6/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__182_i_5
       (.I0(\u1/R5 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [4]),
        .I3(\u1/uk/K_r5 [39]),
        .O(\u1/u6/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__182_i_6
       (.I0(\u1/R5 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r5 [10]),
        .I3(\u1/uk/K_r5 [20]),
        .O(\u1/u6/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__183
       (.I0(\u1/u7/X [41]),
        .I1(\u1/u7/X [40]),
        .I2(\u1/u7/X [39]),
        .I3(\u1/u7/X [38]),
        .I4(\u1/u7/X [42]),
        .I5(\u1/u7/X [37]),
        .O(\u1/out7 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__183_i_1
       (.I0(\u1/R6 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[23] ),
        .I3(\u1/uk/K_r6_reg_n_0_[30] ),
        .O(\u1/u7/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__183_i_2
       (.I0(\u1/R6 [27]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[36] ),
        .I3(\u1/uk/p_45_in ),
        .O(\u1/u7/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__183_i_3
       (.I0(\u1/R6 [26]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[31] ),
        .I3(\u1/uk/K_r6_reg_n_0_[38] ),
        .O(\u1/u7/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__183_i_4
       (.I0(\u1/R6 [25]),
        .I1(decrypt),
        .I2(\u1/uk/p_41_in ),
        .I3(\u1/uk/p_43_in ),
        .O(\u1/u7/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__183_i_5
       (.I0(\u1/R6 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[15] ),
        .I3(\u1/uk/K_r6_reg_n_0_[22] ),
        .O(\u1/u7/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__183_i_6
       (.I0(\u1/R6 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[7] ),
        .I3(\u1/uk/K_r6_reg_n_0_[14] ),
        .O(\u1/u7/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__184
       (.I0(\u1/u7/X [17]),
        .I1(\u1/u7/X [16]),
        .I2(\u1/u7/X [15]),
        .I3(\u1/u7/X [14]),
        .I4(\u1/u7/X [18]),
        .I5(\u1/u7/X [13]),
        .O(\u1/out7 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__184_i_1
       (.I0(\u1/R6 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[26] ),
        .I3(\u1/uk/K_r6_reg_n_0_[33] ),
        .O(\u1/u7/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__184_i_2
       (.I0(\u1/R6 [11]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[11] ),
        .I3(\u1/uk/K_r6_reg_n_0_[18] ),
        .O(\u1/u7/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__184_i_3
       (.I0(\u1/R6 [10]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[10] ),
        .I3(\u1/uk/K_r6_reg_n_0_[17] ),
        .O(\u1/u7/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__184_i_4
       (.I0(\u1/R6 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[34] ),
        .I3(\u1/uk/K_r6_reg_n_0_[41] ),
        .O(\u1/u7/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__184_i_5
       (.I0(\u1/R6 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[39] ),
        .I3(\u1/uk/K_r6_reg_n_0_[46] ),
        .O(\u1/u7/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__184_i_6
       (.I0(\u1/R6 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[5] ),
        .I3(\u1/uk/K_r6_reg_n_0_[12] ),
        .O(\u1/u7/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__185
       (.I0(\u1/u7/X [35]),
        .I1(\u1/u7/X [34]),
        .I2(\u1/u7/X [33]),
        .I3(\u1/u7/X [32]),
        .I4(\u1/u7/X [36]),
        .I5(\u1/u7/X [31]),
        .O(\u1/out7 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__185_i_1
       (.I0(\u1/R6 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[16] ),
        .I3(\u1/uk/K_r6_reg_n_0_[23] ),
        .O(\u1/u7/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__185_i_2
       (.I0(\u1/R6 [23]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[14] ),
        .I3(\u1/uk/K_r6_reg_n_0_[21] ),
        .O(\u1/u7/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__185_i_3
       (.I0(\u1/R6 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[1] ),
        .I3(\u1/uk/K_r6_reg_n_0_[8] ),
        .O(\u1/u7/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__185_i_4
       (.I0(\u1/R6 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[38] ),
        .I3(\u1/uk/K_r6_reg_n_0_[45] ),
        .O(\u1/u7/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__185_i_5
       (.I0(\u1/R6 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[35] ),
        .I3(\u1/uk/p_41_in ),
        .O(\u1/u7/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__185_i_6
       (.I0(\u1/R6 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[50] ),
        .I3(\u1/uk/K_r6_reg_n_0_[2] ),
        .O(\u1/u7/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__186
       (.I0(\u1/u7/X [11]),
        .I1(\u1/u7/X [10]),
        .I2(\u1/u7/X [9]),
        .I3(\u1/u7/X [8]),
        .I4(\u1/u7/X [12]),
        .I5(\u1/u7/X [7]),
        .O(\u1/out7 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__186_i_1
       (.I0(\u1/R6 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[48] ),
        .I3(\u1/uk/K_r6_reg_n_0_[55] ),
        .O(\u1/u7/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__186_i_2
       (.I0(\u1/R6 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[25] ),
        .I3(\u1/uk/K_r6_reg_n_0_[32] ),
        .O(\u1/u7/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__186_i_3
       (.I0(\u1/R6 [6]),
        .I1(decrypt),
        .I2(\u1/uk/p_53_in ),
        .I3(\u1/uk/p_52_in ),
        .O(\u1/u7/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__186_i_4
       (.I0(\u1/R6 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[40] ),
        .I3(\u1/uk/K_r6_reg_n_0_[47] ),
        .O(\u1/u7/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__186_i_5
       (.I0(\u1/R6 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[53] ),
        .I3(\u1/uk/K_r6_reg_n_0_[3] ),
        .O(\u1/u7/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__186_i_6
       (.I0(\u1/R6 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[4] ),
        .I3(\u1/uk/K_r6_reg_n_0_[11] ),
        .O(\u1/u7/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__187
       (.I0(\u1/u7/X [47]),
        .I1(\u1/u7/X [46]),
        .I2(\u1/u7/X [45]),
        .I3(\u1/u7/X [44]),
        .I4(\u1/u7/X [48]),
        .I5(\u1/u7/X [43]),
        .O(\u1/out7 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__187_i_1
       (.I0(\u1/R6 [32]),
        .I1(decrypt),
        .I2(\u1/uk/p_45_in ),
        .I3(\u1/uk/K_r6_reg_n_0_[50] ),
        .O(\u1/u7/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__187_i_2
       (.I0(\u1/R6 [31]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[37] ),
        .I3(\u1/uk/K_r6_reg_n_0_[44] ),
        .O(\u1/u7/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__187_i_3
       (.I0(\u1/R6 [30]),
        .I1(decrypt),
        .I2(\u1/uk/p_43_in ),
        .I3(\u1/uk/K_r6_reg_n_0_[1] ),
        .O(\u1/u7/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__187_i_4
       (.I0(\u1/R6 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[52] ),
        .I3(\u1/uk/K_r6_reg_n_0_ ),
        .O(\u1/u7/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__187_i_5
       (.I0(\u1/R6 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[9] ),
        .I3(\u1/uk/K_r6_reg_n_0_[16] ),
        .O(\u1/u7/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__187_i_6
       (.I0(\u1/R6 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[21] ),
        .I3(\u1/uk/K_r6_reg_n_0_[28] ),
        .O(\u1/u7/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__188
       (.I0(\u1/u7/X [23]),
        .I1(\u1/u7/X [22]),
        .I2(\u1/u7/X [21]),
        .I3(\u1/u7/X [20]),
        .I4(\u1/u7/X [24]),
        .I5(\u1/u7/X [19]),
        .O(\u1/out7 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__188_i_1
       (.I0(\u1/R6 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[17] ),
        .I3(\u1/uk/K_r6_reg_n_0_[24] ),
        .O(\u1/u7/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__188_i_2
       (.I0(\u1/R6 [15]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[41] ),
        .I3(\u1/uk/K_r6_reg_n_0_[48] ),
        .O(\u1/u7/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__188_i_3
       (.I0(\u1/R6 [14]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[33] ),
        .I3(\u1/uk/K_r6_reg_n_0_[40] ),
        .O(\u1/u7/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__188_i_4
       (.I0(\u1/R6 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[32] ),
        .I3(\u1/uk/K_r6_reg_n_0_[39] ),
        .O(\u1/u7/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__188_i_5
       (.I0(\u1/R6 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[54] ),
        .I3(\u1/uk/K_r6_reg_n_0_[4] ),
        .O(\u1/u7/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__188_i_6
       (.I0(\u1/R6 [12]),
        .I1(decrypt),
        .I2(\u1/uk/p_52_in ),
        .I3(\u1/uk/K_r6_reg_n_0_[20] ),
        .O(\u1/u7/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__189
       (.I0(\u1/u7/X [29]),
        .I1(\u1/u7/X [28]),
        .I2(\u1/u7/X [27]),
        .I3(\u1/u7/X [26]),
        .I4(\u1/u7/X [30]),
        .I5(\u1/u7/X [25]),
        .O(\u1/out7 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__189_i_1
       (.I0(\u1/R6 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[28] ),
        .I3(\u1/uk/K_r6_reg_n_0_[35] ),
        .O(\u1/u7/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__189_i_2
       (.I0(\u1/R6 [19]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[44] ),
        .I3(\u1/uk/K_r6_reg_n_0_[51] ),
        .O(\u1/u7/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__189_i_3
       (.I0(\u1/R6 [18]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[2] ),
        .I3(\u1/uk/K_r6_reg_n_0_[9] ),
        .O(\u1/u7/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__189_i_4
       (.I0(\u1/R6 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[8] ),
        .I3(\u1/uk/K_r6_reg_n_0_[15] ),
        .O(\u1/u7/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__189_i_5
       (.I0(\u1/R6 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[29] ),
        .I3(\u1/uk/K_r6_reg_n_0_[36] ),
        .O(\u1/u7/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__189_i_6
       (.I0(\u1/R6 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[45] ),
        .I3(\u1/uk/K_r6_reg_n_0_[52] ),
        .O(\u1/u7/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__18_i_1
       (.I0(\u0/R1 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [3]),
        .I3(\u0/uk/K_r1 [11]),
        .O(\u0/u2/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__18_i_2
       (.I0(\u0/R1 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [12]),
        .I3(\u0/uk/K_r1 [20]),
        .O(\u0/u2/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__18_i_3
       (.I0(\u0/R1 [6]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [18]),
        .I3(\u0/uk/K_r1 [26]),
        .O(\u0/u2/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__18_i_4
       (.I0(\u0/R1 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [27]),
        .I3(\u0/uk/K_r1 [3]),
        .O(\u0/u2/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__18_i_5
       (.I0(\u0/R1 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [40]),
        .I3(\u0/uk/K_r1 [48]),
        .O(\u0/u2/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__18_i_6
       (.I0(\u0/R1 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [48]),
        .I3(\u0/uk/K_r1 [24]),
        .O(\u0/u2/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__19
       (.I0(\u0/u2/X [47]),
        .I1(\u0/u2/X [46]),
        .I2(\u0/u2/X [45]),
        .I3(\u0/u2/X [44]),
        .I4(\u0/u2/X [48]),
        .I5(\u0/u2/X [43]),
        .O(\u0/out2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__190
       (.I0(\u1/u7/X [5]),
        .I1(\u1/u7/X [4]),
        .I2(\u1/u7/X [3]),
        .I3(\u1/u7/X [2]),
        .I4(\u1/u7/X [6]),
        .I5(\u1/u7/X [1]),
        .O(\u1/out7 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__190_i_1
       (.I0(\u1/R6 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[47] ),
        .I3(\u1/uk/K_r6_reg_n_0_[54] ),
        .O(\u1/u7/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__190_i_2
       (.I0(\u1/R6 [3]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[12] ),
        .I3(\u1/uk/K_r6_reg_n_0_[19] ),
        .O(\u1/u7/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__190_i_3
       (.I0(\u1/R6 [2]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[3] ),
        .I3(\u1/uk/K_r6_reg_n_0_[10] ),
        .O(\u1/u7/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__190_i_4
       (.I0(\u1/R6 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[20] ),
        .I3(\u1/uk/K_r6_reg_n_0_[27] ),
        .O(\u1/u7/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__190_i_5
       (.I0(\u1/R6 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[18] ),
        .I3(\u1/uk/K_r6_reg_n_0_[25] ),
        .O(\u1/u7/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__190_i_6
       (.I0(\u1/R6 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r6_reg_n_0_[24] ),
        .I3(\u1/uk/p_53_in ),
        .O(\u1/u7/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__191
       (.I0(\u1/u8/X [41]),
        .I1(\u1/u8/X [40]),
        .I2(\u1/u8/X [39]),
        .I3(\u1/u8/X [38]),
        .I4(\u1/u8/X [42]),
        .I5(\u1/u8/X [37]),
        .O(\u1/out8 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__191_i_1
       (.I0(\u1/R7 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[30] ),
        .I3(\u1/uk/K_r7_reg_n_0_[23] ),
        .O(\u1/u8/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__191_i_2
       (.I0(\u1/R7 [27]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[43] ),
        .I3(\u1/uk/K_r7_reg_n_0_[36] ),
        .O(\u1/u8/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__191_i_3
       (.I0(\u1/R7 [26]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[38] ),
        .I3(\u1/uk/K_r7_reg_n_0_[31] ),
        .O(\u1/u8/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__191_i_4
       (.I0(\u1/R7 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[49] ),
        .I3(\u1/uk/K_r7_reg_n_0_[42] ),
        .O(\u1/u8/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__191_i_5
       (.I0(\u1/R7 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[22] ),
        .I3(\u1/uk/K_r7_reg_n_0_[15] ),
        .O(\u1/u8/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__191_i_6
       (.I0(\u1/R7 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[14] ),
        .I3(\u1/uk/K_r7_reg_n_0_[7] ),
        .O(\u1/u8/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__192
       (.I0(\u1/u8/X [17]),
        .I1(\u1/u8/X [16]),
        .I2(\u1/u8/X [15]),
        .I3(\u1/u8/X [14]),
        .I4(\u1/u8/X [18]),
        .I5(\u1/u8/X [13]),
        .O(\u1/out8 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__192_i_1
       (.I0(\u1/R7 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[33] ),
        .I3(\u1/uk/K_r7_reg_n_0_[26] ),
        .O(\u1/u8/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__192_i_2
       (.I0(\u1/R7 [11]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[18] ),
        .I3(\u1/uk/K_r7_reg_n_0_[11] ),
        .O(\u1/u8/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__192_i_3
       (.I0(\u1/R7 [10]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[17] ),
        .I3(\u1/uk/K_r7_reg_n_0_[10] ),
        .O(\u1/u8/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__192_i_4
       (.I0(\u1/R7 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[41] ),
        .I3(\u1/uk/K_r7_reg_n_0_[34] ),
        .O(\u1/u8/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__192_i_5
       (.I0(\u1/R7 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[46] ),
        .I3(\u1/uk/K_r7_reg_n_0_[39] ),
        .O(\u1/u8/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__192_i_6
       (.I0(\u1/R7 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[12] ),
        .I3(\u1/uk/K_r7_reg_n_0_[5] ),
        .O(\u1/u8/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__193
       (.I0(\u1/u8/X [35]),
        .I1(\u1/u8/X [34]),
        .I2(\u1/u8/X [33]),
        .I3(\u1/u8/X [32]),
        .I4(\u1/u8/X [36]),
        .I5(\u1/u8/X [31]),
        .O(\u1/out8 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__193_i_1
       (.I0(\u1/R7 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[23] ),
        .I3(\u1/uk/K_r7_reg_n_0_[16] ),
        .O(\u1/u8/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__193_i_2
       (.I0(\u1/R7 [23]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[21] ),
        .I3(\u1/uk/K_r7_reg_n_0_[14] ),
        .O(\u1/u8/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__193_i_3
       (.I0(\u1/R7 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[8] ),
        .I3(\u1/uk/K_r7_reg_n_0_[1] ),
        .O(\u1/u8/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__193_i_4
       (.I0(\u1/R7 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[45] ),
        .I3(\u1/uk/K_r7_reg_n_0_[38] ),
        .O(\u1/u8/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__193_i_5
       (.I0(\u1/R7 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[42] ),
        .I3(\u1/uk/K_r7_reg_n_0_[35] ),
        .O(\u1/u8/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__193_i_6
       (.I0(\u1/R7 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[2] ),
        .I3(\u1/uk/K_r7_reg_n_0_[50] ),
        .O(\u1/u8/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__194
       (.I0(\u1/u8/X [11]),
        .I1(\u1/u8/X [10]),
        .I2(\u1/u8/X [9]),
        .I3(\u1/u8/X [8]),
        .I4(\u1/u8/X [12]),
        .I5(\u1/u8/X [7]),
        .O(\u1/out8 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__194_i_1
       (.I0(\u1/R7 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[55] ),
        .I3(\u1/uk/K_r7_reg_n_0_[48] ),
        .O(\u1/u8/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__194_i_2
       (.I0(\u1/R7 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[32] ),
        .I3(\u1/uk/K_r7_reg_n_0_[25] ),
        .O(\u1/u8/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__194_i_3
       (.I0(\u1/R7 [6]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[13] ),
        .I3(\u1/uk/K_r7_reg_n_0_[6] ),
        .O(\u1/u8/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__194_i_4
       (.I0(\u1/R7 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[47] ),
        .I3(\u1/uk/K_r7_reg_n_0_[40] ),
        .O(\u1/u8/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__194_i_5
       (.I0(\u1/R7 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[3] ),
        .I3(\u1/uk/K_r7_reg_n_0_[53] ),
        .O(\u1/u8/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__194_i_6
       (.I0(\u1/R7 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[11] ),
        .I3(\u1/uk/K_r7_reg_n_0_[4] ),
        .O(\u1/u8/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__195
       (.I0(\u1/u8/X [47]),
        .I1(\u1/u8/X [46]),
        .I2(\u1/u8/X [45]),
        .I3(\u1/u8/X [44]),
        .I4(\u1/u8/X [48]),
        .I5(\u1/u8/X [43]),
        .O(\u1/out8 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__195_i_1
       (.I0(\u1/R7 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[50] ),
        .I3(\u1/uk/K_r7_reg_n_0_[43] ),
        .O(\u1/u8/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__195_i_2
       (.I0(\u1/R7 [31]),
        .I1(decrypt),
        .I2(\u1/uk/p_48_in ),
        .I3(\u1/uk/K_r7_reg_n_0_[37] ),
        .O(\u1/u8/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__195_i_3
       (.I0(\u1/R7 [30]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[1] ),
        .I3(\u1/uk/K_r7_reg_n_0_[49] ),
        .O(\u1/u8/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__195_i_4
       (.I0(\u1/R7 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_ ),
        .I3(\u1/uk/K_r7_reg_n_0_[52] ),
        .O(\u1/u8/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__195_i_5
       (.I0(\u1/R7 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[16] ),
        .I3(\u1/uk/K_r7_reg_n_0_[9] ),
        .O(\u1/u8/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__195_i_6
       (.I0(\u1/R7 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[28] ),
        .I3(\u1/uk/K_r7_reg_n_0_[21] ),
        .O(\u1/u8/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__196
       (.I0(\u1/u8/X [23]),
        .I1(\u1/u8/X [22]),
        .I2(\u1/u8/X [21]),
        .I3(\u1/u8/X [20]),
        .I4(\u1/u8/X [24]),
        .I5(\u1/u8/X [19]),
        .O(\u1/out8 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__196_i_1
       (.I0(\u1/R7 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[24] ),
        .I3(\u1/uk/K_r7_reg_n_0_[17] ),
        .O(\u1/u8/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__196_i_2
       (.I0(\u1/R7 [15]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[48] ),
        .I3(\u1/uk/K_r7_reg_n_0_[41] ),
        .O(\u1/u8/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__196_i_3
       (.I0(\u1/R7 [14]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[40] ),
        .I3(\u1/uk/K_r7_reg_n_0_[33] ),
        .O(\u1/u8/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__196_i_4
       (.I0(\u1/R7 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[39] ),
        .I3(\u1/uk/K_r7_reg_n_0_[32] ),
        .O(\u1/u8/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__196_i_5
       (.I0(\u1/R7 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[4] ),
        .I3(\u1/uk/K_r7_reg_n_0_[54] ),
        .O(\u1/u8/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__196_i_6
       (.I0(\u1/R7 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[20] ),
        .I3(\u1/uk/K_r7_reg_n_0_[13] ),
        .O(\u1/u8/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__197
       (.I0(\u1/u8/X [29]),
        .I1(\u1/u8/X [28]),
        .I2(\u1/u8/X [27]),
        .I3(\u1/u8/X [26]),
        .I4(\u1/u8/X [30]),
        .I5(\u1/u8/X [25]),
        .O(\u1/out8 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__197_i_1
       (.I0(\u1/R7 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[35] ),
        .I3(\u1/uk/K_r7_reg_n_0_[28] ),
        .O(\u1/u8/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__197_i_2
       (.I0(\u1/R7 [19]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[51] ),
        .I3(\u1/uk/p_48_in ),
        .O(\u1/u8/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__197_i_3
       (.I0(\u1/R7 [18]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[9] ),
        .I3(\u1/uk/K_r7_reg_n_0_[2] ),
        .O(\u1/u8/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__197_i_4
       (.I0(\u1/R7 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[15] ),
        .I3(\u1/uk/K_r7_reg_n_0_[8] ),
        .O(\u1/u8/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__197_i_5
       (.I0(\u1/R7 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[36] ),
        .I3(\u1/uk/K_r7_reg_n_0_[29] ),
        .O(\u1/u8/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__197_i_6
       (.I0(\u1/R7 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[52] ),
        .I3(\u1/uk/K_r7_reg_n_0_[45] ),
        .O(\u1/u8/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__198
       (.I0(\u1/u8/X [5]),
        .I1(\u1/u8/X [4]),
        .I2(\u1/u8/X [3]),
        .I3(\u1/u8/X [2]),
        .I4(\u1/u8/X [6]),
        .I5(\u1/u8/X [1]),
        .O(\u1/out8 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__198_i_1
       (.I0(\u1/R7 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[54] ),
        .I3(\u1/uk/K_r7_reg_n_0_[47] ),
        .O(\u1/u8/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__198_i_2
       (.I0(\u1/R7 [3]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[19] ),
        .I3(\u1/uk/K_r7_reg_n_0_[12] ),
        .O(\u1/u8/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__198_i_3
       (.I0(\u1/R7 [2]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[10] ),
        .I3(\u1/uk/K_r7_reg_n_0_[3] ),
        .O(\u1/u8/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__198_i_4
       (.I0(\u1/R7 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[27] ),
        .I3(\u1/uk/K_r7_reg_n_0_[20] ),
        .O(\u1/u8/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__198_i_5
       (.I0(\u1/R7 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[25] ),
        .I3(\u1/uk/K_r7_reg_n_0_[18] ),
        .O(\u1/u8/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__198_i_6
       (.I0(\u1/R7 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r7_reg_n_0_[6] ),
        .I3(\u1/uk/K_r7_reg_n_0_[24] ),
        .O(\u1/u8/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__199
       (.I0(\u1/u9/X [41]),
        .I1(\u1/u9/X [40]),
        .I2(\u1/u9/X [39]),
        .I3(\u1/u9/X [38]),
        .I4(\u1/u9/X [42]),
        .I5(\u1/u9/X [37]),
        .O(\u1/out9 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__199_i_1
       (.I0(\u1/R8 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [44]),
        .I3(\u1/uk/K_r8 [9]),
        .O(\u1/u9/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__199_i_2
       (.I0(\u1/R8 [27]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [2]),
        .I3(\u1/uk/K_r8 [22]),
        .O(\u1/u9/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__199_i_3
       (.I0(\u1/R8 [26]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [52]),
        .I3(\u1/uk/K_r8 [44]),
        .O(\u1/u9/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__199_i_4
       (.I0(\u1/R8 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [8]),
        .I3(\u1/uk/K_r8 [28]),
        .O(\u1/u9/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__199_i_5
       (.I0(\u1/R8 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [36]),
        .I3(\u1/uk/K_r8 [1]),
        .O(\u1/u9/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__199_i_6
       (.I0(\u1/R8 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [28]),
        .I3(\u1/uk/K_r8 [52]),
        .O(\u1/u9/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__19_i_1
       (.I0(\u0/R1 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [28]),
        .I3(\u0/uk/K_r1 [38]),
        .O(\u0/u2/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__19_i_2
       (.I0(\u0/R1 [31]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [22]),
        .I3(\u0/uk/K_r1 [28]),
        .O(\u0/u2/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__19_i_3
       (.I0(\u0/R1 [30]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [38]),
        .I3(\u0/uk/K_r1 [16]),
        .O(\u0/u2/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__19_i_4
       (.I0(\u0/R1 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [9]),
        .I3(\u0/uk/K_r1 [15]),
        .O(\u0/u2/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__19_i_5
       (.I0(\u0/R1 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [49]),
        .I3(\u0/uk/K_r1 [0]),
        .O(\u0/u2/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__19_i_6
       (.I0(\u0/R1 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [37]),
        .I3(\u0/uk/K_r1 [43]),
        .O(\u0/u2/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__1_i_1
       (.I0(\u0/IP [56]),
        .I1(decrypt),
        .I2(\u0/key_r [35]),
        .I3(\u0/key_r [28]),
        .O(\u0/u0/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__1_i_2
       (.I0(\u0/IP [55]),
        .I1(decrypt),
        .I2(\u0/key_r [9]),
        .I3(\u0/key_r [2]),
        .O(\u0/u0/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__1_i_3
       (.I0(\u0/IP [54]),
        .I1(decrypt),
        .I2(\u0/key_r [51]),
        .I3(\u0/key_r [44]),
        .O(\u0/u0/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__1_i_4
       (.I0(\u0/IP [53]),
        .I1(decrypt),
        .I2(\u0/key_r [29]),
        .I3(\u0/key_r [22]),
        .O(\u0/u0/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__1_i_5
       (.I0(\u0/IP [57]),
        .I1(decrypt),
        .I2(\u0/key_r [30]),
        .I3(\u0/key_r [23]),
        .O(\u0/u0/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__1_i_6
       (.I0(\u0/IP [52]),
        .I1(decrypt),
        .I2(\u0/key_r [14]),
        .I3(\u0/key_r [7]),
        .O(\u0/u0/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__2
       (.I0(\u0/u0/X [11]),
        .I1(\u0/u0/X [10]),
        .I2(\u0/u0/X [9]),
        .I3(\u0/u0/X [8]),
        .I4(\u0/u0/X [12]),
        .I5(\u0/u0/X [7]),
        .O(\u0/out0 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__20
       (.I0(\u0/u2/X [23]),
        .I1(\u0/u2/X [22]),
        .I2(\u0/u2/X [21]),
        .I3(\u0/u2/X [20]),
        .I4(\u0/u2/X [24]),
        .I5(\u0/u2/X [19]),
        .O(\u0/out2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__200
       (.I0(\u1/u9/X [17]),
        .I1(\u1/u9/X [16]),
        .I2(\u1/u9/X [15]),
        .I3(\u1/u9/X [14]),
        .I4(\u1/u9/X [18]),
        .I5(\u1/u9/X [13]),
        .O(\u1/out9 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__200_i_1
       (.I0(\u1/R8 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [47]),
        .I3(\u1/uk/K_r8 [12]),
        .O(\u1/u9/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__200_i_2
       (.I0(\u1/R8 [11]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [32]),
        .I3(\u1/uk/K_r8 [54]),
        .O(\u1/u9/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__200_i_3
       (.I0(\u1/R8 [10]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [6]),
        .I3(\u1/uk/K_r8 [53]),
        .O(\u1/u9/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__200_i_4
       (.I0(\u1/R8 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [55]),
        .I3(\u1/uk/K_r8 [20]),
        .O(\u1/u9/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__200_i_5
       (.I0(\u1/R8 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [3]),
        .I3(\u1/uk/K_r8 [25]),
        .O(\u1/u9/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__200_i_6
       (.I0(\u1/R8 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [26]),
        .I3(\u1/uk/K_r8 [48]),
        .O(\u1/u9/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__201
       (.I0(\u1/u9/X [35]),
        .I1(\u1/u9/X [34]),
        .I2(\u1/u9/X [33]),
        .I3(\u1/u9/X [32]),
        .I4(\u1/u9/X [36]),
        .I5(\u1/u9/X [31]),
        .O(\u1/out9 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__201_i_1
       (.I0(\u1/R8 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [37]),
        .I3(\u1/uk/K_r8 [2]),
        .O(\u1/u9/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__201_i_2
       (.I0(\u1/R8 [23]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [35]),
        .I3(\u1/uk/K_r8 [0]),
        .O(\u1/u9/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__201_i_3
       (.I0(\u1/R8 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [22]),
        .I3(\u1/uk/K_r8 [42]),
        .O(\u1/u9/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__201_i_4
       (.I0(\u1/R8 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [0]),
        .I3(\u1/uk/K_r8 [51]),
        .O(\u1/u9/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__201_i_5
       (.I0(\u1/R8 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [1]),
        .I3(\u1/uk/K_r8 [21]),
        .O(\u1/u9/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__201_i_6
       (.I0(\u1/R8 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [16]),
        .I3(\u1/uk/K_r8 [36]),
        .O(\u1/u9/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__202
       (.I0(\u1/u9/X [11]),
        .I1(\u1/u9/X [10]),
        .I2(\u1/u9/X [9]),
        .I3(\u1/u9/X [8]),
        .I4(\u1/u9/X [12]),
        .I5(\u1/u9/X [7]),
        .O(\u1/out9 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__202_i_1
       (.I0(\u1/R8 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [12]),
        .I3(\u1/uk/K_r8 [34]),
        .O(\u1/u9/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__202_i_2
       (.I0(\u1/R8 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [46]),
        .I3(\u1/uk/K_r8 [11]),
        .O(\u1/u9/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__202_i_3
       (.I0(\u1/R8 [6]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [27]),
        .I3(\u1/uk/K_r8 [17]),
        .O(\u1/u9/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__202_i_4
       (.I0(\u1/R8 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [4]),
        .I3(\u1/uk/K_r8 [26]),
        .O(\u1/u9/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__202_i_5
       (.I0(\u1/R8 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [17]),
        .I3(\u1/uk/K_r8 [39]),
        .O(\u1/u9/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__202_i_6
       (.I0(\u1/R8 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [25]),
        .I3(\u1/uk/K_r8 [47]),
        .O(\u1/u9/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__203
       (.I0(\u1/u9/X [47]),
        .I1(\u1/u9/X [46]),
        .I2(\u1/u9/X [45]),
        .I3(\u1/u9/X [44]),
        .I4(\u1/u9/X [48]),
        .I5(\u1/u9/X [43]),
        .O(\u1/out9 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__203_i_1
       (.I0(\u1/R8 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [9]),
        .I3(\u1/uk/K_r8 [29]),
        .O(\u1/u9/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__203_i_2
       (.I0(\u1/R8 [31]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [31]),
        .I3(\u1/uk/K_r8 [23]),
        .O(\u1/u9/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__203_i_3
       (.I0(\u1/R8 [30]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [15]),
        .I3(\u1/uk/K_r8 [35]),
        .O(\u1/u9/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__203_i_4
       (.I0(\u1/R8 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [14]),
        .I3(\u1/uk/K_r8 [38]),
        .O(\u1/u9/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__203_i_5
       (.I0(\u1/R8 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [30]),
        .I3(\u1/uk/K_r8 [50]),
        .O(\u1/u9/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__203_i_6
       (.I0(\u1/R8 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [42]),
        .I3(\u1/uk/K_r8 [7]),
        .O(\u1/u9/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__204
       (.I0(\u1/u9/X [23]),
        .I1(\u1/u9/X [22]),
        .I2(\u1/u9/X [21]),
        .I3(\u1/u9/X [20]),
        .I4(\u1/u9/X [24]),
        .I5(\u1/u9/X [19]),
        .O(\u1/out9 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__204_i_1
       (.I0(\u1/R8 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [13]),
        .I3(\u1/uk/K_r8 [3]),
        .O(\u1/u9/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__204_i_2
       (.I0(\u1/R8 [15]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [5]),
        .I3(\u1/uk/K_r8 [27]),
        .O(\u1/u9/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__204_i_3
       (.I0(\u1/R8 [14]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [54]),
        .I3(\u1/uk/K_r8 [19]),
        .O(\u1/u9/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__204_i_4
       (.I0(\u1/R8 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [53]),
        .I3(\u1/uk/K_r8 [18]),
        .O(\u1/u9/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__204_i_5
       (.I0(\u1/R8 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [18]),
        .I3(\u1/uk/K_r8 [40]),
        .O(\u1/u9/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__204_i_6
       (.I0(\u1/R8 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [34]),
        .I3(\u1/uk/K_r8 [24]),
        .O(\u1/u9/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__205
       (.I0(\u1/u9/X [29]),
        .I1(\u1/u9/X [28]),
        .I2(\u1/u9/X [27]),
        .I3(\u1/u9/X [26]),
        .I4(\u1/u9/X [30]),
        .I5(\u1/u9/X [25]),
        .O(\u1/out9 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__205_i_1
       (.I0(\u1/R8 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [49]),
        .I3(\u1/uk/K_r8 [14]),
        .O(\u1/u9/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__205_i_2
       (.I0(\u1/R8 [19]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [38]),
        .I3(\u1/uk/K_r8 [30]),
        .O(\u1/u9/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__205_i_3
       (.I0(\u1/R8 [18]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [23]),
        .I3(\u1/uk/K_r8 [43]),
        .O(\u1/u9/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__205_i_4
       (.I0(\u1/R8 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [29]),
        .I3(\u1/uk/K_r8 [49]),
        .O(\u1/u9/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__205_i_5
       (.I0(\u1/R8 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [50]),
        .I3(\u1/uk/K_r8 [15]),
        .O(\u1/u9/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__205_i_6
       (.I0(\u1/R8 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [7]),
        .I3(\u1/uk/K_r8 [31]),
        .O(\u1/u9/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__206
       (.I0(\u1/u9/X [5]),
        .I1(\u1/u9/X [4]),
        .I2(\u1/u9/X [3]),
        .I3(\u1/u9/X [2]),
        .I4(\u1/u9/X [6]),
        .I5(\u1/u9/X [1]),
        .O(\u1/out9 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__206_i_1
       (.I0(\u1/R8 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [11]),
        .I3(\u1/uk/K_r8 [33]),
        .O(\u1/u9/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__206_i_2
       (.I0(\u1/R8 [3]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [33]),
        .I3(\u1/uk/K_r8 [55]),
        .O(\u1/u9/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__206_i_3
       (.I0(\u1/R8 [2]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [24]),
        .I3(\u1/uk/K_r8 [46]),
        .O(\u1/u9/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__206_i_4
       (.I0(\u1/R8 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [41]),
        .I3(\u1/uk/K_r8 [6]),
        .O(\u1/u9/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__206_i_5
       (.I0(\u1/R8 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [39]),
        .I3(\u1/uk/K_r8 [4]),
        .O(\u1/u9/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__206_i_6
       (.I0(\u1/R8 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r8 [20]),
        .I3(\u1/uk/K_r8 [10]),
        .O(\u1/u9/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__207
       (.I0(\u1/u10/X [41]),
        .I1(\u1/u10/X [40]),
        .I2(\u1/u10/X [39]),
        .I3(\u1/u10/X [38]),
        .I4(\u1/u10/X [42]),
        .I5(\u1/u10/X [37]),
        .O(\u1/out10 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__207_i_1
       (.I0(\u1/R9 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [31]),
        .I3(\u1/uk/K_r9 [50]),
        .O(\u1/u10/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__207_i_2
       (.I0(\u1/R9 [27]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [16]),
        .I3(\u1/uk/K_r9 [8]),
        .O(\u1/u10/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__207_i_3
       (.I0(\u1/R9 [26]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [7]),
        .I3(\u1/uk/K_r9 [30]),
        .O(\u1/u10/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__207_i_4
       (.I0(\u1/R9 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [22]),
        .I3(\u1/uk/K_r9 [14]),
        .O(\u1/u10/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__207_i_5
       (.I0(\u1/R9 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [50]),
        .I3(\u1/uk/K_r9 [42]),
        .O(\u1/u10/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__207_i_6
       (.I0(\u1/R9 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [42]),
        .I3(\u1/uk/K_r9 [38]),
        .O(\u1/u10/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__208
       (.I0(\u1/u10/X [17]),
        .I1(\u1/u10/X [16]),
        .I2(\u1/u10/X [15]),
        .I3(\u1/u10/X [14]),
        .I4(\u1/u10/X [18]),
        .I5(\u1/u10/X [13]),
        .O(\u1/out10 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__208_i_1
       (.I0(\u1/R9 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [4]),
        .I3(\u1/uk/K_r9 [55]),
        .O(\u1/u10/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__208_i_2
       (.I0(\u1/R9 [11]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [46]),
        .I3(\u1/uk/K_r9 [40]),
        .O(\u1/u10/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__208_i_3
       (.I0(\u1/R9 [10]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [20]),
        .I3(\u1/uk/K_r9 [39]),
        .O(\u1/u10/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__208_i_4
       (.I0(\u1/R9 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [12]),
        .I3(\u1/uk/K_r9 [6]),
        .O(\u1/u10/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__208_i_5
       (.I0(\u1/R9 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [17]),
        .I3(\u1/uk/K_r9 [11]),
        .O(\u1/u10/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__208_i_6
       (.I0(\u1/R9 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [40]),
        .I3(\u1/uk/K_r9 [34]),
        .O(\u1/u10/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__209
       (.I0(\u1/u10/X [35]),
        .I1(\u1/u10/X [34]),
        .I2(\u1/u10/X [33]),
        .I3(\u1/u10/X [32]),
        .I4(\u1/u10/X [36]),
        .I5(\u1/u10/X [31]),
        .O(\u1/out10 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__209_i_1
       (.I0(\u1/R9 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [51]),
        .I3(\u1/uk/K_r9 [43]),
        .O(\u1/u10/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__209_i_2
       (.I0(\u1/R9 [23]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [49]),
        .I3(\u1/uk/K_r9 [45]),
        .O(\u1/u10/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__209_i_3
       (.I0(\u1/R9 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [36]),
        .I3(\u1/uk/K_r9 [28]),
        .O(\u1/u10/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__209_i_4
       (.I0(\u1/R9 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [14]),
        .I3(\u1/uk/K_r9 [37]),
        .O(\u1/u10/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__209_i_5
       (.I0(\u1/R9 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [15]),
        .I3(\u1/uk/K_r9 [7]),
        .O(\u1/u10/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__209_i_6
       (.I0(\u1/R9 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [30]),
        .I3(\u1/uk/K_r9 [22]),
        .O(\u1/u10/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__20_i_1
       (.I0(\u0/R1 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [4]),
        .I3(\u0/uk/K_r1 [12]),
        .O(\u0/u2/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__20_i_2
       (.I0(\u0/R1 [15]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [53]),
        .I3(\u0/uk/K_r1 [4]),
        .O(\u0/u2/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__20_i_3
       (.I0(\u0/R1 [14]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [20]),
        .I3(\u0/uk/K_r1 [53]),
        .O(\u0/u2/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__20_i_4
       (.I0(\u0/R1 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [19]),
        .I3(\u0/uk/K_r1 [27]),
        .O(\u0/u2/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__20_i_5
       (.I0(\u0/R1 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [41]),
        .I3(\u0/uk/K_r1 [17]),
        .O(\u0/u2/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__20_i_6
       (.I0(\u0/R1 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [25]),
        .I3(\u0/uk/K_r1 [33]),
        .O(\u0/u2/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__21
       (.I0(\u0/u2/X [29]),
        .I1(\u0/u2/X [28]),
        .I2(\u0/u2/X [27]),
        .I3(\u0/u2/X [26]),
        .I4(\u0/u2/X [30]),
        .I5(\u0/u2/X [25]),
        .O(\u0/out2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__210
       (.I0(\u1/u10/X [11]),
        .I1(\u1/u10/X [10]),
        .I2(\u1/u10/X [9]),
        .I3(\u1/u10/X [8]),
        .I4(\u1/u10/X [12]),
        .I5(\u1/u10/X [7]),
        .O(\u1/out10 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__210_i_1
       (.I0(\u1/R9 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [26]),
        .I3(\u1/uk/K_r9 [20]),
        .O(\u1/u10/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__210_i_2
       (.I0(\u1/R9 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [3]),
        .I3(\u1/uk/K_r9 [54]),
        .O(\u1/u10/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__210_i_3
       (.I0(\u1/R9 [6]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [41]),
        .I3(\u1/uk/K_r9 [3]),
        .O(\u1/u10/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__210_i_4
       (.I0(\u1/R9 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [18]),
        .I3(\u1/uk/K_r9 [12]),
        .O(\u1/u10/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__210_i_5
       (.I0(\u1/R9 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [6]),
        .I3(\u1/uk/K_r9 [25]),
        .O(\u1/u10/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__210_i_6
       (.I0(\u1/R9 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [39]),
        .I3(\u1/uk/K_r9 [33]),
        .O(\u1/u10/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__211
       (.I0(\u1/u10/X [47]),
        .I1(\u1/u10/X [46]),
        .I2(\u1/u10/X [45]),
        .I3(\u1/u10/X [44]),
        .I4(\u1/u10/X [48]),
        .I5(\u1/u10/X [43]),
        .O(\u1/out10 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__211_i_1
       (.I0(\u1/R9 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [23]),
        .I3(\u1/uk/K_r9 [15]),
        .O(\u1/u10/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__211_i_2
       (.I0(\u1/R9 [31]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [45]),
        .I3(\u1/uk/K_r9 [9]),
        .O(\u1/u10/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__211_i_3
       (.I0(\u1/R9 [30]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [29]),
        .I3(\u1/uk/K_r9 [21]),
        .O(\u1/u10/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__211_i_4
       (.I0(\u1/R9 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [28]),
        .I3(\u1/uk/K_r9 [51]),
        .O(\u1/u10/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__211_i_5
       (.I0(\u1/R9 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [44]),
        .I3(\u1/uk/K_r9 [36]),
        .O(\u1/u10/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__211_i_6
       (.I0(\u1/R9 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [1]),
        .I3(\u1/uk/K_r9 [52]),
        .O(\u1/u10/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__212
       (.I0(\u1/u10/X [23]),
        .I1(\u1/u10/X [22]),
        .I2(\u1/u10/X [21]),
        .I3(\u1/u10/X [20]),
        .I4(\u1/u10/X [24]),
        .I5(\u1/u10/X [19]),
        .O(\u1/out10 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__212_i_1
       (.I0(\u1/R9 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [27]),
        .I3(\u1/uk/K_r9 [46]),
        .O(\u1/u10/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__212_i_2
       (.I0(\u1/R9 [15]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [19]),
        .I3(\u1/uk/K_r9 [13]),
        .O(\u1/u10/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__212_i_3
       (.I0(\u1/R9 [14]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [11]),
        .I3(\u1/uk/K_r9 [5]),
        .O(\u1/u10/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__212_i_4
       (.I0(\u1/R9 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [10]),
        .I3(\u1/uk/K_r9 [4]),
        .O(\u1/u10/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__212_i_5
       (.I0(\u1/R9 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [32]),
        .I3(\u1/uk/K_r9 [26]),
        .O(\u1/u10/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__212_i_6
       (.I0(\u1/R9 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [48]),
        .I3(\u1/uk/K_r9 [10]),
        .O(\u1/u10/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__213
       (.I0(\u1/u10/X [29]),
        .I1(\u1/u10/X [28]),
        .I2(\u1/u10/X [27]),
        .I3(\u1/u10/X [26]),
        .I4(\u1/u10/X [30]),
        .I5(\u1/u10/X [25]),
        .O(\u1/out10 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__213_i_1
       (.I0(\u1/R9 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [8]),
        .I3(\u1/uk/K_r9 [0]),
        .O(\u1/u10/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__213_i_2
       (.I0(\u1/R9 [19]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [52]),
        .I3(\u1/uk/K_r9 [16]),
        .O(\u1/u10/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__213_i_3
       (.I0(\u1/R9 [18]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [37]),
        .I3(\u1/uk/K_r9 [29]),
        .O(\u1/u10/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__213_i_4
       (.I0(\u1/R9 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [43]),
        .I3(\u1/uk/K_r9 [35]),
        .O(\u1/u10/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__213_i_5
       (.I0(\u1/R9 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [9]),
        .I3(\u1/uk/K_r9 [1]),
        .O(\u1/u10/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__213_i_6
       (.I0(\u1/R9 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [21]),
        .I3(\u1/uk/K_r9 [44]),
        .O(\u1/u10/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__214
       (.I0(\u1/u10/X [5]),
        .I1(\u1/u10/X [4]),
        .I2(\u1/u10/X [3]),
        .I3(\u1/u10/X [2]),
        .I4(\u1/u10/X [6]),
        .I5(\u1/u10/X [1]),
        .O(\u1/out10 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__214_i_1
       (.I0(\u1/R9 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [25]),
        .I3(\u1/uk/K_r9 [19]),
        .O(\u1/u10/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__214_i_2
       (.I0(\u1/R9 [3]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [47]),
        .I3(\u1/uk/K_r9 [41]),
        .O(\u1/u10/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__214_i_3
       (.I0(\u1/R9 [2]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [13]),
        .I3(\u1/uk/K_r9 [32]),
        .O(\u1/u10/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__214_i_4
       (.I0(\u1/R9 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [55]),
        .I3(\u1/uk/K_r9 [17]),
        .O(\u1/u10/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__214_i_5
       (.I0(\u1/R9 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [53]),
        .I3(\u1/uk/K_r9 [47]),
        .O(\u1/u10/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__214_i_6
       (.I0(\u1/R9 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r9 [34]),
        .I3(\u1/uk/K_r9 [53]),
        .O(\u1/u10/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__215
       (.I0(\u1/u11/X [41]),
        .I1(\u1/u11/X [40]),
        .I2(\u1/u11/X [39]),
        .I3(\u1/u11/X [38]),
        .I4(\u1/u11/X [42]),
        .I5(\u1/u11/X [37]),
        .O(\u1/out11 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__215_i_1
       (.I0(\u1/R10_reg_n_0_[28] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [45]),
        .I3(\u1/uk/K_r10 [36]),
        .O(\u1/u11/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__215_i_2
       (.I0(\u1/R10_reg_n_0_[27] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [30]),
        .I3(\u1/uk/K_r10 [49]),
        .O(\u1/u11/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__215_i_3
       (.I0(\u1/R10_reg_n_0_[26] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [21]),
        .I3(\u1/uk/K_r10 [16]),
        .O(\u1/u11/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__215_i_4
       (.I0(\u1/R10_reg_n_0_[25] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [36]),
        .I3(\u1/uk/K_r10 [0]),
        .O(\u1/u11/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__215_i_5
       (.I0(\u1/R10_reg_n_0_[29] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [9]),
        .I3(\u1/uk/K_r10 [28]),
        .O(\u1/u11/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__215_i_6
       (.I0(\u1/R10_reg_n_0_[24] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [1]),
        .I3(\u1/uk/K_r10 [51]),
        .O(\u1/u11/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__216
       (.I0(\u1/u11/X [17]),
        .I1(\u1/u11/X [16]),
        .I2(\u1/u11/X [15]),
        .I3(\u1/u11/X [14]),
        .I4(\u1/u11/X [18]),
        .I5(\u1/u11/X [13]),
        .O(\u1/out11 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__216_i_1
       (.I0(\u1/R10_reg_n_0_[12] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [18]),
        .I3(\u1/uk/K_r10 [41]),
        .O(\u1/u11/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__216_i_2
       (.I0(\u1/R10_reg_n_0_[11] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [3]),
        .I3(\u1/uk/K_r10 [26]),
        .O(\u1/u11/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__216_i_3
       (.I0(\u1/R10_reg_n_0_ ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [34]),
        .I3(\u1/uk/K_r10 [25]),
        .O(\u1/u11/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__216_i_4
       (.I0(\u1/R10_reg_n_0_[9] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [26]),
        .I3(\u1/uk/K_r10 [17]),
        .O(\u1/u11/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__216_i_5
       (.I0(\u1/R10_reg_n_0_[13] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [6]),
        .I3(\u1/uk/K_r10 [54]),
        .O(\u1/u11/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__216_i_6
       (.I0(\u1/R10_reg_n_0_[8] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [54]),
        .I3(\u1/uk/K_r10 [20]),
        .O(\u1/u11/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__217
       (.I0(\u1/u11/X [35]),
        .I1(\u1/u11/X [34]),
        .I2(\u1/u11/X [33]),
        .I3(\u1/u11/X [32]),
        .I4(\u1/u11/X [36]),
        .I5(\u1/u11/X [31]),
        .O(\u1/out11 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__217_i_1
       (.I0(\u1/R10_reg_n_0_[24] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [38]),
        .I3(\u1/uk/K_r10 [29]),
        .O(\u1/u11/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__217_i_2
       (.I0(\u1/R10_reg_n_0_[23] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [8]),
        .I3(\u1/uk/K_r10 [31]),
        .O(\u1/u11/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__217_i_3
       (.I0(\u1/R10_reg_n_0_[22] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [50]),
        .I3(\u1/uk/K_r10 [14]),
        .O(\u1/u11/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__217_i_4
       (.I0(\u1/R10_reg_n_0_[21] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [28]),
        .I3(\u1/uk/K_r10 [23]),
        .O(\u1/u11/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__217_i_5
       (.I0(\u1/R10_reg_n_0_[25] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [29]),
        .I3(\u1/uk/K_r10 [52]),
        .O(\u1/u11/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__217_i_6
       (.I0(\u1/R10_reg_n_0_[20] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [44]),
        .I3(\u1/uk/K_r10 [8]),
        .O(\u1/u11/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__218
       (.I0(\u1/u11/X [11]),
        .I1(\u1/u11/X [10]),
        .I2(\u1/u11/X [9]),
        .I3(\u1/u11/X [8]),
        .I4(\u1/u11/X [12]),
        .I5(\u1/u11/X [7]),
        .O(\u1/out11 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__218_i_1
       (.I0(\u1/R10_reg_n_0_[8] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [40]),
        .I3(\u1/uk/K_r10 [6]),
        .O(\u1/u11/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__218_i_2
       (.I0(\u1/R10_reg_n_0_[7] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [17]),
        .I3(\u1/uk/K_r10 [40]),
        .O(\u1/u11/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__218_i_3
       (.I0(\u1/R10_reg_n_0_[6] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [55]),
        .I3(\u1/uk/K_r10 [46]),
        .O(\u1/u11/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__218_i_4
       (.I0(\u1/R10_reg_n_0_[5] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [32]),
        .I3(\u1/uk/K_r10 [55]),
        .O(\u1/u11/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__218_i_5
       (.I0(\u1/R10_reg_n_0_[9] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [20]),
        .I3(\u1/uk/K_r10 [11]),
        .O(\u1/u11/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__218_i_6
       (.I0(\u1/R10_reg_n_0_[4] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [53]),
        .I3(\u1/uk/K_r10 [19]),
        .O(\u1/u11/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__219
       (.I0(\u1/u11/X [47]),
        .I1(\u1/u11/X [46]),
        .I2(\u1/u11/X [45]),
        .I3(\u1/u11/X [44]),
        .I4(\u1/u11/X [48]),
        .I5(\u1/u11/X [43]),
        .O(\u1/out11 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__219_i_1
       (.I0(\u1/R10_reg_n_0_[32] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [37]),
        .I3(\u1/uk/K_r10 [1]),
        .O(\u1/u11/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__219_i_2
       (.I0(\u1/R10_reg_n_0_[31] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [0]),
        .I3(\u1/uk/K_r10 [50]),
        .O(\u1/u11/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__219_i_3
       (.I0(\u1/R10_reg_n_0_[30] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [43]),
        .I3(\u1/uk/K_r10 [7]),
        .O(\u1/u11/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__219_i_4
       (.I0(\u1/R10_reg_n_0_[29] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [42]),
        .I3(\u1/uk/K_r10 [37]),
        .O(\u1/u11/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__219_i_5
       (.I0(\u1/R10_reg_n_0_[1] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [31]),
        .I3(\u1/uk/K_r10 [22]),
        .O(\u1/u11/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__219_i_6
       (.I0(\u1/R10_reg_n_0_[28] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [15]),
        .I3(\u1/uk/K_r10 [38]),
        .O(\u1/u11/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__21_i_1
       (.I0(\u0/R1 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [44]),
        .I3(\u0/uk/K_r1 [50]),
        .O(\u0/u2/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__21_i_2
       (.I0(\u0/R1 [19]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [29]),
        .I3(\u0/uk/K_r1 [35]),
        .O(\u0/u2/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__21_i_3
       (.I0(\u0/R1 [18]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [42]),
        .I3(\u0/uk/K_r1 [52]),
        .O(\u0/u2/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__21_i_4
       (.I0(\u0/R1 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [52]),
        .I3(\u0/uk/K_r1 [30]),
        .O(\u0/u2/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__21_i_5
       (.I0(\u0/R1 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [14]),
        .I3(\u0/uk/K_r1 [51]),
        .O(\u0/u2/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__21_i_6
       (.I0(\u0/R1 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [2]),
        .I3(\u0/uk/K_r1 [8]),
        .O(\u0/u2/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__22
       (.I0(\u0/u2/X [5]),
        .I1(\u0/u2/X [4]),
        .I2(\u0/u2/X [3]),
        .I3(\u0/u2/X [2]),
        .I4(\u0/u2/X [6]),
        .I5(\u0/u2/X [1]),
        .O(\u0/out2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__220
       (.I0(\u1/u11/X [23]),
        .I1(\u1/u11/X [22]),
        .I2(\u1/u11/X [21]),
        .I3(\u1/u11/X [20]),
        .I4(\u1/u11/X [24]),
        .I5(\u1/u11/X [19]),
        .O(\u1/out11 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__220_i_1
       (.I0(\u1/R10_reg_n_0_[16] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [41]),
        .I3(\u1/uk/K_r10 [32]),
        .O(\u1/u11/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__220_i_2
       (.I0(\u1/R10_reg_n_0_[15] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [33]),
        .I3(\u1/uk/K_r10 [24]),
        .O(\u1/u11/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__220_i_3
       (.I0(\u1/R10_reg_n_0_[14] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [25]),
        .I3(\u1/uk/K_r10 [48]),
        .O(\u1/u11/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__220_i_4
       (.I0(\u1/R10_reg_n_0_[13] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [24]),
        .I3(\u1/uk/K_r10 [47]),
        .O(\u1/u11/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__220_i_5
       (.I0(\u1/R10_reg_n_0_[17] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [46]),
        .I3(\u1/uk/K_r10 [12]),
        .O(\u1/u11/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__220_i_6
       (.I0(\u1/R10_reg_n_0_[12] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [5]),
        .I3(\u1/uk/K_r10 [53]),
        .O(\u1/u11/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__221
       (.I0(\u1/u11/X [29]),
        .I1(\u1/u11/X [28]),
        .I2(\u1/u11/X [27]),
        .I3(\u1/u11/X [26]),
        .I4(\u1/u11/X [30]),
        .I5(\u1/u11/X [25]),
        .O(\u1/out11 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__221_i_1
       (.I0(\u1/R10_reg_n_0_[20] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [22]),
        .I3(\u1/uk/K_r10 [45]),
        .O(\u1/u11/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__221_i_2
       (.I0(\u1/R10_reg_n_0_[19] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [7]),
        .I3(\u1/uk/K_r10 [2]),
        .O(\u1/u11/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__221_i_3
       (.I0(\u1/R10_reg_n_0_[18] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [51]),
        .I3(\u1/uk/K_r10 [15]),
        .O(\u1/u11/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__221_i_4
       (.I0(\u1/R10_reg_n_0_[17] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [2]),
        .I3(\u1/uk/K_r10 [21]),
        .O(\u1/u11/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__221_i_5
       (.I0(\u1/R10_reg_n_0_[21] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [23]),
        .I3(\u1/uk/K_r10 [42]),
        .O(\u1/u11/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__221_i_6
       (.I0(\u1/R10_reg_n_0_[16] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [35]),
        .I3(\u1/uk/K_r10 [30]),
        .O(\u1/u11/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__222
       (.I0(\u1/u11/X [5]),
        .I1(\u1/u11/X [4]),
        .I2(\u1/u11/X [3]),
        .I3(\u1/u11/X [2]),
        .I4(\u1/u11/X [6]),
        .I5(\u1/u11/X [1]),
        .O(\u1/out11 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__222_i_1
       (.I0(\u1/R10_reg_n_0_[4] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [39]),
        .I3(\u1/uk/K_r10 [5]),
        .O(\u1/u11/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__222_i_2
       (.I0(\u1/R10_reg_n_0_[3] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [4]),
        .I3(\u1/uk/K_r10 [27]),
        .O(\u1/u11/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__222_i_3
       (.I0(\u1/R10_reg_n_0_[2] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [27]),
        .I3(\u1/uk/K_r10 [18]),
        .O(\u1/u11/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__222_i_4
       (.I0(\u1/R10_reg_n_0_[1] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [12]),
        .I3(\u1/uk/K_r10 [3]),
        .O(\u1/u11/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__222_i_5
       (.I0(\u1/R10_reg_n_0_[5] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [10]),
        .I3(\u1/uk/K_r10 [33]),
        .O(\u1/u11/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__222_i_6
       (.I0(\u1/R10_reg_n_0_[32] ),
        .I1(decrypt),
        .I2(\u1/uk/K_r10 [48]),
        .I3(\u1/uk/K_r10 [39]),
        .O(\u1/u11/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__223
       (.I0(\u1/u12/X [41]),
        .I1(\u1/u12/X [40]),
        .I2(\u1/u12/X [39]),
        .I3(\u1/u12/X [38]),
        .I4(\u1/u12/X [42]),
        .I5(\u1/u12/X [37]),
        .O(\u1/out12 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__223_i_1
       (.I0(\u1/R11 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [0]),
        .I3(\u1/uk/K_r11 [22]),
        .O(\u1/u12/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__223_i_2
       (.I0(\u1/R11 [27]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [44]),
        .I3(\u1/uk/K_r11 [35]),
        .O(\u1/u12/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__223_i_3
       (.I0(\u1/R11 [26]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [35]),
        .I3(\u1/uk/K_r11 [2]),
        .O(\u1/u12/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__223_i_4
       (.I0(\u1/R11 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [50]),
        .I3(\u1/uk/K_r11 [45]),
        .O(\u1/u12/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__223_i_5
       (.I0(\u1/R11 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [23]),
        .I3(\u1/uk/K_r11 [14]),
        .O(\u1/u12/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__223_i_6
       (.I0(\u1/R11 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [15]),
        .I3(\u1/uk/K_r11 [37]),
        .O(\u1/u12/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__224
       (.I0(\u1/u12/X [17]),
        .I1(\u1/u12/X [16]),
        .I2(\u1/u12/X [15]),
        .I3(\u1/u12/X [14]),
        .I4(\u1/u12/X [18]),
        .I5(\u1/u12/X [13]),
        .O(\u1/out12 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__224_i_1
       (.I0(\u1/R11 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [32]),
        .I3(\u1/uk/K_r11 [27]),
        .O(\u1/u12/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__224_i_2
       (.I0(\u1/R11 [11]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [17]),
        .I3(\u1/uk/K_r11 [12]),
        .O(\u1/u12/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__224_i_3
       (.I0(\u1/R11 [10]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [48]),
        .I3(\u1/uk/K_r11 [11]),
        .O(\u1/u12/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__224_i_4
       (.I0(\u1/R11 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [40]),
        .I3(\u1/uk/K_r11 [3]),
        .O(\u1/u12/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__224_i_5
       (.I0(\u1/R11 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [20]),
        .I3(\u1/uk/K_r11 [40]),
        .O(\u1/u12/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__224_i_6
       (.I0(\u1/R11 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [11]),
        .I3(\u1/uk/K_r11 [6]),
        .O(\u1/u12/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__225
       (.I0(\u1/u12/X [35]),
        .I1(\u1/u12/X [34]),
        .I2(\u1/u12/X [33]),
        .I3(\u1/u12/X [32]),
        .I4(\u1/u12/X [36]),
        .I5(\u1/u12/X [31]),
        .O(\u1/out12 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__225_i_1
       (.I0(\u1/R11 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [52]),
        .I3(\u1/uk/K_r11 [15]),
        .O(\u1/u12/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__225_i_2
       (.I0(\u1/R11 [23]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [22]),
        .I3(\u1/uk/K_r11 [44]),
        .O(\u1/u12/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__225_i_3
       (.I0(\u1/R11 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [9]),
        .I3(\u1/uk/K_r11 [0]),
        .O(\u1/u12/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__225_i_4
       (.I0(\u1/R11 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [42]),
        .I3(\u1/uk/K_r11 [9]),
        .O(\u1/u12/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__225_i_5
       (.I0(\u1/R11 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [43]),
        .I3(\u1/uk/K_r11 [38]),
        .O(\u1/u12/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__225_i_6
       (.I0(\u1/R11 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [31]),
        .I3(\u1/uk/K_r11 [49]),
        .O(\u1/u12/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__226
       (.I0(\u1/u12/X [11]),
        .I1(\u1/u12/X [10]),
        .I2(\u1/u12/X [9]),
        .I3(\u1/u12/X [8]),
        .I4(\u1/u12/X [12]),
        .I5(\u1/u12/X [7]),
        .O(\u1/out12 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__226_i_1
       (.I0(\u1/R11 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [54]),
        .I3(\u1/uk/K_r11 [17]),
        .O(\u1/u12/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__226_i_2
       (.I0(\u1/R11 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [6]),
        .I3(\u1/uk/K_r11 [26]),
        .O(\u1/u12/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__226_i_3
       (.I0(\u1/R11 [6]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [12]),
        .I3(\u1/uk/K_r11 [32]),
        .O(\u1/u12/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__226_i_4
       (.I0(\u1/R11 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [46]),
        .I3(\u1/uk/K_r11 [41]),
        .O(\u1/u12/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__226_i_5
       (.I0(\u1/R11 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [34]),
        .I3(\u1/uk/K_r11 [54]),
        .O(\u1/u12/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__226_i_6
       (.I0(\u1/R11 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [10]),
        .I3(\u1/uk/K_r11 [5]),
        .O(\u1/u12/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__227
       (.I0(\u1/u12/X [47]),
        .I1(\u1/u12/X [46]),
        .I2(\u1/u12/X [45]),
        .I3(\u1/u12/X [44]),
        .I4(\u1/u12/X [48]),
        .I5(\u1/u12/X [43]),
        .O(\u1/out12 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__227_i_1
       (.I0(\u1/R11 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [51]),
        .I3(\u1/uk/K_r11 [42]),
        .O(\u1/u12/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__227_i_2
       (.I0(\u1/R11 [31]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [14]),
        .I3(\u1/uk/K_r11 [36]),
        .O(\u1/u12/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__227_i_3
       (.I0(\u1/R11 [30]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [2]),
        .I3(\u1/uk/K_r11 [52]),
        .O(\u1/u12/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__227_i_4
       (.I0(\u1/R11 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [1]),
        .I3(\u1/uk/K_r11 [23]),
        .O(\u1/u12/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__227_i_5
       (.I0(\u1/R11 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [45]),
        .I3(\u1/uk/K_r11 [8]),
        .O(\u1/u12/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__227_i_6
       (.I0(\u1/R11 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [29]),
        .I3(\u1/uk/K_r11 [51]),
        .O(\u1/u12/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__228
       (.I0(\u1/u12/X [23]),
        .I1(\u1/u12/X [22]),
        .I2(\u1/u12/X [21]),
        .I3(\u1/u12/X [20]),
        .I4(\u1/u12/X [24]),
        .I5(\u1/u12/X [19]),
        .O(\u1/out12 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__228_i_1
       (.I0(\u1/R11 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [55]),
        .I3(\u1/uk/K_r11 [18]),
        .O(\u1/u12/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__228_i_2
       (.I0(\u1/R11 [15]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [47]),
        .I3(\u1/uk/K_r11 [10]),
        .O(\u1/u12/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__228_i_3
       (.I0(\u1/R11 [14]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [39]),
        .I3(\u1/uk/K_r11 [34]),
        .O(\u1/u12/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__228_i_4
       (.I0(\u1/R11 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [13]),
        .I3(\u1/uk/K_r11 [33]),
        .O(\u1/u12/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__228_i_5
       (.I0(\u1/R11 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [3]),
        .I3(\u1/uk/K_r11 [55]),
        .O(\u1/u12/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__228_i_6
       (.I0(\u1/R11 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [19]),
        .I3(\u1/uk/K_r11 [39]),
        .O(\u1/u12/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__229
       (.I0(\u1/u12/X [29]),
        .I1(\u1/u12/X [28]),
        .I2(\u1/u12/X [27]),
        .I3(\u1/u12/X [26]),
        .I4(\u1/u12/X [30]),
        .I5(\u1/u12/X [25]),
        .O(\u1/out12 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__229_i_1
       (.I0(\u1/R11 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [36]),
        .I3(\u1/uk/K_r11 [31]),
        .O(\u1/u12/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__229_i_2
       (.I0(\u1/R11 [19]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [21]),
        .I3(\u1/uk/K_r11 [43]),
        .O(\u1/u12/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__229_i_3
       (.I0(\u1/R11 [18]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [38]),
        .I3(\u1/uk/K_r11 [1]),
        .O(\u1/u12/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__229_i_4
       (.I0(\u1/R11 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [16]),
        .I3(\u1/uk/K_r11 [7]),
        .O(\u1/u12/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__229_i_5
       (.I0(\u1/R11 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [37]),
        .I3(\u1/uk/K_r11 [28]),
        .O(\u1/u12/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__229_i_6
       (.I0(\u1/R11 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [49]),
        .I3(\u1/uk/K_r11 [16]),
        .O(\u1/u12/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__22_i_1
       (.I0(\u0/R1 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [34]),
        .I3(\u0/uk/K_r1 [10]),
        .O(\u0/u2/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__22_i_2
       (.I0(\u0/R1 [3]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [24]),
        .I3(\u0/uk/K_r1 [32]),
        .O(\u0/u2/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__22_i_3
       (.I0(\u0/R1 [2]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [47]),
        .I3(\u0/uk/K_r1 [55]),
        .O(\u0/u2/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__22_i_4
       (.I0(\u0/R1 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [32]),
        .I3(\u0/uk/K_r1 [40]),
        .O(\u0/u2/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__22_i_5
       (.I0(\u0/R1 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [5]),
        .I3(\u0/uk/K_r1 [13]),
        .O(\u0/u2/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__22_i_6
       (.I0(\u0/R1 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r1 [11]),
        .I3(\u0/uk/K_r1 [19]),
        .O(\u0/u2/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__23
       (.I0(\u0/u3/X [41]),
        .I1(\u0/u3/X [40]),
        .I2(\u0/u3/X [39]),
        .I3(\u0/u3/X [38]),
        .I4(\u0/u3/X [42]),
        .I5(\u0/u3/X [37]),
        .O(\u0/out3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__230
       (.I0(\u1/u12/X [5]),
        .I1(\u1/u12/X [4]),
        .I2(\u1/u12/X [3]),
        .I3(\u1/u12/X [2]),
        .I4(\u1/u12/X [6]),
        .I5(\u1/u12/X [1]),
        .O(\u1/out12 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__230_i_1
       (.I0(\u1/R11 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [53]),
        .I3(\u1/uk/K_r11 [48]),
        .O(\u1/u12/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__230_i_2
       (.I0(\u1/R11 [3]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [18]),
        .I3(\u1/uk/K_r11 [13]),
        .O(\u1/u12/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__230_i_3
       (.I0(\u1/R11 [2]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [41]),
        .I3(\u1/uk/K_r11 [4]),
        .O(\u1/u12/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__230_i_4
       (.I0(\u1/R11 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [26]),
        .I3(\u1/uk/K_r11 [46]),
        .O(\u1/u12/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__230_i_5
       (.I0(\u1/R11 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [24]),
        .I3(\u1/uk/K_r11 [19]),
        .O(\u1/u12/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__230_i_6
       (.I0(\u1/R11 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r11 [5]),
        .I3(\u1/uk/K_r11 [25]),
        .O(\u1/u12/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__231
       (.I0(\u1/u13/X [41]),
        .I1(\u1/u13/X [40]),
        .I2(\u1/u13/X [39]),
        .I3(\u1/u13/X [38]),
        .I4(\u1/u13/X [42]),
        .I5(\u1/u13/X [37]),
        .O(\u1/out13 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__231_i_1
       (.I0(\u1/R12 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [14]),
        .I3(\u1/uk/K_r12 [8]),
        .O(\u1/u13/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__231_i_2
       (.I0(\u1/R12 [27]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [31]),
        .I3(\u1/uk/K_r12 [21]),
        .O(\u1/u13/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__231_i_3
       (.I0(\u1/R12 [26]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [49]),
        .I3(\u1/uk/K_r12 [43]),
        .O(\u1/u13/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__231_i_4
       (.I0(\u1/R12 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [9]),
        .I3(\u1/uk/K_r12 [31]),
        .O(\u1/u13/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__231_i_5
       (.I0(\u1/R12 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [37]),
        .I3(\u1/uk/K_r12 [0]),
        .O(\u1/u13/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__231_i_6
       (.I0(\u1/R12 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [29]),
        .I3(\u1/uk/K_r12 [23]),
        .O(\u1/u13/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__232
       (.I0(\u1/u13/X [17]),
        .I1(\u1/u13/X [16]),
        .I2(\u1/u13/X [15]),
        .I3(\u1/u13/X [14]),
        .I4(\u1/u13/X [18]),
        .I5(\u1/u13/X [13]),
        .O(\u1/out13 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__232_i_1
       (.I0(\u1/R12 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [46]),
        .I3(\u1/uk/K_r12 [13]),
        .O(\u1/u13/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__232_i_2
       (.I0(\u1/R12 [11]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [6]),
        .I3(\u1/uk/K_r12 [55]),
        .O(\u1/u13/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__232_i_3
       (.I0(\u1/R12 [10]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [5]),
        .I3(\u1/uk/K_r12 [54]),
        .O(\u1/u13/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__232_i_4
       (.I0(\u1/R12 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [54]),
        .I3(\u1/uk/K_r12 [46]),
        .O(\u1/u13/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__232_i_5
       (.I0(\u1/R12 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [34]),
        .I3(\u1/uk/K_r12 [26]),
        .O(\u1/u13/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__232_i_6
       (.I0(\u1/R12 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [25]),
        .I3(\u1/uk/K_r12 [17]),
        .O(\u1/u13/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__233
       (.I0(\u1/u13/X [35]),
        .I1(\u1/u13/X [34]),
        .I2(\u1/u13/X [33]),
        .I3(\u1/u13/X [32]),
        .I4(\u1/u13/X [36]),
        .I5(\u1/u13/X [31]),
        .O(\u1/out13 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__233_i_1
       (.I0(\u1/R12 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [7]),
        .I3(\u1/uk/K_r12 [1]),
        .O(\u1/u13/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__233_i_2
       (.I0(\u1/R12 [23]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [36]),
        .I3(\u1/uk/K_r12 [30]),
        .O(\u1/u13/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__233_i_3
       (.I0(\u1/R12 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [23]),
        .I3(\u1/uk/K_r12 [45]),
        .O(\u1/u13/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__233_i_4
       (.I0(\u1/R12 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [1]),
        .I3(\u1/uk/K_r12 [50]),
        .O(\u1/u13/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__233_i_5
       (.I0(\u1/R12 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [2]),
        .I3(\u1/uk/K_r12 [51]),
        .O(\u1/u13/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__233_i_6
       (.I0(\u1/R12 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [45]),
        .I3(\u1/uk/K_r12 [35]),
        .O(\u1/u13/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__234
       (.I0(\u1/u13/X [11]),
        .I1(\u1/u13/X [10]),
        .I2(\u1/u13/X [9]),
        .I3(\u1/u13/X [8]),
        .I4(\u1/u13/X [12]),
        .I5(\u1/u13/X [7]),
        .O(\u1/out13 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__234_i_1
       (.I0(\u1/R12 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [11]),
        .I3(\u1/uk/K_r12 [3]),
        .O(\u1/u13/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__234_i_2
       (.I0(\u1/R12 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [20]),
        .I3(\u1/uk/K_r12 [12]),
        .O(\u1/u13/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__234_i_3
       (.I0(\u1/R12 [6]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [26]),
        .I3(\u1/uk/K_r12 [18]),
        .O(\u1/u13/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__234_i_4
       (.I0(\u1/R12 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [3]),
        .I3(\u1/uk/K_r12 [27]),
        .O(\u1/u13/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__234_i_5
       (.I0(\u1/R12 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [48]),
        .I3(\u1/uk/K_r12 [40]),
        .O(\u1/u13/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__234_i_6
       (.I0(\u1/R12 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [24]),
        .I3(\u1/uk/K_r12 [48]),
        .O(\u1/u13/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__235
       (.I0(\u1/u13/X [47]),
        .I1(\u1/u13/X [46]),
        .I2(\u1/u13/X [45]),
        .I3(\u1/u13/X [44]),
        .I4(\u1/u13/X [48]),
        .I5(\u1/u13/X [43]),
        .O(\u1/out13 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__235_i_1
       (.I0(\u1/R12 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [38]),
        .I3(\u1/uk/K_r12 [28]),
        .O(\u1/u13/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__235_i_2
       (.I0(\u1/R12 [31]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [28]),
        .I3(\u1/uk/K_r12 [22]),
        .O(\u1/u13/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__235_i_3
       (.I0(\u1/R12 [30]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [16]),
        .I3(\u1/uk/K_r12 [38]),
        .O(\u1/u13/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__235_i_4
       (.I0(\u1/R12 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [15]),
        .I3(\u1/uk/K_r12 [9]),
        .O(\u1/u13/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__235_i_5
       (.I0(\u1/R12 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [0]),
        .I3(\u1/uk/K_r12 [49]),
        .O(\u1/u13/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__235_i_6
       (.I0(\u1/R12 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [43]),
        .I3(\u1/uk/K_r12 [37]),
        .O(\u1/u13/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__236
       (.I0(\u1/u13/X [23]),
        .I1(\u1/u13/X [22]),
        .I2(\u1/u13/X [21]),
        .I3(\u1/u13/X [20]),
        .I4(\u1/u13/X [24]),
        .I5(\u1/u13/X [19]),
        .O(\u1/out13 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__236_i_1
       (.I0(\u1/R12 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [12]),
        .I3(\u1/uk/K_r12 [4]),
        .O(\u1/u13/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__236_i_2
       (.I0(\u1/R12 [15]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [4]),
        .I3(\u1/uk/K_r12 [53]),
        .O(\u1/u13/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__236_i_3
       (.I0(\u1/R12 [14]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [53]),
        .I3(\u1/uk/K_r12 [20]),
        .O(\u1/u13/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__236_i_4
       (.I0(\u1/R12 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [27]),
        .I3(\u1/uk/K_r12 [19]),
        .O(\u1/u13/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__236_i_5
       (.I0(\u1/R12 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [17]),
        .I3(\u1/uk/K_r12 [41]),
        .O(\u1/u13/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__236_i_6
       (.I0(\u1/R12 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [33]),
        .I3(\u1/uk/K_r12 [25]),
        .O(\u1/u13/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__237
       (.I0(\u1/u13/X [29]),
        .I1(\u1/u13/X [28]),
        .I2(\u1/u13/X [27]),
        .I3(\u1/u13/X [26]),
        .I4(\u1/u13/X [30]),
        .I5(\u1/u13/X [25]),
        .O(\u1/out13 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__237_i_1
       (.I0(\u1/R12 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [50]),
        .I3(\u1/uk/K_r12 [44]),
        .O(\u1/u13/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__237_i_2
       (.I0(\u1/R12 [19]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [35]),
        .I3(\u1/uk/K_r12 [29]),
        .O(\u1/u13/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__237_i_3
       (.I0(\u1/R12 [18]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [52]),
        .I3(\u1/uk/K_r12 [42]),
        .O(\u1/u13/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__237_i_4
       (.I0(\u1/R12 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [30]),
        .I3(\u1/uk/K_r12 [52]),
        .O(\u1/u13/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__237_i_5
       (.I0(\u1/R12 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [51]),
        .I3(\u1/uk/K_r12 [14]),
        .O(\u1/u13/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__237_i_6
       (.I0(\u1/R12 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [8]),
        .I3(\u1/uk/K_r12 [2]),
        .O(\u1/u13/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__238
       (.I0(\u1/u13/X [5]),
        .I1(\u1/u13/X [4]),
        .I2(\u1/u13/X [3]),
        .I3(\u1/u13/X [2]),
        .I4(\u1/u13/X [6]),
        .I5(\u1/u13/X [1]),
        .O(\u1/out13 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__238_i_1
       (.I0(\u1/R12 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [10]),
        .I3(\u1/uk/K_r12 [34]),
        .O(\u1/u13/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__238_i_2
       (.I0(\u1/R12 [3]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [32]),
        .I3(\u1/uk/K_r12 [24]),
        .O(\u1/u13/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__238_i_3
       (.I0(\u1/R12 [2]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [55]),
        .I3(\u1/uk/K_r12 [47]),
        .O(\u1/u13/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__238_i_4
       (.I0(\u1/R12 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [40]),
        .I3(\u1/uk/K_r12 [32]),
        .O(\u1/u13/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__238_i_5
       (.I0(\u1/R12 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [13]),
        .I3(\u1/uk/K_r12 [5]),
        .O(\u1/u13/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__238_i_6
       (.I0(\u1/R12 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r12 [19]),
        .I3(\u1/uk/K_r12 [11]),
        .O(\u1/u13/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__239
       (.I0(\u1/u14/X [41]),
        .I1(\u1/u14/X [40]),
        .I2(\u1/u14/X [39]),
        .I3(\u1/u14/X [38]),
        .I4(\u1/u14/X [42]),
        .I5(\u1/u14/X [37]),
        .O(\u1/out14 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__239_i_1
       (.I0(\u1/R13 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [28]),
        .I3(\u1/uk/K_r13 [49]),
        .O(\u1/u14/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__239_i_2
       (.I0(\u1/R13 [27]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [45]),
        .I3(\u1/uk/K_r13 [7]),
        .O(\u1/u14/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__239_i_3
       (.I0(\u1/R13 [26]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [8]),
        .I3(\u1/uk/K_r13 [29]),
        .O(\u1/u14/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__239_i_4
       (.I0(\u1/R13 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [23]),
        .I3(\u1/uk/K_r13 [44]),
        .O(\u1/u14/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__239_i_5
       (.I0(\u1/R13 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [51]),
        .I3(\u1/uk/K_r13 [45]),
        .O(\u1/u14/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__239_i_6
       (.I0(\u1/R13 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [43]),
        .I3(\u1/uk/K_r13 [9]),
        .O(\u1/u14/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__23_i_1
       (.I0(\u0/R2 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [22]),
        .I3(\u0/uk/K_r2 [0]),
        .O(\u0/u3/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__23_i_2
       (.I0(\u0/R2 [27]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [35]),
        .I3(\u0/uk/K_r2 [44]),
        .O(\u0/u3/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__23_i_3
       (.I0(\u0/R2 [26]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [2]),
        .I3(\u0/uk/K_r2 [35]),
        .O(\u0/u3/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__23_i_4
       (.I0(\u0/R2 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [45]),
        .I3(\u0/uk/K_r2 [50]),
        .O(\u0/u3/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__23_i_5
       (.I0(\u0/R2 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [14]),
        .I3(\u0/uk/K_r2 [23]),
        .O(\u0/u3/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__23_i_6
       (.I0(\u0/R2 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [37]),
        .I3(\u0/uk/K_r2 [15]),
        .O(\u0/u3/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__24
       (.I0(\u0/u3/X [17]),
        .I1(\u0/u3/X [16]),
        .I2(\u0/u3/X [15]),
        .I3(\u0/u3/X [14]),
        .I4(\u0/u3/X [18]),
        .I5(\u0/u3/X [13]),
        .O(\u0/out3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__240
       (.I0(\u1/u14/X [17]),
        .I1(\u1/u14/X [16]),
        .I2(\u1/u14/X [15]),
        .I3(\u1/u14/X [14]),
        .I4(\u1/u14/X [18]),
        .I5(\u1/u14/X [13]),
        .O(\u1/out14 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__240_i_1
       (.I0(\u1/R13 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [3]),
        .I3(\u1/uk/K_r13 [24]),
        .O(\u1/u14/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__240_i_2
       (.I0(\u1/R13 [11]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [20]),
        .I3(\u1/uk/K_r13 [41]),
        .O(\u1/u14/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__240_i_3
       (.I0(\u1/R13 [10]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [19]),
        .I3(\u1/uk/K_r13 [40]),
        .O(\u1/u14/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__240_i_4
       (.I0(\u1/R13 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [11]),
        .I3(\u1/uk/K_r13 [32]),
        .O(\u1/u14/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__240_i_5
       (.I0(\u1/R13 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [48]),
        .I3(\u1/uk/K_r13 [12]),
        .O(\u1/u14/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__240_i_6
       (.I0(\u1/R13 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [39]),
        .I3(\u1/uk/K_r13 [3]),
        .O(\u1/u14/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__241
       (.I0(\u1/u14/X [35]),
        .I1(\u1/u14/X [34]),
        .I2(\u1/u14/X [33]),
        .I3(\u1/u14/X [32]),
        .I4(\u1/u14/X [36]),
        .I5(\u1/u14/X [31]),
        .O(\u1/out14 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__241_i_1
       (.I0(\u1/R13 [24]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [21]),
        .I3(\u1/uk/K_r13 [42]),
        .O(\u1/u14/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__241_i_2
       (.I0(\u1/R13 [23]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [50]),
        .I3(\u1/uk/K_r13 [16]),
        .O(\u1/u14/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__241_i_3
       (.I0(\u1/R13 [22]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [37]),
        .I3(\u1/uk/K_r13 [31]),
        .O(\u1/u14/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__241_i_4
       (.I0(\u1/R13 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [15]),
        .I3(\u1/uk/K_r13 [36]),
        .O(\u1/u14/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__241_i_5
       (.I0(\u1/R13 [25]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [16]),
        .I3(\u1/uk/K_r13 [37]),
        .O(\u1/u14/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__241_i_6
       (.I0(\u1/R13 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [0]),
        .I3(\u1/uk/K_r13 [21]),
        .O(\u1/u14/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__242
       (.I0(\u1/u14/X [11]),
        .I1(\u1/u14/X [10]),
        .I2(\u1/u14/X [9]),
        .I3(\u1/u14/X [8]),
        .I4(\u1/u14/X [12]),
        .I5(\u1/u14/X [7]),
        .O(\u1/out14 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__242_i_1
       (.I0(\u1/R13 [8]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [25]),
        .I3(\u1/uk/K_r13 [46]),
        .O(\u1/u14/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__242_i_2
       (.I0(\u1/R13 [7]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [34]),
        .I3(\u1/uk/K_r13 [55]),
        .O(\u1/u14/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__242_i_3
       (.I0(\u1/R13 [6]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [40]),
        .I3(\u1/uk/K_r13 [4]),
        .O(\u1/u14/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__242_i_4
       (.I0(\u1/R13 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [17]),
        .I3(\u1/uk/K_r13 [13]),
        .O(\u1/u14/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__242_i_5
       (.I0(\u1/R13 [9]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [5]),
        .I3(\u1/uk/K_r13 [26]),
        .O(\u1/u14/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__242_i_6
       (.I0(\u1/R13 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [13]),
        .I3(\u1/uk/K_r13 [34]),
        .O(\u1/u14/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__243
       (.I0(\u1/u14/X [47]),
        .I1(\u1/u14/X [46]),
        .I2(\u1/u14/X [45]),
        .I3(\u1/u14/X [44]),
        .I4(\u1/u14/X [48]),
        .I5(\u1/u14/X [43]),
        .O(\u1/out14 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__243_i_1
       (.I0(\u1/R13 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [52]),
        .I3(\u1/uk/K_r13 [14]),
        .O(\u1/u14/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__243_i_2
       (.I0(\u1/R13 [31]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [42]),
        .I3(\u1/uk/K_r13 [8]),
        .O(\u1/u14/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__243_i_3
       (.I0(\u1/R13 [30]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [30]),
        .I3(\u1/uk/K_r13 [51]),
        .O(\u1/u14/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__243_i_4
       (.I0(\u1/R13 [29]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [29]),
        .I3(\u1/uk/K_r13 [50]),
        .O(\u1/u14/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__243_i_5
       (.I0(\u1/R13 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [14]),
        .I3(\u1/uk/K_r13 [35]),
        .O(\u1/u14/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__243_i_6
       (.I0(\u1/R13 [28]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [2]),
        .I3(\u1/uk/K_r13 [23]),
        .O(\u1/u14/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__244
       (.I0(\u1/u14/X [23]),
        .I1(\u1/u14/X [22]),
        .I2(\u1/u14/X [21]),
        .I3(\u1/u14/X [20]),
        .I4(\u1/u14/X [24]),
        .I5(\u1/u14/X [19]),
        .O(\u1/out14 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__244_i_1
       (.I0(\u1/R13 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [26]),
        .I3(\u1/uk/K_r13 [47]),
        .O(\u1/u14/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__244_i_2
       (.I0(\u1/R13 [15]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [18]),
        .I3(\u1/uk/K_r13 [39]),
        .O(\u1/u14/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__244_i_3
       (.I0(\u1/R13 [14]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [10]),
        .I3(\u1/uk/K_r13 [6]),
        .O(\u1/u14/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__244_i_4
       (.I0(\u1/R13 [13]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [41]),
        .I3(\u1/uk/K_r13 [5]),
        .O(\u1/u14/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__244_i_5
       (.I0(\u1/R13 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [6]),
        .I3(\u1/uk/K_r13 [27]),
        .O(\u1/u14/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__244_i_6
       (.I0(\u1/R13 [12]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [47]),
        .I3(\u1/uk/K_r13 [11]),
        .O(\u1/u14/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__245
       (.I0(\u1/u14/X [29]),
        .I1(\u1/u14/X [28]),
        .I2(\u1/u14/X [27]),
        .I3(\u1/u14/X [26]),
        .I4(\u1/u14/X [30]),
        .I5(\u1/u14/X [25]),
        .O(\u1/out14 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__245_i_1
       (.I0(\u1/R13 [20]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [9]),
        .I3(\u1/uk/K_r13 [30]),
        .O(\u1/u14/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__245_i_2
       (.I0(\u1/R13 [19]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [49]),
        .I3(\u1/uk/K_r13 [15]),
        .O(\u1/u14/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__245_i_3
       (.I0(\u1/R13 [18]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [7]),
        .I3(\u1/uk/K_r13 [28]),
        .O(\u1/u14/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__245_i_4
       (.I0(\u1/R13 [17]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [44]),
        .I3(\u1/uk/K_r13 [38]),
        .O(\u1/u14/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__245_i_5
       (.I0(\u1/R13 [21]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [38]),
        .I3(\u1/uk/K_r13 [0]),
        .O(\u1/u14/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__245_i_6
       (.I0(\u1/R13 [16]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [22]),
        .I3(\u1/uk/K_r13 [43]),
        .O(\u1/u14/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__246
       (.I0(\u1/u14/X [5]),
        .I1(\u1/u14/X [4]),
        .I2(\u1/u14/X [3]),
        .I3(\u1/u14/X [2]),
        .I4(\u1/u14/X [6]),
        .I5(\u1/u14/X [1]),
        .O(\u1/out14 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__246_i_1
       (.I0(\u1/R13 [4]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [24]),
        .I3(\u1/uk/K_r13 [20]),
        .O(\u1/u14/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__246_i_2
       (.I0(\u1/R13 [3]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [46]),
        .I3(\u1/uk/K_r13 [10]),
        .O(\u1/u14/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__246_i_3
       (.I0(\u1/R13 [2]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [12]),
        .I3(\u1/uk/K_r13 [33]),
        .O(\u1/u14/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__246_i_4
       (.I0(\u1/R13 [1]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [54]),
        .I3(\u1/uk/K_r13 [18]),
        .O(\u1/u14/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__246_i_5
       (.I0(\u1/R13 [5]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [27]),
        .I3(\u1/uk/K_r13 [48]),
        .O(\u1/u14/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__246_i_6
       (.I0(\u1/R13 [32]),
        .I1(decrypt),
        .I2(\u1/uk/K_r13 [33]),
        .I3(\u1/uk/K_r13 [54]),
        .O(\u1/u14/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__247
       (.I0(\u1/u15/X [41]),
        .I1(\u1/u15/X [40]),
        .I2(\u1/u15/X [39]),
        .I3(\u1/u15/X [38]),
        .I4(\u1/u15/X [42]),
        .I5(\u1/u15/X [37]),
        .O(\u1/out15 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__247_i_1
       (.I0(\u1/FP [60]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[35] ),
        .I3(\u1/uk/K_r14_reg_n_0_[42] ),
        .O(\u1/u15/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__247_i_2
       (.I0(\u1/FP [59]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[52] ),
        .I3(\u1/uk/K_r14_reg_n_0_ ),
        .O(\u1/u15/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__247_i_3
       (.I0(\u1/FP [58]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[15] ),
        .I3(\u1/uk/K_r14_reg_n_0_[22] ),
        .O(\u1/u15/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__247_i_4
       (.I0(\u1/FP [57]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[30] ),
        .I3(\u1/uk/K_r14_reg_n_0_[37] ),
        .O(\u1/u15/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__247_i_5
       (.I0(\u1/FP [61]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[31] ),
        .I3(\u1/uk/K_r14_reg_n_0_[38] ),
        .O(\u1/u15/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__247_i_6
       (.I0(\u1/FP [56]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[50] ),
        .I3(\u1/uk/K_r14_reg_n_0_[2] ),
        .O(\u1/u15/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__248
       (.I0(\u1/u15/X [17]),
        .I1(\u1/u15/X [16]),
        .I2(\u1/u15/X [15]),
        .I3(\u1/u15/X [14]),
        .I4(\u1/u15/X [18]),
        .I5(\u1/u15/X [13]),
        .O(\u1/out15 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__248_i_1
       (.I0(\u1/FP [44]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[10] ),
        .I3(\u1/uk/K_r14_reg_n_0_[17] ),
        .O(\u1/u15/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__248_i_2
       (.I0(\u1/FP [43]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[27] ),
        .I3(\u1/uk/K_r14_reg_n_0_[34] ),
        .O(\u1/u15/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__248_i_3
       (.I0(\u1/FP [42]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[26] ),
        .I3(\u1/uk/K_r14_reg_n_0_[33] ),
        .O(\u1/u15/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__248_i_4
       (.I0(\u1/FP [41]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[18] ),
        .I3(\u1/uk/K_r14_reg_n_0_[25] ),
        .O(\u1/u15/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__248_i_5
       (.I0(\u1/FP [45]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[55] ),
        .I3(\u1/uk/K_r14_reg_n_0_[5] ),
        .O(\u1/u15/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__248_i_6
       (.I0(\u1/FP [40]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[46] ),
        .I3(\u1/uk/K_r14_reg_n_0_[53] ),
        .O(\u1/u15/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__249
       (.I0(\u1/u15/X [35]),
        .I1(\u1/u15/X [34]),
        .I2(\u1/u15/X [33]),
        .I3(\u1/u15/X [32]),
        .I4(\u1/u15/X [36]),
        .I5(\u1/u15/X [31]),
        .O(\u1/out15 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__249_i_1
       (.I0(\u1/FP [56]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[28] ),
        .I3(\u1/uk/K_r14_reg_n_0_[35] ),
        .O(\u1/u15/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__249_i_2
       (.I0(\u1/FP [55]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[2] ),
        .I3(\u1/uk/K_r14_reg_n_0_[9] ),
        .O(\u1/u15/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__249_i_3
       (.I0(\u1/FP [54]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[44] ),
        .I3(\u1/uk/K_r14_reg_n_0_[51] ),
        .O(\u1/u15/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__249_i_4
       (.I0(\u1/FP [53]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[22] ),
        .I3(\u1/uk/K_r14_reg_n_0_[29] ),
        .O(\u1/u15/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__249_i_5
       (.I0(\u1/FP [57]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[23] ),
        .I3(\u1/uk/K_r14_reg_n_0_[30] ),
        .O(\u1/u15/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__249_i_6
       (.I0(\u1/FP [52]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[7] ),
        .I3(\u1/uk/K_r14_reg_n_0_[14] ),
        .O(\u1/u15/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__24_i_1
       (.I0(\u0/R2 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [27]),
        .I3(\u0/uk/K_r2 [32]),
        .O(\u0/u3/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__24_i_2
       (.I0(\u0/R2 [11]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [12]),
        .I3(\u0/uk/K_r2 [17]),
        .O(\u0/u3/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__24_i_3
       (.I0(\u0/R2 [10]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [11]),
        .I3(\u0/uk/K_r2 [48]),
        .O(\u0/u3/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__24_i_4
       (.I0(\u0/R2 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [3]),
        .I3(\u0/uk/K_r2 [40]),
        .O(\u0/u3/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__24_i_5
       (.I0(\u0/R2 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [40]),
        .I3(\u0/uk/K_r2 [20]),
        .O(\u0/u3/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__24_i_6
       (.I0(\u0/R2 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [6]),
        .I3(\u0/uk/K_r2 [11]),
        .O(\u0/u3/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__25
       (.I0(\u0/u3/X [35]),
        .I1(\u0/u3/X [34]),
        .I2(\u0/u3/X [33]),
        .I3(\u0/u3/X [32]),
        .I4(\u0/u3/X [36]),
        .I5(\u0/u3/X [31]),
        .O(\u0/out3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__250
       (.I0(\u1/u15/X [11]),
        .I1(\u1/u15/X [10]),
        .I2(\u1/u15/X [9]),
        .I3(\u1/u15/X [8]),
        .I4(\u1/u15/X [12]),
        .I5(\u1/u15/X [7]),
        .O(\u1/out15 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__250_i_1
       (.I0(\u1/FP [40]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[32] ),
        .I3(\u1/uk/K_r14_reg_n_0_[39] ),
        .O(\u1/u15/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__250_i_2
       (.I0(\u1/FP [39]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[41] ),
        .I3(\u1/uk/K_r14_reg_n_0_[48] ),
        .O(\u1/u15/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__250_i_3
       (.I0(\u1/FP [38]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[47] ),
        .I3(\u1/uk/K_r14_reg_n_0_[54] ),
        .O(\u1/u15/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__250_i_4
       (.I0(\u1/FP [37]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[24] ),
        .I3(\u1/uk/K_r14_reg_n_0_[6] ),
        .O(\u1/u15/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__250_i_5
       (.I0(\u1/FP [41]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[12] ),
        .I3(\u1/uk/K_r14_reg_n_0_[19] ),
        .O(\u1/u15/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__250_i_6
       (.I0(\u1/FP [36]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[20] ),
        .I3(\u1/uk/K_r14_reg_n_0_[27] ),
        .O(\u1/u15/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__251
       (.I0(\u1/u15/X [47]),
        .I1(\u1/u15/X [46]),
        .I2(\u1/u15/X [45]),
        .I3(\u1/u15/X [44]),
        .I4(\u1/u15/X [48]),
        .I5(\u1/u15/X [43]),
        .O(\u1/out15 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__251_i_1
       (.I0(\u1/FP [64]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_ ),
        .I3(\u1/uk/K_r14_reg_n_0_[7] ),
        .O(\u1/u15/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__251_i_2
       (.I0(\u1/FP [63]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[49] ),
        .I3(\u1/uk/K_r14_reg_n_0_[1] ),
        .O(\u1/u15/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__251_i_3
       (.I0(\u1/FP [62]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[37] ),
        .I3(\u1/uk/K_r14_reg_n_0_[44] ),
        .O(\u1/u15/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__251_i_4
       (.I0(\u1/FP [61]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[36] ),
        .I3(\u1/uk/K_r14_reg_n_0_[43] ),
        .O(\u1/u15/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__251_i_5
       (.I0(\u1/FP [33]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[21] ),
        .I3(\u1/uk/K_r14_reg_n_0_[28] ),
        .O(\u1/u15/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__251_i_6
       (.I0(\u1/FP [60]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[9] ),
        .I3(\u1/uk/K_r14_reg_n_0_[16] ),
        .O(\u1/u15/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__252
       (.I0(\u1/u15/X [23]),
        .I1(\u1/u15/X [22]),
        .I2(\u1/u15/X [21]),
        .I3(\u1/u15/X [20]),
        .I4(\u1/u15/X [24]),
        .I5(\u1/u15/X [19]),
        .O(\u1/out15 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__252_i_1
       (.I0(\u1/FP [48]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[33] ),
        .I3(\u1/uk/K_r14_reg_n_0_[40] ),
        .O(\u1/u15/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__252_i_2
       (.I0(\u1/FP [47]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[25] ),
        .I3(\u1/uk/K_r14_reg_n_0_[32] ),
        .O(\u1/u15/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__252_i_3
       (.I0(\u1/FP [46]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[17] ),
        .I3(\u1/uk/K_r14_reg_n_0_[24] ),
        .O(\u1/u15/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__252_i_4
       (.I0(\u1/FP [45]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[48] ),
        .I3(\u1/uk/K_r14_reg_n_0_[55] ),
        .O(\u1/u15/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__252_i_5
       (.I0(\u1/FP [49]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[13] ),
        .I3(\u1/uk/K_r14_reg_n_0_[20] ),
        .O(\u1/u15/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__252_i_6
       (.I0(\u1/FP [44]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[54] ),
        .I3(\u1/uk/K_r14_reg_n_0_[4] ),
        .O(\u1/u15/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__253
       (.I0(\u1/u15/X [29]),
        .I1(\u1/u15/X [28]),
        .I2(\u1/u15/X [27]),
        .I3(\u1/u15/X [26]),
        .I4(\u1/u15/X [30]),
        .I5(\u1/u15/X [25]),
        .O(\u1/out15 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__253_i_1
       (.I0(\u1/FP [52]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[16] ),
        .I3(\u1/uk/K_r14_reg_n_0_[23] ),
        .O(\u1/u15/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__253_i_2
       (.I0(\u1/FP [51]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[1] ),
        .I3(\u1/uk/K_r14_reg_n_0_[8] ),
        .O(\u1/u15/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__253_i_3
       (.I0(\u1/FP [50]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[14] ),
        .I3(\u1/uk/K_r14_reg_n_0_[21] ),
        .O(\u1/u15/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__253_i_4
       (.I0(\u1/FP [49]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[51] ),
        .I3(\u1/uk/K_r14_reg_n_0_[31] ),
        .O(\u1/u15/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__253_i_5
       (.I0(\u1/FP [53]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[45] ),
        .I3(\u1/uk/K_r14_reg_n_0_[52] ),
        .O(\u1/u15/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__253_i_6
       (.I0(\u1/FP [48]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[29] ),
        .I3(\u1/uk/K_r14_reg_n_0_[36] ),
        .O(\u1/u15/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__254
       (.I0(\u1/u15/X [5]),
        .I1(\u1/u15/X [4]),
        .I2(\u1/u15/X [3]),
        .I3(\u1/u15/X [2]),
        .I4(\u1/u15/X [6]),
        .I5(\u1/u15/X [1]),
        .O(\u1/out15 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__254_i_1
       (.I0(\u1/FP [36]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[6] ),
        .I3(\u1/uk/K_r14_reg_n_0_[13] ),
        .O(\u1/u15/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__254_i_2
       (.I0(\u1/FP [35]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[53] ),
        .I3(\u1/uk/K_r14_reg_n_0_[3] ),
        .O(\u1/u15/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__254_i_3
       (.I0(\u1/FP [34]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[19] ),
        .I3(\u1/uk/K_r14_reg_n_0_[26] ),
        .O(\u1/u15/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__254_i_4
       (.I0(\u1/FP [33]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[4] ),
        .I3(\u1/uk/K_r14_reg_n_0_[11] ),
        .O(\u1/u15/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__254_i_5
       (.I0(\u1/FP [37]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[34] ),
        .I3(\u1/uk/K_r14_reg_n_0_[41] ),
        .O(\u1/u15/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h596A)) 
    g0_b0__254_i_6
       (.I0(\u1/FP [64]),
        .I1(decrypt),
        .I2(\u1/uk/K_r14_reg_n_0_[40] ),
        .I3(\u1/uk/K_r14_reg_n_0_[47] ),
        .O(\u1/u15/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__255
       (.I0(\u2/u0/X [41]),
        .I1(\u2/u0/X [40]),
        .I2(\u2/u0/X [39]),
        .I3(\u2/u0/X [38]),
        .I4(\u2/u0/X [42]),
        .I5(\u2/u0/X [37]),
        .O(\u2/out0 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__255_i_1
       (.I0(\u2/IP [60]),
        .I1(decrypt),
        .I2(\u2/key_r [42]),
        .I3(\u2/key_r [35]),
        .O(\u2/u0/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__255_i_2
       (.I0(\u2/IP [59]),
        .I1(decrypt),
        .I2(\u2/key_r [0]),
        .I3(\u2/key_r [52]),
        .O(\u2/u0/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__255_i_3
       (.I0(\u2/IP [58]),
        .I1(decrypt),
        .I2(\u2/key_r [22]),
        .I3(\u2/key_r [15]),
        .O(\u2/u0/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__255_i_4
       (.I0(\u2/IP [57]),
        .I1(decrypt),
        .I2(\u2/key_r [37]),
        .I3(\u2/key_r [30]),
        .O(\u2/u0/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__255_i_5
       (.I0(\u2/IP [61]),
        .I1(decrypt),
        .I2(\u2/key_r [38]),
        .I3(\u2/key_r [31]),
        .O(\u2/u0/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__255_i_6
       (.I0(\u2/IP [56]),
        .I1(decrypt),
        .I2(\u2/key_r [2]),
        .I3(\u2/key_r [50]),
        .O(\u2/u0/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__256
       (.I0(\u2/u0/X [17]),
        .I1(\u2/u0/X [16]),
        .I2(\u2/u0/X [15]),
        .I3(\u2/u0/X [14]),
        .I4(\u2/u0/X [18]),
        .I5(\u2/u0/X [13]),
        .O(\u2/out0 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__256_i_1
       (.I0(\u2/IP [44]),
        .I1(decrypt),
        .I2(\u2/key_r [17]),
        .I3(\u2/key_r [10]),
        .O(\u2/u0/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__256_i_2
       (.I0(\u2/IP [43]),
        .I1(decrypt),
        .I2(\u2/key_r [34]),
        .I3(\u2/key_r [27]),
        .O(\u2/u0/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__256_i_3
       (.I0(\u2/IP [42]),
        .I1(decrypt),
        .I2(\u2/key_r [33]),
        .I3(\u2/key_r [26]),
        .O(\u2/u0/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__256_i_4
       (.I0(\u2/IP [41]),
        .I1(decrypt),
        .I2(\u2/key_r [25]),
        .I3(\u2/key_r [18]),
        .O(\u2/u0/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__256_i_5
       (.I0(\u2/IP [45]),
        .I1(decrypt),
        .I2(\u2/key_r [5]),
        .I3(\u2/key_r [55]),
        .O(\u2/u0/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__256_i_6
       (.I0(\u2/IP [40]),
        .I1(decrypt),
        .I2(\u2/key_r [53]),
        .I3(\u2/key_r [46]),
        .O(\u2/u0/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__257
       (.I0(\u2/u0/X [35]),
        .I1(\u2/u0/X [34]),
        .I2(\u2/u0/X [33]),
        .I3(\u2/u0/X [32]),
        .I4(\u2/u0/X [36]),
        .I5(\u2/u0/X [31]),
        .O(\u2/out0 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__257_i_1
       (.I0(\u2/IP [56]),
        .I1(decrypt),
        .I2(\u2/key_r [35]),
        .I3(\u2/key_r [28]),
        .O(\u2/u0/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__257_i_2
       (.I0(\u2/IP [55]),
        .I1(decrypt),
        .I2(\u2/key_r [9]),
        .I3(\u2/key_r [2]),
        .O(\u2/u0/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__257_i_3
       (.I0(\u2/IP [54]),
        .I1(decrypt),
        .I2(\u2/key_r [51]),
        .I3(\u2/key_r [44]),
        .O(\u2/u0/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__257_i_4
       (.I0(\u2/IP [53]),
        .I1(decrypt),
        .I2(\u2/key_r [29]),
        .I3(\u2/key_r [22]),
        .O(\u2/u0/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__257_i_5
       (.I0(\u2/IP [57]),
        .I1(decrypt),
        .I2(\u2/key_r [30]),
        .I3(\u2/key_r [23]),
        .O(\u2/u0/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__257_i_6
       (.I0(\u2/IP [52]),
        .I1(decrypt),
        .I2(\u2/key_r [14]),
        .I3(\u2/key_r [7]),
        .O(\u2/u0/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__258
       (.I0(\u2/u0/X [11]),
        .I1(\u2/u0/X [10]),
        .I2(\u2/u0/X [9]),
        .I3(\u2/u0/X [8]),
        .I4(\u2/u0/X [12]),
        .I5(\u2/u0/X [7]),
        .O(\u2/out0 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__258_i_1
       (.I0(\u2/IP [40]),
        .I1(decrypt),
        .I2(\u2/key_r [39]),
        .I3(\u2/key_r [32]),
        .O(\u2/u0/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__258_i_2
       (.I0(\u2/IP [39]),
        .I1(decrypt),
        .I2(\u2/key_r [48]),
        .I3(\u2/key_r [41]),
        .O(\u2/u0/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__258_i_3
       (.I0(\u2/IP [38]),
        .I1(decrypt),
        .I2(\u2/key_r [54]),
        .I3(\u2/key_r [47]),
        .O(\u2/u0/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__258_i_4
       (.I0(\u2/IP [37]),
        .I1(decrypt),
        .I2(\u2/key_r [6]),
        .I3(\u2/key_r [24]),
        .O(\u2/u0/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__258_i_5
       (.I0(\u2/IP [41]),
        .I1(decrypt),
        .I2(\u2/key_r [19]),
        .I3(\u2/key_r [12]),
        .O(\u2/u0/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__258_i_6
       (.I0(\u2/IP [36]),
        .I1(decrypt),
        .I2(\u2/key_r [27]),
        .I3(\u2/key_r [20]),
        .O(\u2/u0/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__259
       (.I0(\u2/u0/X [47]),
        .I1(\u2/u0/X [46]),
        .I2(\u2/u0/X [45]),
        .I3(\u2/u0/X [44]),
        .I4(\u2/u0/X [48]),
        .I5(\u2/u0/X [43]),
        .O(\u2/out0 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__259_i_1
       (.I0(\u2/IP [64]),
        .I1(decrypt),
        .I2(\u2/key_r [7]),
        .I3(\u2/key_r [0]),
        .O(\u2/u0/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__259_i_2
       (.I0(\u2/IP [63]),
        .I1(decrypt),
        .I2(\u2/key_r [1]),
        .I3(\u2/key_r [49]),
        .O(\u2/u0/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__259_i_3
       (.I0(\u2/IP [62]),
        .I1(decrypt),
        .I2(\u2/key_r [44]),
        .I3(\u2/key_r [37]),
        .O(\u2/u0/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__259_i_4
       (.I0(\u2/IP [61]),
        .I1(decrypt),
        .I2(\u2/key_r [43]),
        .I3(\u2/key_r [36]),
        .O(\u2/u0/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__259_i_5
       (.I0(\u2/IP [33]),
        .I1(decrypt),
        .I2(\u2/key_r [28]),
        .I3(\u2/key_r [21]),
        .O(\u2/u0/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__259_i_6
       (.I0(\u2/IP [60]),
        .I1(decrypt),
        .I2(\u2/key_r [16]),
        .I3(\u2/key_r [9]),
        .O(\u2/u0/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__25_i_1
       (.I0(\u0/R2 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [15]),
        .I3(\u0/uk/K_r2 [52]),
        .O(\u0/u3/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__25_i_2
       (.I0(\u0/R2 [23]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [44]),
        .I3(\u0/uk/K_r2 [22]),
        .O(\u0/u3/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__25_i_3
       (.I0(\u0/R2 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [0]),
        .I3(\u0/uk/K_r2 [9]),
        .O(\u0/u3/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__25_i_4
       (.I0(\u0/R2 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [9]),
        .I3(\u0/uk/K_r2 [42]),
        .O(\u0/u3/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__25_i_5
       (.I0(\u0/R2 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [38]),
        .I3(\u0/uk/K_r2 [43]),
        .O(\u0/u3/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__25_i_6
       (.I0(\u0/R2 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [49]),
        .I3(\u0/uk/K_r2 [31]),
        .O(\u0/u3/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__26
       (.I0(\u0/u3/X [11]),
        .I1(\u0/u3/X [10]),
        .I2(\u0/u3/X [9]),
        .I3(\u0/u3/X [8]),
        .I4(\u0/u3/X [12]),
        .I5(\u0/u3/X [7]),
        .O(\u0/out3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__260
       (.I0(\u2/u0/X [23]),
        .I1(\u2/u0/X [22]),
        .I2(\u2/u0/X [21]),
        .I3(\u2/u0/X [20]),
        .I4(\u2/u0/X [24]),
        .I5(\u2/u0/X [19]),
        .O(\u2/out0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__260_i_1
       (.I0(\u2/IP [48]),
        .I1(decrypt),
        .I2(\u2/key_r [40]),
        .I3(\u2/key_r [33]),
        .O(\u2/u0/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__260_i_2
       (.I0(\u2/IP [47]),
        .I1(decrypt),
        .I2(\u2/key_r [32]),
        .I3(\u2/key_r [25]),
        .O(\u2/u0/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__260_i_3
       (.I0(\u2/IP [46]),
        .I1(decrypt),
        .I2(\u2/key_r [24]),
        .I3(\u2/key_r [17]),
        .O(\u2/u0/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__260_i_4
       (.I0(\u2/IP [45]),
        .I1(decrypt),
        .I2(\u2/key_r [55]),
        .I3(\u2/key_r [48]),
        .O(\u2/u0/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__260_i_5
       (.I0(\u2/IP [49]),
        .I1(decrypt),
        .I2(\u2/key_r [20]),
        .I3(\u2/key_r [13]),
        .O(\u2/u0/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__260_i_6
       (.I0(\u2/IP [44]),
        .I1(decrypt),
        .I2(\u2/key_r [4]),
        .I3(\u2/key_r [54]),
        .O(\u2/u0/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__261
       (.I0(\u2/u0/X [29]),
        .I1(\u2/u0/X [28]),
        .I2(\u2/u0/X [27]),
        .I3(\u2/u0/X [26]),
        .I4(\u2/u0/X [30]),
        .I5(\u2/u0/X [25]),
        .O(\u2/out0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__261_i_1
       (.I0(\u2/IP [52]),
        .I1(decrypt),
        .I2(\u2/key_r [23]),
        .I3(\u2/key_r [16]),
        .O(\u2/u0/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__261_i_2
       (.I0(\u2/IP [51]),
        .I1(decrypt),
        .I2(\u2/key_r [8]),
        .I3(\u2/key_r [1]),
        .O(\u2/u0/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__261_i_3
       (.I0(\u2/IP [50]),
        .I1(decrypt),
        .I2(\u2/key_r [21]),
        .I3(\u2/key_r [14]),
        .O(\u2/u0/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__261_i_4
       (.I0(\u2/IP [49]),
        .I1(decrypt),
        .I2(\u2/key_r [31]),
        .I3(\u2/key_r [51]),
        .O(\u2/u0/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__261_i_5
       (.I0(\u2/IP [53]),
        .I1(decrypt),
        .I2(\u2/key_r [52]),
        .I3(\u2/key_r [45]),
        .O(\u2/u0/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__261_i_6
       (.I0(\u2/IP [48]),
        .I1(decrypt),
        .I2(\u2/key_r [36]),
        .I3(\u2/key_r [29]),
        .O(\u2/u0/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__262
       (.I0(\u2/u0/X [5]),
        .I1(\u2/u0/X [4]),
        .I2(\u2/u0/X [3]),
        .I3(\u2/u0/X [2]),
        .I4(\u2/u0/X [6]),
        .I5(\u2/u0/X [1]),
        .O(\u2/out0 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__262_i_1
       (.I0(\u2/IP [36]),
        .I1(decrypt),
        .I2(\u2/key_r [13]),
        .I3(\u2/key_r [6]),
        .O(\u2/u0/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__262_i_2
       (.I0(\u2/IP [35]),
        .I1(decrypt),
        .I2(\u2/key_r [3]),
        .I3(\u2/key_r [53]),
        .O(\u2/u0/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__262_i_3
       (.I0(\u2/IP [34]),
        .I1(decrypt),
        .I2(\u2/key_r [26]),
        .I3(\u2/key_r [19]),
        .O(\u2/u0/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__262_i_4
       (.I0(\u2/IP [33]),
        .I1(decrypt),
        .I2(\u2/key_r [11]),
        .I3(\u2/key_r [4]),
        .O(\u2/u0/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__262_i_5
       (.I0(\u2/IP [37]),
        .I1(decrypt),
        .I2(\u2/key_r [41]),
        .I3(\u2/key_r [34]),
        .O(\u2/u0/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__262_i_6
       (.I0(\u2/IP [64]),
        .I1(decrypt),
        .I2(\u2/key_r [47]),
        .I3(\u2/key_r [40]),
        .O(\u2/u0/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__263
       (.I0(\u2/u1/X [41]),
        .I1(\u2/u1/X [40]),
        .I2(\u2/u1/X [39]),
        .I3(\u2/u1/X [38]),
        .I4(\u2/u1/X [42]),
        .I5(\u2/u1/X [37]),
        .O(\u2/out1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__263_i_1
       (.I0(\u2/R0 [28]),
        .I1(decrypt),
        .I2(\u2/uk/p_34_in ),
        .I3(\u2/uk/p_20_in ),
        .O(\u2/u1/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__263_i_2
       (.I0(\u2/R0 [27]),
        .I1(decrypt),
        .I2(\u2/uk/p_21_in ),
        .I3(\u2/uk/p_33_in ),
        .O(\u2/u1/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__263_i_3
       (.I0(\u2/R0 [26]),
        .I1(decrypt),
        .I2(\u2/uk/p_31_in ),
        .I3(\u2/uk/p_32_in ),
        .O(\u2/u1/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__263_i_4
       (.I0(\u2/R0 [25]),
        .I1(decrypt),
        .I2(\u2/uk/p_19_in ),
        .I3(\u2/uk/p_30_in ),
        .O(\u2/u1/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__263_i_5
       (.I0(\u2/R0 [29]),
        .I1(decrypt),
        .I2(\u2/uk/p_33_in ),
        .I3(\u2/uk/p_35_in ),
        .O(\u2/u1/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__263_i_6
       (.I0(\u2/R0 [24]),
        .I1(decrypt),
        .I2(\u2/uk/p_23_in ),
        .I3(\u2/uk/p_17_in ),
        .O(\u2/u1/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__264
       (.I0(\u2/u1/X [17]),
        .I1(\u2/u1/X [16]),
        .I2(\u2/u1/X [15]),
        .I3(\u2/u1/X [14]),
        .I4(\u2/u1/X [18]),
        .I5(\u2/u1/X [13]),
        .O(\u2/out1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__264_i_1
       (.I0(\u2/R0 [12]),
        .I1(decrypt),
        .I2(\u2/uk/p_3_in ),
        .I3(\u2/uk/p_11_in ),
        .O(\u2/u1/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__264_i_2
       (.I0(\u2/R0 [11]),
        .I1(decrypt),
        .I2(\u2/uk/p_13_in ),
        .I3(\u2/uk/p_2_in ),
        .O(\u2/u1/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__264_i_3
       (.I0(\u2/R0 [10]),
        .I1(decrypt),
        .I2(\u2/uk/p_8_in ),
        .I3(\u2/uk/K_r0_reg_n_0_[19] ),
        .O(\u2/u1/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__264_i_4
       (.I0(\u2/R0 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r0_reg_n_0_[32] ),
        .I3(\u2/uk/p_14_in ),
        .O(\u2/u1/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__264_i_5
       (.I0(\u2/R0 [13]),
        .I1(decrypt),
        .I2(\u2/uk/p_38_in ),
        .I3(\u2/uk/p_4_in ),
        .O(\u2/u1/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__264_i_6
       (.I0(\u2/R0 [8]),
        .I1(decrypt),
        .I2(\u2/uk/p_11_in ),
        .I3(\u2/uk/p_12_in ),
        .O(\u2/u1/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__265
       (.I0(\u2/u1/X [35]),
        .I1(\u2/u1/X [34]),
        .I2(\u2/u1/X [33]),
        .I3(\u2/u1/X [32]),
        .I4(\u2/u1/X [36]),
        .I5(\u2/u1/X [31]),
        .O(\u2/out1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__265_i_1
       (.I0(\u2/R0 [24]),
        .I1(decrypt),
        .I2(\u2/uk/p_29_in ),
        .I3(\u2/uk/p_24_in ),
        .O(\u2/u1/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__265_i_2
       (.I0(\u2/R0 [23]),
        .I1(decrypt),
        .I2(\u2/uk/p_27_in ),
        .I3(\u2/uk/p_28_in ),
        .O(\u2/u1/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__265_i_3
       (.I0(\u2/R0 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r0_reg_n_0_[31] ),
        .I3(\u2/uk/p_26_in ),
        .O(\u2/u1/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__265_i_4
       (.I0(\u2/R0 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r0_reg_n_0_[36] ),
        .I3(\u2/uk/p_25_in ),
        .O(\u2/u1/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__265_i_5
       (.I0(\u2/R0 [25]),
        .I1(decrypt),
        .I2(\u2/uk/p_26_in ),
        .I3(\u2/uk/p_27_in ),
        .O(\u2/u1/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__265_i_6
       (.I0(\u2/R0 [20]),
        .I1(decrypt),
        .I2(\u2/uk/p_24_in ),
        .I3(\u2/uk/K_r0_reg_n_0_ ),
        .O(\u2/u1/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__266
       (.I0(\u2/u1/X [11]),
        .I1(\u2/u1/X [10]),
        .I2(\u2/u1/X [9]),
        .I3(\u2/u1/X [8]),
        .I4(\u2/u1/X [12]),
        .I5(\u2/u1/X [7]),
        .O(\u2/out1 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__266_i_1
       (.I0(\u2/R0 [8]),
        .I1(decrypt),
        .I2(\u2/uk/p_1_in ),
        .I3(\u2/uk/K_r0_reg_n_0_[25] ),
        .O(\u2/u1/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__266_i_2
       (.I0(\u2/R0 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r0_reg_n_0_[55] ),
        .I3(\u2/uk/p_6_in ),
        .O(\u2/u1/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__266_i_3
       (.I0(\u2/R0 [6]),
        .I1(decrypt),
        .I2(\u2/uk/K_r0_reg_n_0_[4] ),
        .I3(\u2/uk/p_8_in ),
        .O(\u2/u1/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__266_i_4
       (.I0(\u2/R0 [5]),
        .I1(decrypt),
        .I2(\u2/uk/p_7_in ),
        .I3(\u2/uk/K_r0_reg_n_0_[17] ),
        .O(\u2/u1/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__266_i_5
       (.I0(\u2/R0 [9]),
        .I1(decrypt),
        .I2(\u2/uk/p_9_in ),
        .I3(\u2/uk/p_10_in ),
        .O(\u2/u1/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__266_i_6
       (.I0(\u2/R0 [4]),
        .I1(decrypt),
        .I2(\u2/uk/p_6_in ),
        .I3(\u2/uk/p_7_in ),
        .O(\u2/u1/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__267
       (.I0(\u2/u1/X [47]),
        .I1(\u2/u1/X [46]),
        .I2(\u2/u1/X [45]),
        .I3(\u2/u1/X [44]),
        .I4(\u2/u1/X [48]),
        .I5(\u2/u1/X [43]),
        .O(\u2/out1 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__267_i_1
       (.I0(\u2/R0 [32]),
        .I1(decrypt),
        .I2(\u2/uk/p_36_in ),
        .I3(\u2/uk/K_r0_reg_n_0_[52] ),
        .O(\u2/u1/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__267_i_2
       (.I0(\u2/R0 [31]),
        .I1(decrypt),
        .I2(\u2/uk/p_32_in ),
        .I3(\u2/uk/p_29_in ),
        .O(\u2/u1/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__267_i_3
       (.I0(\u2/R0 [30]),
        .I1(decrypt),
        .I2(\u2/uk/p_35_in ),
        .I3(\u2/uk/p_22_in ),
        .O(\u2/u1/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__267_i_4
       (.I0(\u2/R0 [29]),
        .I1(decrypt),
        .I2(\u2/uk/p_28_in ),
        .I3(\u2/uk/p_31_in ),
        .O(\u2/u1/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__267_i_5
       (.I0(\u2/R0 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r0_reg_n_0_[35] ),
        .I3(\u2/uk/p_36_in ),
        .O(\u2/u1/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__267_i_6
       (.I0(\u2/R0 [28]),
        .I1(decrypt),
        .I2(\u2/uk/p_30_in ),
        .I3(\u2/uk/K_r0_reg_n_0_[2] ),
        .O(\u2/u1/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__268
       (.I0(\u2/u1/X [23]),
        .I1(\u2/u1/X [22]),
        .I2(\u2/u1/X [21]),
        .I3(\u2/u1/X [20]),
        .I4(\u2/u1/X [24]),
        .I5(\u2/u1/X [19]),
        .O(\u2/out1 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__268_i_1
       (.I0(\u2/R0 [16]),
        .I1(decrypt),
        .I2(\u2/uk/p_15_in ),
        .I3(\u2/uk/p_9_in ),
        .O(\u2/u1/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__268_i_2
       (.I0(\u2/R0 [15]),
        .I1(decrypt),
        .I2(\u2/uk/p_12_in ),
        .I3(\u2/uk/p_37_in ),
        .O(\u2/u1/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__268_i_3
       (.I0(\u2/R0 [14]),
        .I1(decrypt),
        .I2(\u2/uk/p_16_in ),
        .I3(\u2/uk/p_0_in ),
        .O(\u2/u1/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__268_i_4
       (.I0(\u2/R0 [13]),
        .I1(decrypt),
        .I2(\u2/uk/p_10_in ),
        .I3(\u2/uk/p_13_in ),
        .O(\u2/u1/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__268_i_5
       (.I0(\u2/R0 [17]),
        .I1(decrypt),
        .I2(\u2/uk/p_5_in ),
        .I3(\u2/uk/p_16_in ),
        .O(\u2/u1/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__268_i_6
       (.I0(\u2/R0 [12]),
        .I1(decrypt),
        .I2(\u2/uk/p_14_in ),
        .I3(\u2/uk/p_15_in ),
        .O(\u2/u1/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__269
       (.I0(\u2/u1/X [29]),
        .I1(\u2/u1/X [28]),
        .I2(\u2/u1/X [27]),
        .I3(\u2/u1/X [26]),
        .I4(\u2/u1/X [30]),
        .I5(\u2/u1/X [25]),
        .O(\u2/out1 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__269_i_1
       (.I0(\u2/R0 [20]),
        .I1(decrypt),
        .I2(\u2/uk/p_22_in ),
        .I3(\u2/uk/p_23_in ),
        .O(\u2/u1/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__269_i_2
       (.I0(\u2/R0 [19]),
        .I1(decrypt),
        .I2(\u2/uk/p_25_in ),
        .I3(\u2/uk/p_34_in ),
        .O(\u2/u1/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__269_i_3
       (.I0(\u2/R0 [18]),
        .I1(decrypt),
        .I2(\u2/uk/p_20_in ),
        .I3(\u2/uk/p_21_in ),
        .O(\u2/u1/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__269_i_4
       (.I0(\u2/R0 [17]),
        .I1(decrypt),
        .I2(\u2/uk/p_18_in ),
        .I3(\u2/uk/p_19_in ),
        .O(\u2/u1/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__269_i_5
       (.I0(\u2/R0 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r0_reg_n_0_ ),
        .I3(\u2/uk/p_18_in ),
        .O(\u2/u1/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__269_i_6
       (.I0(\u2/R0 [16]),
        .I1(decrypt),
        .I2(\u2/uk/p_17_in ),
        .I3(\u2/uk/K_r0_reg_n_0_[22] ),
        .O(\u2/u1/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__26_i_1
       (.I0(\u0/R2 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [17]),
        .I3(\u0/uk/K_r2 [54]),
        .O(\u0/u3/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__26_i_2
       (.I0(\u0/R2 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [26]),
        .I3(\u0/uk/K_r2 [6]),
        .O(\u0/u3/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__26_i_3
       (.I0(\u0/R2 [6]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [32]),
        .I3(\u0/uk/K_r2 [12]),
        .O(\u0/u3/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__26_i_4
       (.I0(\u0/R2 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [41]),
        .I3(\u0/uk/K_r2 [46]),
        .O(\u0/u3/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__26_i_5
       (.I0(\u0/R2 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [54]),
        .I3(\u0/uk/K_r2 [34]),
        .O(\u0/u3/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__26_i_6
       (.I0(\u0/R2 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [5]),
        .I3(\u0/uk/K_r2 [10]),
        .O(\u0/u3/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__27
       (.I0(\u0/u3/X [47]),
        .I1(\u0/u3/X [46]),
        .I2(\u0/u3/X [45]),
        .I3(\u0/u3/X [44]),
        .I4(\u0/u3/X [48]),
        .I5(\u0/u3/X [43]),
        .O(\u0/out3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__270
       (.I0(\u2/u1/X [5]),
        .I1(\u2/u1/X [4]),
        .I2(\u2/u1/X [3]),
        .I3(\u2/u1/X [2]),
        .I4(\u2/u1/X [6]),
        .I5(\u2/u1/X [1]),
        .O(\u2/out1 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__270_i_1
       (.I0(\u2/R0 [4]),
        .I1(decrypt),
        .I2(\u2/uk/p_2_in ),
        .I3(\u2/uk/p_3_in ),
        .O(\u2/u1/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__270_i_2
       (.I0(\u2/R0 [3]),
        .I1(decrypt),
        .I2(\u2/uk/p_0_in ),
        .I3(\u2/uk/p_1_in ),
        .O(\u2/u1/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__270_i_3
       (.I0(\u2/R0 [2]),
        .I1(decrypt),
        .I2(\u2/uk/p_39_in ),
        .I3(\u2/uk/p_38_in ),
        .O(\u2/u1/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__270_i_4
       (.I0(\u2/R0 [1]),
        .I1(decrypt),
        .I2(\u2/uk/p_37_in ),
        .I3(\u2/uk/p_40_in ),
        .O(\u2/u1/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__270_i_5
       (.I0(\u2/R0 [5]),
        .I1(decrypt),
        .I2(\u2/uk/p_4_in ),
        .I3(\u2/uk/p_5_in ),
        .O(\u2/u1/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__270_i_6
       (.I0(\u2/R0 [32]),
        .I1(decrypt),
        .I2(\u2/uk/p_40_in ),
        .I3(\u2/uk/p_39_in ),
        .O(\u2/u1/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__271
       (.I0(\u2/u2/X [41]),
        .I1(\u2/u2/X [40]),
        .I2(\u2/u2/X [39]),
        .I3(\u2/u2/X [38]),
        .I4(\u2/u2/X [42]),
        .I5(\u2/u2/X [37]),
        .O(\u2/out2 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__271_i_1
       (.I0(\u2/R1 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [8]),
        .I3(\u2/uk/K_r1 [14]),
        .O(\u2/u2/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__271_i_2
       (.I0(\u2/R1 [27]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [21]),
        .I3(\u2/uk/K_r1 [31]),
        .O(\u2/u2/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__271_i_3
       (.I0(\u2/R1 [26]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [43]),
        .I3(\u2/uk/K_r1 [49]),
        .O(\u2/u2/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__271_i_4
       (.I0(\u2/R1 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [31]),
        .I3(\u2/uk/K_r1 [9]),
        .O(\u2/u2/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__271_i_5
       (.I0(\u2/R1 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [0]),
        .I3(\u2/uk/K_r1 [37]),
        .O(\u2/u2/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__271_i_6
       (.I0(\u2/R1 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [23]),
        .I3(\u2/uk/K_r1 [29]),
        .O(\u2/u2/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__272
       (.I0(\u2/u2/X [17]),
        .I1(\u2/u2/X [16]),
        .I2(\u2/u2/X [15]),
        .I3(\u2/u2/X [14]),
        .I4(\u2/u2/X [18]),
        .I5(\u2/u2/X [13]),
        .O(\u2/out2 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__272_i_1
       (.I0(\u2/R1 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [13]),
        .I3(\u2/uk/K_r1 [46]),
        .O(\u2/u2/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__272_i_2
       (.I0(\u2/R1 [11]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [55]),
        .I3(\u2/uk/K_r1 [6]),
        .O(\u2/u2/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__272_i_3
       (.I0(\u2/R1 [10]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [54]),
        .I3(\u2/uk/K_r1 [5]),
        .O(\u2/u2/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__272_i_4
       (.I0(\u2/R1 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [46]),
        .I3(\u2/uk/K_r1 [54]),
        .O(\u2/u2/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__272_i_5
       (.I0(\u2/R1 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [26]),
        .I3(\u2/uk/K_r1 [34]),
        .O(\u2/u2/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__272_i_6
       (.I0(\u2/R1 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [17]),
        .I3(\u2/uk/K_r1 [25]),
        .O(\u2/u2/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__273
       (.I0(\u2/u2/X [35]),
        .I1(\u2/u2/X [34]),
        .I2(\u2/u2/X [33]),
        .I3(\u2/u2/X [32]),
        .I4(\u2/u2/X [36]),
        .I5(\u2/u2/X [31]),
        .O(\u2/out2 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__273_i_1
       (.I0(\u2/R1 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [1]),
        .I3(\u2/uk/K_r1 [7]),
        .O(\u2/u2/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__273_i_2
       (.I0(\u2/R1 [23]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [30]),
        .I3(\u2/uk/K_r1 [36]),
        .O(\u2/u2/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__273_i_3
       (.I0(\u2/R1 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [45]),
        .I3(\u2/uk/K_r1 [23]),
        .O(\u2/u2/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__273_i_4
       (.I0(\u2/R1 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [50]),
        .I3(\u2/uk/K_r1 [1]),
        .O(\u2/u2/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__273_i_5
       (.I0(\u2/R1 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [51]),
        .I3(\u2/uk/K_r1 [2]),
        .O(\u2/u2/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__273_i_6
       (.I0(\u2/R1 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [35]),
        .I3(\u2/uk/K_r1 [45]),
        .O(\u2/u2/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__274
       (.I0(\u2/u2/X [11]),
        .I1(\u2/u2/X [10]),
        .I2(\u2/u2/X [9]),
        .I3(\u2/u2/X [8]),
        .I4(\u2/u2/X [12]),
        .I5(\u2/u2/X [7]),
        .O(\u2/out2 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__274_i_1
       (.I0(\u2/R1 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [3]),
        .I3(\u2/uk/K_r1 [11]),
        .O(\u2/u2/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__274_i_2
       (.I0(\u2/R1 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [12]),
        .I3(\u2/uk/K_r1 [20]),
        .O(\u2/u2/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__274_i_3
       (.I0(\u2/R1 [6]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [18]),
        .I3(\u2/uk/K_r1 [26]),
        .O(\u2/u2/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__274_i_4
       (.I0(\u2/R1 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [27]),
        .I3(\u2/uk/K_r1 [3]),
        .O(\u2/u2/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__274_i_5
       (.I0(\u2/R1 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [40]),
        .I3(\u2/uk/K_r1 [48]),
        .O(\u2/u2/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__274_i_6
       (.I0(\u2/R1 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [48]),
        .I3(\u2/uk/K_r1 [24]),
        .O(\u2/u2/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__275
       (.I0(\u2/u2/X [47]),
        .I1(\u2/u2/X [46]),
        .I2(\u2/u2/X [45]),
        .I3(\u2/u2/X [44]),
        .I4(\u2/u2/X [48]),
        .I5(\u2/u2/X [43]),
        .O(\u2/out2 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__275_i_1
       (.I0(\u2/R1 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [28]),
        .I3(\u2/uk/K_r1 [38]),
        .O(\u2/u2/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__275_i_2
       (.I0(\u2/R1 [31]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [22]),
        .I3(\u2/uk/K_r1 [28]),
        .O(\u2/u2/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__275_i_3
       (.I0(\u2/R1 [30]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [38]),
        .I3(\u2/uk/K_r1 [16]),
        .O(\u2/u2/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__275_i_4
       (.I0(\u2/R1 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [9]),
        .I3(\u2/uk/K_r1 [15]),
        .O(\u2/u2/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__275_i_5
       (.I0(\u2/R1 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [49]),
        .I3(\u2/uk/K_r1 [0]),
        .O(\u2/u2/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__275_i_6
       (.I0(\u2/R1 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [37]),
        .I3(\u2/uk/K_r1 [43]),
        .O(\u2/u2/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__276
       (.I0(\u2/u2/X [23]),
        .I1(\u2/u2/X [22]),
        .I2(\u2/u2/X [21]),
        .I3(\u2/u2/X [20]),
        .I4(\u2/u2/X [24]),
        .I5(\u2/u2/X [19]),
        .O(\u2/out2 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__276_i_1
       (.I0(\u2/R1 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [4]),
        .I3(\u2/uk/K_r1 [12]),
        .O(\u2/u2/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__276_i_2
       (.I0(\u2/R1 [15]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [53]),
        .I3(\u2/uk/K_r1 [4]),
        .O(\u2/u2/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__276_i_3
       (.I0(\u2/R1 [14]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [20]),
        .I3(\u2/uk/K_r1 [53]),
        .O(\u2/u2/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__276_i_4
       (.I0(\u2/R1 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [19]),
        .I3(\u2/uk/K_r1 [27]),
        .O(\u2/u2/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__276_i_5
       (.I0(\u2/R1 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [41]),
        .I3(\u2/uk/K_r1 [17]),
        .O(\u2/u2/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__276_i_6
       (.I0(\u2/R1 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [25]),
        .I3(\u2/uk/K_r1 [33]),
        .O(\u2/u2/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__277
       (.I0(\u2/u2/X [29]),
        .I1(\u2/u2/X [28]),
        .I2(\u2/u2/X [27]),
        .I3(\u2/u2/X [26]),
        .I4(\u2/u2/X [30]),
        .I5(\u2/u2/X [25]),
        .O(\u2/out2 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__277_i_1
       (.I0(\u2/R1 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [44]),
        .I3(\u2/uk/K_r1 [50]),
        .O(\u2/u2/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__277_i_2
       (.I0(\u2/R1 [19]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [29]),
        .I3(\u2/uk/K_r1 [35]),
        .O(\u2/u2/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__277_i_3
       (.I0(\u2/R1 [18]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [42]),
        .I3(\u2/uk/K_r1 [52]),
        .O(\u2/u2/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__277_i_4
       (.I0(\u2/R1 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [52]),
        .I3(\u2/uk/K_r1 [30]),
        .O(\u2/u2/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__277_i_5
       (.I0(\u2/R1 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [14]),
        .I3(\u2/uk/K_r1 [51]),
        .O(\u2/u2/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__277_i_6
       (.I0(\u2/R1 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [2]),
        .I3(\u2/uk/K_r1 [8]),
        .O(\u2/u2/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__278
       (.I0(\u2/u2/X [5]),
        .I1(\u2/u2/X [4]),
        .I2(\u2/u2/X [3]),
        .I3(\u2/u2/X [2]),
        .I4(\u2/u2/X [6]),
        .I5(\u2/u2/X [1]),
        .O(\u2/out2 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__278_i_1
       (.I0(\u2/R1 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [34]),
        .I3(\u2/uk/K_r1 [10]),
        .O(\u2/u2/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__278_i_2
       (.I0(\u2/R1 [3]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [24]),
        .I3(\u2/uk/K_r1 [32]),
        .O(\u2/u2/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__278_i_3
       (.I0(\u2/R1 [2]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [47]),
        .I3(\u2/uk/K_r1 [55]),
        .O(\u2/u2/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__278_i_4
       (.I0(\u2/R1 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [32]),
        .I3(\u2/uk/K_r1 [40]),
        .O(\u2/u2/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__278_i_5
       (.I0(\u2/R1 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [5]),
        .I3(\u2/uk/K_r1 [13]),
        .O(\u2/u2/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__278_i_6
       (.I0(\u2/R1 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r1 [11]),
        .I3(\u2/uk/K_r1 [19]),
        .O(\u2/u2/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__279
       (.I0(\u2/u3/X [41]),
        .I1(\u2/u3/X [40]),
        .I2(\u2/u3/X [39]),
        .I3(\u2/u3/X [38]),
        .I4(\u2/u3/X [42]),
        .I5(\u2/u3/X [37]),
        .O(\u2/out3 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__279_i_1
       (.I0(\u2/R2 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [22]),
        .I3(\u2/uk/K_r2 [0]),
        .O(\u2/u3/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__279_i_2
       (.I0(\u2/R2 [27]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [35]),
        .I3(\u2/uk/K_r2 [44]),
        .O(\u2/u3/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__279_i_3
       (.I0(\u2/R2 [26]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [2]),
        .I3(\u2/uk/K_r2 [35]),
        .O(\u2/u3/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__279_i_4
       (.I0(\u2/R2 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [45]),
        .I3(\u2/uk/K_r2 [50]),
        .O(\u2/u3/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__279_i_5
       (.I0(\u2/R2 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [14]),
        .I3(\u2/uk/K_r2 [23]),
        .O(\u2/u3/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__279_i_6
       (.I0(\u2/R2 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [37]),
        .I3(\u2/uk/K_r2 [15]),
        .O(\u2/u3/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__27_i_1
       (.I0(\u0/R2 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [42]),
        .I3(\u0/uk/K_r2 [51]),
        .O(\u0/u3/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__27_i_2
       (.I0(\u0/R2 [31]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [36]),
        .I3(\u0/uk/K_r2 [14]),
        .O(\u0/u3/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__27_i_3
       (.I0(\u0/R2 [30]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [52]),
        .I3(\u0/uk/K_r2 [2]),
        .O(\u0/u3/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__27_i_4
       (.I0(\u0/R2 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [23]),
        .I3(\u0/uk/K_r2 [1]),
        .O(\u0/u3/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__27_i_5
       (.I0(\u0/R2 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [8]),
        .I3(\u0/uk/K_r2 [45]),
        .O(\u0/u3/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__27_i_6
       (.I0(\u0/R2 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [51]),
        .I3(\u0/uk/K_r2 [29]),
        .O(\u0/u3/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__28
       (.I0(\u0/u3/X [23]),
        .I1(\u0/u3/X [22]),
        .I2(\u0/u3/X [21]),
        .I3(\u0/u3/X [20]),
        .I4(\u0/u3/X [24]),
        .I5(\u0/u3/X [19]),
        .O(\u0/out3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__280
       (.I0(\u2/u3/X [17]),
        .I1(\u2/u3/X [16]),
        .I2(\u2/u3/X [15]),
        .I3(\u2/u3/X [14]),
        .I4(\u2/u3/X [18]),
        .I5(\u2/u3/X [13]),
        .O(\u2/out3 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__280_i_1
       (.I0(\u2/R2 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [27]),
        .I3(\u2/uk/K_r2 [32]),
        .O(\u2/u3/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__280_i_2
       (.I0(\u2/R2 [11]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [12]),
        .I3(\u2/uk/K_r2 [17]),
        .O(\u2/u3/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__280_i_3
       (.I0(\u2/R2 [10]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [11]),
        .I3(\u2/uk/K_r2 [48]),
        .O(\u2/u3/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__280_i_4
       (.I0(\u2/R2 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [3]),
        .I3(\u2/uk/K_r2 [40]),
        .O(\u2/u3/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__280_i_5
       (.I0(\u2/R2 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [40]),
        .I3(\u2/uk/K_r2 [20]),
        .O(\u2/u3/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__280_i_6
       (.I0(\u2/R2 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [6]),
        .I3(\u2/uk/K_r2 [11]),
        .O(\u2/u3/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__281
       (.I0(\u2/u3/X [35]),
        .I1(\u2/u3/X [34]),
        .I2(\u2/u3/X [33]),
        .I3(\u2/u3/X [32]),
        .I4(\u2/u3/X [36]),
        .I5(\u2/u3/X [31]),
        .O(\u2/out3 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__281_i_1
       (.I0(\u2/R2 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [15]),
        .I3(\u2/uk/K_r2 [52]),
        .O(\u2/u3/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__281_i_2
       (.I0(\u2/R2 [23]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [44]),
        .I3(\u2/uk/K_r2 [22]),
        .O(\u2/u3/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__281_i_3
       (.I0(\u2/R2 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [0]),
        .I3(\u2/uk/K_r2 [9]),
        .O(\u2/u3/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__281_i_4
       (.I0(\u2/R2 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [9]),
        .I3(\u2/uk/K_r2 [42]),
        .O(\u2/u3/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__281_i_5
       (.I0(\u2/R2 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [38]),
        .I3(\u2/uk/K_r2 [43]),
        .O(\u2/u3/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__281_i_6
       (.I0(\u2/R2 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [49]),
        .I3(\u2/uk/K_r2 [31]),
        .O(\u2/u3/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__282
       (.I0(\u2/u3/X [11]),
        .I1(\u2/u3/X [10]),
        .I2(\u2/u3/X [9]),
        .I3(\u2/u3/X [8]),
        .I4(\u2/u3/X [12]),
        .I5(\u2/u3/X [7]),
        .O(\u2/out3 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__282_i_1
       (.I0(\u2/R2 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [17]),
        .I3(\u2/uk/K_r2 [54]),
        .O(\u2/u3/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__282_i_2
       (.I0(\u2/R2 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [26]),
        .I3(\u2/uk/K_r2 [6]),
        .O(\u2/u3/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__282_i_3
       (.I0(\u2/R2 [6]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [32]),
        .I3(\u2/uk/K_r2 [12]),
        .O(\u2/u3/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__282_i_4
       (.I0(\u2/R2 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [41]),
        .I3(\u2/uk/K_r2 [46]),
        .O(\u2/u3/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__282_i_5
       (.I0(\u2/R2 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [54]),
        .I3(\u2/uk/K_r2 [34]),
        .O(\u2/u3/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__282_i_6
       (.I0(\u2/R2 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [5]),
        .I3(\u2/uk/K_r2 [10]),
        .O(\u2/u3/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__283
       (.I0(\u2/u3/X [47]),
        .I1(\u2/u3/X [46]),
        .I2(\u2/u3/X [45]),
        .I3(\u2/u3/X [44]),
        .I4(\u2/u3/X [48]),
        .I5(\u2/u3/X [43]),
        .O(\u2/out3 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__283_i_1
       (.I0(\u2/R2 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [42]),
        .I3(\u2/uk/K_r2 [51]),
        .O(\u2/u3/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__283_i_2
       (.I0(\u2/R2 [31]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [36]),
        .I3(\u2/uk/K_r2 [14]),
        .O(\u2/u3/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__283_i_3
       (.I0(\u2/R2 [30]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [52]),
        .I3(\u2/uk/K_r2 [2]),
        .O(\u2/u3/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__283_i_4
       (.I0(\u2/R2 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [23]),
        .I3(\u2/uk/K_r2 [1]),
        .O(\u2/u3/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__283_i_5
       (.I0(\u2/R2 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [8]),
        .I3(\u2/uk/K_r2 [45]),
        .O(\u2/u3/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__283_i_6
       (.I0(\u2/R2 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [51]),
        .I3(\u2/uk/K_r2 [29]),
        .O(\u2/u3/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__284
       (.I0(\u2/u3/X [23]),
        .I1(\u2/u3/X [22]),
        .I2(\u2/u3/X [21]),
        .I3(\u2/u3/X [20]),
        .I4(\u2/u3/X [24]),
        .I5(\u2/u3/X [19]),
        .O(\u2/out3 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__284_i_1
       (.I0(\u2/R2 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [18]),
        .I3(\u2/uk/K_r2 [55]),
        .O(\u2/u3/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__284_i_2
       (.I0(\u2/R2 [15]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [10]),
        .I3(\u2/uk/K_r2 [47]),
        .O(\u2/u3/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__284_i_3
       (.I0(\u2/R2 [14]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [34]),
        .I3(\u2/uk/K_r2 [39]),
        .O(\u2/u3/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__284_i_4
       (.I0(\u2/R2 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [33]),
        .I3(\u2/uk/K_r2 [13]),
        .O(\u2/u3/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__284_i_5
       (.I0(\u2/R2 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [55]),
        .I3(\u2/uk/K_r2 [3]),
        .O(\u2/u3/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__284_i_6
       (.I0(\u2/R2 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [39]),
        .I3(\u2/uk/K_r2 [19]),
        .O(\u2/u3/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__285
       (.I0(\u2/u3/X [29]),
        .I1(\u2/u3/X [28]),
        .I2(\u2/u3/X [27]),
        .I3(\u2/u3/X [26]),
        .I4(\u2/u3/X [30]),
        .I5(\u2/u3/X [25]),
        .O(\u2/out3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__285_i_1
       (.I0(\u2/R2 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [31]),
        .I3(\u2/uk/K_r2 [36]),
        .O(\u2/u3/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__285_i_2
       (.I0(\u2/R2 [19]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [43]),
        .I3(\u2/uk/K_r2 [21]),
        .O(\u2/u3/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__285_i_3
       (.I0(\u2/R2 [18]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [1]),
        .I3(\u2/uk/K_r2 [38]),
        .O(\u2/u3/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__285_i_4
       (.I0(\u2/R2 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [7]),
        .I3(\u2/uk/K_r2 [16]),
        .O(\u2/u3/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__285_i_5
       (.I0(\u2/R2 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [28]),
        .I3(\u2/uk/K_r2 [37]),
        .O(\u2/u3/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__285_i_6
       (.I0(\u2/R2 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [16]),
        .I3(\u2/uk/K_r2 [49]),
        .O(\u2/u3/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__286
       (.I0(\u2/u3/X [5]),
        .I1(\u2/u3/X [4]),
        .I2(\u2/u3/X [3]),
        .I3(\u2/u3/X [2]),
        .I4(\u2/u3/X [6]),
        .I5(\u2/u3/X [1]),
        .O(\u2/out3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__286_i_1
       (.I0(\u2/R2 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [48]),
        .I3(\u2/uk/K_r2 [53]),
        .O(\u2/u3/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__286_i_2
       (.I0(\u2/R2 [3]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [13]),
        .I3(\u2/uk/K_r2 [18]),
        .O(\u2/u3/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__286_i_3
       (.I0(\u2/R2 [2]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [4]),
        .I3(\u2/uk/K_r2 [41]),
        .O(\u2/u3/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__286_i_4
       (.I0(\u2/R2 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [46]),
        .I3(\u2/uk/K_r2 [26]),
        .O(\u2/u3/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__286_i_5
       (.I0(\u2/R2 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [19]),
        .I3(\u2/uk/K_r2 [24]),
        .O(\u2/u3/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__286_i_6
       (.I0(\u2/R2 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r2 [25]),
        .I3(\u2/uk/K_r2 [5]),
        .O(\u2/u3/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__287
       (.I0(\u2/u4/X [41]),
        .I1(\u2/u4/X [40]),
        .I2(\u2/u4/X [39]),
        .I3(\u2/u4/X [38]),
        .I4(\u2/u4/X [42]),
        .I5(\u2/u4/X [37]),
        .O(\u2/out4 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__287_i_1
       (.I0(\u2/R3 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [36]),
        .I3(\u2/uk/K_r3 [45]),
        .O(\u2/u4/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__287_i_2
       (.I0(\u2/R3 [27]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [49]),
        .I3(\u2/uk/K_r3 [30]),
        .O(\u2/u4/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__287_i_3
       (.I0(\u2/R3 [26]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [16]),
        .I3(\u2/uk/K_r3 [21]),
        .O(\u2/u4/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__287_i_4
       (.I0(\u2/R3 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [0]),
        .I3(\u2/uk/K_r3 [36]),
        .O(\u2/u4/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__287_i_5
       (.I0(\u2/R3 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [28]),
        .I3(\u2/uk/K_r3 [9]),
        .O(\u2/u4/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__287_i_6
       (.I0(\u2/R3 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [51]),
        .I3(\u2/uk/K_r3 [1]),
        .O(\u2/u4/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__288
       (.I0(\u2/u4/X [17]),
        .I1(\u2/u4/X [16]),
        .I2(\u2/u4/X [15]),
        .I3(\u2/u4/X [14]),
        .I4(\u2/u4/X [18]),
        .I5(\u2/u4/X [13]),
        .O(\u2/out4 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__288_i_1
       (.I0(\u2/R3 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [41]),
        .I3(\u2/uk/K_r3 [18]),
        .O(\u2/u4/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__288_i_2
       (.I0(\u2/R3 [11]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [26]),
        .I3(\u2/uk/K_r3 [3]),
        .O(\u2/u4/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__288_i_3
       (.I0(\u2/R3 [10]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [25]),
        .I3(\u2/uk/K_r3 [34]),
        .O(\u2/u4/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__288_i_4
       (.I0(\u2/R3 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [17]),
        .I3(\u2/uk/K_r3 [26]),
        .O(\u2/u4/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__288_i_5
       (.I0(\u2/R3 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [54]),
        .I3(\u2/uk/K_r3 [6]),
        .O(\u2/u4/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__288_i_6
       (.I0(\u2/R3 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [20]),
        .I3(\u2/uk/K_r3 [54]),
        .O(\u2/u4/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__289
       (.I0(\u2/u4/X [35]),
        .I1(\u2/u4/X [34]),
        .I2(\u2/u4/X [33]),
        .I3(\u2/u4/X [32]),
        .I4(\u2/u4/X [36]),
        .I5(\u2/u4/X [31]),
        .O(\u2/out4 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__289_i_1
       (.I0(\u2/R3 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [29]),
        .I3(\u2/uk/K_r3 [38]),
        .O(\u2/u4/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__289_i_2
       (.I0(\u2/R3 [23]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [31]),
        .I3(\u2/uk/K_r3 [8]),
        .O(\u2/u4/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__289_i_3
       (.I0(\u2/R3 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [14]),
        .I3(\u2/uk/K_r3 [50]),
        .O(\u2/u4/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__289_i_4
       (.I0(\u2/R3 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [23]),
        .I3(\u2/uk/K_r3 [28]),
        .O(\u2/u4/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__289_i_5
       (.I0(\u2/R3 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [52]),
        .I3(\u2/uk/K_r3 [29]),
        .O(\u2/u4/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__289_i_6
       (.I0(\u2/R3 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [8]),
        .I3(\u2/uk/K_r3 [44]),
        .O(\u2/u4/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__28_i_1
       (.I0(\u0/R2 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [18]),
        .I3(\u0/uk/K_r2 [55]),
        .O(\u0/u3/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__28_i_2
       (.I0(\u0/R2 [15]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [10]),
        .I3(\u0/uk/K_r2 [47]),
        .O(\u0/u3/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__28_i_3
       (.I0(\u0/R2 [14]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [34]),
        .I3(\u0/uk/K_r2 [39]),
        .O(\u0/u3/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__28_i_4
       (.I0(\u0/R2 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [33]),
        .I3(\u0/uk/K_r2 [13]),
        .O(\u0/u3/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__28_i_5
       (.I0(\u0/R2 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [55]),
        .I3(\u0/uk/K_r2 [3]),
        .O(\u0/u3/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__28_i_6
       (.I0(\u0/R2 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [39]),
        .I3(\u0/uk/K_r2 [19]),
        .O(\u0/u3/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__29
       (.I0(\u0/u3/X [29]),
        .I1(\u0/u3/X [28]),
        .I2(\u0/u3/X [27]),
        .I3(\u0/u3/X [26]),
        .I4(\u0/u3/X [30]),
        .I5(\u0/u3/X [25]),
        .O(\u0/out3 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__290
       (.I0(\u2/u4/X [11]),
        .I1(\u2/u4/X [10]),
        .I2(\u2/u4/X [9]),
        .I3(\u2/u4/X [8]),
        .I4(\u2/u4/X [12]),
        .I5(\u2/u4/X [7]),
        .O(\u2/out4 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__290_i_1
       (.I0(\u2/R3 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [6]),
        .I3(\u2/uk/K_r3 [40]),
        .O(\u2/u4/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__290_i_2
       (.I0(\u2/R3 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [40]),
        .I3(\u2/uk/K_r3 [17]),
        .O(\u2/u4/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__290_i_3
       (.I0(\u2/R3 [6]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [46]),
        .I3(\u2/uk/K_r3 [55]),
        .O(\u2/u4/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__290_i_4
       (.I0(\u2/R3 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [55]),
        .I3(\u2/uk/K_r3 [32]),
        .O(\u2/u4/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__290_i_5
       (.I0(\u2/R3 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [11]),
        .I3(\u2/uk/K_r3 [20]),
        .O(\u2/u4/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__290_i_6
       (.I0(\u2/R3 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [19]),
        .I3(\u2/uk/K_r3 [53]),
        .O(\u2/u4/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__291
       (.I0(\u2/u4/X [47]),
        .I1(\u2/u4/X [46]),
        .I2(\u2/u4/X [45]),
        .I3(\u2/u4/X [44]),
        .I4(\u2/u4/X [48]),
        .I5(\u2/u4/X [43]),
        .O(\u2/out4 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__291_i_1
       (.I0(\u2/R3 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [1]),
        .I3(\u2/uk/K_r3 [37]),
        .O(\u2/u4/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__291_i_2
       (.I0(\u2/R3 [31]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [50]),
        .I3(\u2/uk/K_r3 [0]),
        .O(\u2/u4/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__291_i_3
       (.I0(\u2/R3 [30]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [7]),
        .I3(\u2/uk/K_r3 [43]),
        .O(\u2/u4/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__291_i_4
       (.I0(\u2/R3 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [37]),
        .I3(\u2/uk/K_r3 [42]),
        .O(\u2/u4/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__291_i_5
       (.I0(\u2/R3 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [22]),
        .I3(\u2/uk/K_r3 [31]),
        .O(\u2/u4/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__291_i_6
       (.I0(\u2/R3 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [38]),
        .I3(\u2/uk/K_r3 [15]),
        .O(\u2/u4/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__292
       (.I0(\u2/u4/X [23]),
        .I1(\u2/u4/X [22]),
        .I2(\u2/u4/X [21]),
        .I3(\u2/u4/X [20]),
        .I4(\u2/u4/X [24]),
        .I5(\u2/u4/X [19]),
        .O(\u2/out4 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__292_i_1
       (.I0(\u2/R3 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [32]),
        .I3(\u2/uk/K_r3 [41]),
        .O(\u2/u4/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__292_i_2
       (.I0(\u2/R3 [15]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [24]),
        .I3(\u2/uk/K_r3 [33]),
        .O(\u2/u4/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__292_i_3
       (.I0(\u2/R3 [14]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [48]),
        .I3(\u2/uk/K_r3 [25]),
        .O(\u2/u4/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__292_i_4
       (.I0(\u2/R3 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [47]),
        .I3(\u2/uk/K_r3 [24]),
        .O(\u2/u4/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__292_i_5
       (.I0(\u2/R3 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [12]),
        .I3(\u2/uk/K_r3 [46]),
        .O(\u2/u4/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__292_i_6
       (.I0(\u2/R3 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [53]),
        .I3(\u2/uk/K_r3 [5]),
        .O(\u2/u4/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__293
       (.I0(\u2/u4/X [29]),
        .I1(\u2/u4/X [28]),
        .I2(\u2/u4/X [27]),
        .I3(\u2/u4/X [26]),
        .I4(\u2/u4/X [30]),
        .I5(\u2/u4/X [25]),
        .O(\u2/out4 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__293_i_1
       (.I0(\u2/R3 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [45]),
        .I3(\u2/uk/K_r3 [22]),
        .O(\u2/u4/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__293_i_2
       (.I0(\u2/R3 [19]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [2]),
        .I3(\u2/uk/K_r3 [7]),
        .O(\u2/u4/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__293_i_3
       (.I0(\u2/R3 [18]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [15]),
        .I3(\u2/uk/K_r3 [51]),
        .O(\u2/u4/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__293_i_4
       (.I0(\u2/R3 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [21]),
        .I3(\u2/uk/K_r3 [2]),
        .O(\u2/u4/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__293_i_5
       (.I0(\u2/R3 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [42]),
        .I3(\u2/uk/K_r3 [23]),
        .O(\u2/u4/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__293_i_6
       (.I0(\u2/R3 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [30]),
        .I3(\u2/uk/K_r3 [35]),
        .O(\u2/u4/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__294
       (.I0(\u2/u4/X [5]),
        .I1(\u2/u4/X [4]),
        .I2(\u2/u4/X [3]),
        .I3(\u2/u4/X [2]),
        .I4(\u2/u4/X [6]),
        .I5(\u2/u4/X [1]),
        .O(\u2/out4 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__294_i_1
       (.I0(\u2/R3 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [5]),
        .I3(\u2/uk/K_r3 [39]),
        .O(\u2/u4/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__294_i_2
       (.I0(\u2/R3 [3]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [27]),
        .I3(\u2/uk/K_r3 [4]),
        .O(\u2/u4/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__294_i_3
       (.I0(\u2/R3 [2]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [18]),
        .I3(\u2/uk/K_r3 [27]),
        .O(\u2/u4/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__294_i_4
       (.I0(\u2/R3 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [3]),
        .I3(\u2/uk/K_r3 [12]),
        .O(\u2/u4/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__294_i_5
       (.I0(\u2/R3 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [33]),
        .I3(\u2/uk/K_r3 [10]),
        .O(\u2/u4/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__294_i_6
       (.I0(\u2/R3 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r3 [39]),
        .I3(\u2/uk/K_r3 [48]),
        .O(\u2/u4/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__295
       (.I0(\u2/u5/X [41]),
        .I1(\u2/u5/X [40]),
        .I2(\u2/u5/X [39]),
        .I3(\u2/u5/X [38]),
        .I4(\u2/u5/X [42]),
        .I5(\u2/u5/X [37]),
        .O(\u2/out5 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__295_i_1
       (.I0(\u2/R4 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[50] ),
        .I3(\u2/uk/K_r4_reg_n_0_[31] ),
        .O(\u2/u5/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__295_i_2
       (.I0(\u2/R4 [27]),
        .I1(decrypt),
        .I2(\u2/uk/p_42_in ),
        .I3(\u2/uk/K_r4_reg_n_0_[16] ),
        .O(\u2/u5/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__295_i_3
       (.I0(\u2/R4 [26]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[30] ),
        .I3(\u2/uk/K_r4_reg_n_0_[7] ),
        .O(\u2/u5/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__295_i_4
       (.I0(\u2/R4 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[14] ),
        .I3(\u2/uk/K_r4_reg_n_0_[22] ),
        .O(\u2/u5/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__295_i_5
       (.I0(\u2/R4 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[42] ),
        .I3(\u2/uk/K_r4_reg_n_0_[50] ),
        .O(\u2/u5/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__295_i_6
       (.I0(\u2/R4 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[38] ),
        .I3(\u2/uk/K_r4_reg_n_0_[42] ),
        .O(\u2/u5/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__296
       (.I0(\u2/u5/X [17]),
        .I1(\u2/u5/X [16]),
        .I2(\u2/u5/X [15]),
        .I3(\u2/u5/X [14]),
        .I4(\u2/u5/X [18]),
        .I5(\u2/u5/X [13]),
        .O(\u2/out5 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__296_i_1
       (.I0(\u2/R4 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[55] ),
        .I3(\u2/uk/K_r4_reg_n_0_[4] ),
        .O(\u2/u5/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__296_i_2
       (.I0(\u2/R4 [11]),
        .I1(decrypt),
        .I2(\u2/uk/p_49_in ),
        .I3(\u2/uk/p_47_in ),
        .O(\u2/u5/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__296_i_3
       (.I0(\u2/R4 [10]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[39] ),
        .I3(\u2/uk/K_r4_reg_n_0_[20] ),
        .O(\u2/u5/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__296_i_4
       (.I0(\u2/R4 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[6] ),
        .I3(\u2/uk/K_r4_reg_n_0_[12] ),
        .O(\u2/u5/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__296_i_5
       (.I0(\u2/R4 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[11] ),
        .I3(\u2/uk/K_r4_reg_n_0_[17] ),
        .O(\u2/u5/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__296_i_6
       (.I0(\u2/R4 [8]),
        .I1(decrypt),
        .I2(\u2/uk/p_50_in ),
        .I3(\u2/uk/p_49_in ),
        .O(\u2/u5/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__297
       (.I0(\u2/u5/X [35]),
        .I1(\u2/u5/X [34]),
        .I2(\u2/u5/X [33]),
        .I3(\u2/u5/X [32]),
        .I4(\u2/u5/X [36]),
        .I5(\u2/u5/X [31]),
        .O(\u2/out5 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__297_i_1
       (.I0(\u2/R4 [24]),
        .I1(decrypt),
        .I2(\u2/uk/p_44_in ),
        .I3(\u2/uk/K_r4_reg_n_0_[51] ),
        .O(\u2/u5/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__297_i_2
       (.I0(\u2/R4 [23]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[45] ),
        .I3(\u2/uk/K_r4_reg_n_0_[49] ),
        .O(\u2/u5/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__297_i_3
       (.I0(\u2/R4 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[28] ),
        .I3(\u2/uk/K_r4_reg_n_0_[36] ),
        .O(\u2/u5/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__297_i_4
       (.I0(\u2/R4 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[37] ),
        .I3(\u2/uk/K_r4_reg_n_0_[14] ),
        .O(\u2/u5/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__297_i_5
       (.I0(\u2/R4 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[7] ),
        .I3(\u2/uk/K_r4_reg_n_0_[15] ),
        .O(\u2/u5/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__297_i_6
       (.I0(\u2/R4 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[22] ),
        .I3(\u2/uk/K_r4_reg_n_0_[30] ),
        .O(\u2/u5/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__298
       (.I0(\u2/u5/X [11]),
        .I1(\u2/u5/X [10]),
        .I2(\u2/u5/X [9]),
        .I3(\u2/u5/X [8]),
        .I4(\u2/u5/X [12]),
        .I5(\u2/u5/X [7]),
        .O(\u2/out5 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__298_i_1
       (.I0(\u2/R4 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[20] ),
        .I3(\u2/uk/K_r4_reg_n_0_[26] ),
        .O(\u2/u5/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__298_i_2
       (.I0(\u2/R4 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[54] ),
        .I3(\u2/uk/K_r4_reg_n_0_[3] ),
        .O(\u2/u5/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__298_i_3
       (.I0(\u2/R4 [6]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[3] ),
        .I3(\u2/uk/K_r4_reg_n_0_[41] ),
        .O(\u2/u5/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__298_i_4
       (.I0(\u2/R4 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[12] ),
        .I3(\u2/uk/K_r4_reg_n_0_[18] ),
        .O(\u2/u5/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__298_i_5
       (.I0(\u2/R4 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[25] ),
        .I3(\u2/uk/K_r4_reg_n_0_[6] ),
        .O(\u2/u5/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__298_i_6
       (.I0(\u2/R4 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[33] ),
        .I3(\u2/uk/K_r4_reg_n_0_[39] ),
        .O(\u2/u5/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__299
       (.I0(\u2/u5/X [47]),
        .I1(\u2/u5/X [46]),
        .I2(\u2/u5/X [45]),
        .I3(\u2/u5/X [44]),
        .I4(\u2/u5/X [48]),
        .I5(\u2/u5/X [43]),
        .O(\u2/out5 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__299_i_1
       (.I0(\u2/R4 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[15] ),
        .I3(\u2/uk/K_r4_reg_n_0_[23] ),
        .O(\u2/u5/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__299_i_2
       (.I0(\u2/R4 [31]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[9] ),
        .I3(\u2/uk/K_r4_reg_n_0_[45] ),
        .O(\u2/u5/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__299_i_3
       (.I0(\u2/R4 [30]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[21] ),
        .I3(\u2/uk/K_r4_reg_n_0_[29] ),
        .O(\u2/u5/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__299_i_4
       (.I0(\u2/R4 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[51] ),
        .I3(\u2/uk/K_r4_reg_n_0_[28] ),
        .O(\u2/u5/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__299_i_5
       (.I0(\u2/R4 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[36] ),
        .I3(\u2/uk/K_r4_reg_n_0_[44] ),
        .O(\u2/u5/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__299_i_6
       (.I0(\u2/R4 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[52] ),
        .I3(\u2/uk/K_r4_reg_n_0_[1] ),
        .O(\u2/u5/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__29_i_1
       (.I0(\u0/R2 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [31]),
        .I3(\u0/uk/K_r2 [36]),
        .O(\u0/u3/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__29_i_2
       (.I0(\u0/R2 [19]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [43]),
        .I3(\u0/uk/K_r2 [21]),
        .O(\u0/u3/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__29_i_3
       (.I0(\u0/R2 [18]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [1]),
        .I3(\u0/uk/K_r2 [38]),
        .O(\u0/u3/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__29_i_4
       (.I0(\u0/R2 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [7]),
        .I3(\u0/uk/K_r2 [16]),
        .O(\u0/u3/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__29_i_5
       (.I0(\u0/R2 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [28]),
        .I3(\u0/uk/K_r2 [37]),
        .O(\u0/u3/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__29_i_6
       (.I0(\u0/R2 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [16]),
        .I3(\u0/uk/K_r2 [49]),
        .O(\u0/u3/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__2_i_1
       (.I0(\u0/IP [40]),
        .I1(decrypt),
        .I2(\u0/key_r [39]),
        .I3(\u0/key_r [32]),
        .O(\u0/u0/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__2_i_2
       (.I0(\u0/IP [39]),
        .I1(decrypt),
        .I2(\u0/key_r [48]),
        .I3(\u0/key_r [41]),
        .O(\u0/u0/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__2_i_3
       (.I0(\u0/IP [38]),
        .I1(decrypt),
        .I2(\u0/key_r [54]),
        .I3(\u0/key_r [47]),
        .O(\u0/u0/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__2_i_4
       (.I0(\u0/IP [37]),
        .I1(decrypt),
        .I2(\u0/key_r [6]),
        .I3(\u0/key_r [24]),
        .O(\u0/u0/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__2_i_5
       (.I0(\u0/IP [41]),
        .I1(decrypt),
        .I2(\u0/key_r [19]),
        .I3(\u0/key_r [12]),
        .O(\u0/u0/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__2_i_6
       (.I0(\u0/IP [36]),
        .I1(decrypt),
        .I2(\u0/key_r [27]),
        .I3(\u0/key_r [20]),
        .O(\u0/u0/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__3
       (.I0(\u0/u0/X [47]),
        .I1(\u0/u0/X [46]),
        .I2(\u0/u0/X [45]),
        .I3(\u0/u0/X [44]),
        .I4(\u0/u0/X [48]),
        .I5(\u0/u0/X [43]),
        .O(\u0/out0 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__30
       (.I0(\u0/u3/X [5]),
        .I1(\u0/u3/X [4]),
        .I2(\u0/u3/X [3]),
        .I3(\u0/u3/X [2]),
        .I4(\u0/u3/X [6]),
        .I5(\u0/u3/X [1]),
        .O(\u0/out3 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__300
       (.I0(\u2/u5/X [23]),
        .I1(\u2/u5/X [22]),
        .I2(\u2/u5/X [21]),
        .I3(\u2/u5/X [20]),
        .I4(\u2/u5/X [24]),
        .I5(\u2/u5/X [19]),
        .O(\u2/out5 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__300_i_1
       (.I0(\u2/R4 [16]),
        .I1(decrypt),
        .I2(\u2/uk/p_47_in ),
        .I3(\u2/uk/K_r4_reg_n_0_[27] ),
        .O(\u2/u5/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__300_i_2
       (.I0(\u2/R4 [15]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[13] ),
        .I3(\u2/uk/K_r4_reg_n_0_[19] ),
        .O(\u2/u5/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__300_i_3
       (.I0(\u2/R4 [14]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[5] ),
        .I3(\u2/uk/K_r4_reg_n_0_[11] ),
        .O(\u2/u5/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__300_i_4
       (.I0(\u2/R4 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[4] ),
        .I3(\u2/uk/K_r4_reg_n_0_[10] ),
        .O(\u2/u5/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__300_i_5
       (.I0(\u2/R4 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[26] ),
        .I3(\u2/uk/K_r4_reg_n_0_[32] ),
        .O(\u2/u5/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__300_i_6
       (.I0(\u2/R4 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[10] ),
        .I3(\u2/uk/K_r4_reg_n_0_[48] ),
        .O(\u2/u5/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__301
       (.I0(\u2/u5/X [29]),
        .I1(\u2/u5/X [28]),
        .I2(\u2/u5/X [27]),
        .I3(\u2/u5/X [26]),
        .I4(\u2/u5/X [30]),
        .I5(\u2/u5/X [25]),
        .O(\u2/out5 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__301_i_1
       (.I0(\u2/R4 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_ ),
        .I3(\u2/uk/p_42_in ),
        .O(\u2/u5/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__301_i_2
       (.I0(\u2/R4 [19]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[16] ),
        .I3(\u2/uk/K_r4_reg_n_0_[52] ),
        .O(\u2/u5/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__301_i_3
       (.I0(\u2/R4 [18]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[29] ),
        .I3(\u2/uk/K_r4_reg_n_0_[37] ),
        .O(\u2/u5/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__301_i_4
       (.I0(\u2/R4 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[35] ),
        .I3(\u2/uk/p_44_in ),
        .O(\u2/u5/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__301_i_5
       (.I0(\u2/R4 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[1] ),
        .I3(\u2/uk/K_r4_reg_n_0_[9] ),
        .O(\u2/u5/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__301_i_6
       (.I0(\u2/R4 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[44] ),
        .I3(\u2/uk/K_r4_reg_n_0_[21] ),
        .O(\u2/u5/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__302
       (.I0(\u2/u5/X [5]),
        .I1(\u2/u5/X [4]),
        .I2(\u2/u5/X [3]),
        .I3(\u2/u5/X [2]),
        .I4(\u2/u5/X [6]),
        .I5(\u2/u5/X [1]),
        .O(\u2/out5 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__302_i_1
       (.I0(\u2/R4 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[19] ),
        .I3(\u2/uk/K_r4_reg_n_0_[25] ),
        .O(\u2/u5/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__302_i_2
       (.I0(\u2/R4 [3]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[41] ),
        .I3(\u2/uk/K_r4_reg_n_0_[47] ),
        .O(\u2/u5/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__302_i_3
       (.I0(\u2/R4 [2]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[32] ),
        .I3(\u2/uk/K_r4_reg_n_0_[13] ),
        .O(\u2/u5/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__302_i_4
       (.I0(\u2/R4 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[17] ),
        .I3(\u2/uk/K_r4_reg_n_0_[55] ),
        .O(\u2/u5/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__302_i_5
       (.I0(\u2/R4 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r4_reg_n_0_[47] ),
        .I3(\u2/uk/p_51_in ),
        .O(\u2/u5/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__302_i_6
       (.I0(\u2/R4 [32]),
        .I1(decrypt),
        .I2(\u2/uk/p_51_in ),
        .I3(\u2/uk/p_50_in ),
        .O(\u2/u5/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__303
       (.I0(\u2/u6/X [41]),
        .I1(\u2/u6/X [40]),
        .I2(\u2/u6/X [39]),
        .I3(\u2/u6/X [38]),
        .I4(\u2/u6/X [42]),
        .I5(\u2/u6/X [37]),
        .O(\u2/out6 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__303_i_1
       (.I0(\u2/R5 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [9]),
        .I3(\u2/uk/K_r5 [44]),
        .O(\u2/u6/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__303_i_2
       (.I0(\u2/R5 [27]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [22]),
        .I3(\u2/uk/K_r5 [2]),
        .O(\u2/u6/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__303_i_3
       (.I0(\u2/R5 [26]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [44]),
        .I3(\u2/uk/K_r5 [52]),
        .O(\u2/u6/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__303_i_4
       (.I0(\u2/R5 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [28]),
        .I3(\u2/uk/K_r5 [8]),
        .O(\u2/u6/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__303_i_5
       (.I0(\u2/R5 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [1]),
        .I3(\u2/uk/K_r5 [36]),
        .O(\u2/u6/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__303_i_6
       (.I0(\u2/R5 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [52]),
        .I3(\u2/uk/K_r5 [28]),
        .O(\u2/u6/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__304
       (.I0(\u2/u6/X [17]),
        .I1(\u2/u6/X [16]),
        .I2(\u2/u6/X [15]),
        .I3(\u2/u6/X [14]),
        .I4(\u2/u6/X [18]),
        .I5(\u2/u6/X [13]),
        .O(\u2/out6 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__304_i_1
       (.I0(\u2/R5 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [12]),
        .I3(\u2/uk/K_r5 [47]),
        .O(\u2/u6/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__304_i_2
       (.I0(\u2/R5 [11]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [54]),
        .I3(\u2/uk/K_r5 [32]),
        .O(\u2/u6/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__304_i_3
       (.I0(\u2/R5 [10]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [53]),
        .I3(\u2/uk/K_r5 [6]),
        .O(\u2/u6/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__304_i_4
       (.I0(\u2/R5 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [20]),
        .I3(\u2/uk/K_r5 [55]),
        .O(\u2/u6/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__304_i_5
       (.I0(\u2/R5 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [25]),
        .I3(\u2/uk/K_r5 [3]),
        .O(\u2/u6/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__304_i_6
       (.I0(\u2/R5 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [48]),
        .I3(\u2/uk/K_r5 [26]),
        .O(\u2/u6/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__305
       (.I0(\u2/u6/X [35]),
        .I1(\u2/u6/X [34]),
        .I2(\u2/u6/X [33]),
        .I3(\u2/u6/X [32]),
        .I4(\u2/u6/X [36]),
        .I5(\u2/u6/X [31]),
        .O(\u2/out6 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__305_i_1
       (.I0(\u2/R5 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [2]),
        .I3(\u2/uk/K_r5 [37]),
        .O(\u2/u6/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__305_i_2
       (.I0(\u2/R5 [23]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [0]),
        .I3(\u2/uk/K_r5 [35]),
        .O(\u2/u6/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__305_i_3
       (.I0(\u2/R5 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [42]),
        .I3(\u2/uk/K_r5 [22]),
        .O(\u2/u6/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__305_i_4
       (.I0(\u2/R5 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [51]),
        .I3(\u2/uk/K_r5 [0]),
        .O(\u2/u6/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__305_i_5
       (.I0(\u2/R5 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [21]),
        .I3(\u2/uk/K_r5 [1]),
        .O(\u2/u6/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__305_i_6
       (.I0(\u2/R5 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [36]),
        .I3(\u2/uk/K_r5 [16]),
        .O(\u2/u6/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__306
       (.I0(\u2/u6/X [11]),
        .I1(\u2/u6/X [10]),
        .I2(\u2/u6/X [9]),
        .I3(\u2/u6/X [8]),
        .I4(\u2/u6/X [12]),
        .I5(\u2/u6/X [7]),
        .O(\u2/out6 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__306_i_1
       (.I0(\u2/R5 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [34]),
        .I3(\u2/uk/K_r5 [12]),
        .O(\u2/u6/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__306_i_2
       (.I0(\u2/R5 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [11]),
        .I3(\u2/uk/K_r5 [46]),
        .O(\u2/u6/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__306_i_3
       (.I0(\u2/R5 [6]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [17]),
        .I3(\u2/uk/K_r5 [27]),
        .O(\u2/u6/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__306_i_4
       (.I0(\u2/R5 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [26]),
        .I3(\u2/uk/K_r5 [4]),
        .O(\u2/u6/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__306_i_5
       (.I0(\u2/R5 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [39]),
        .I3(\u2/uk/K_r5 [17]),
        .O(\u2/u6/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__306_i_6
       (.I0(\u2/R5 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [47]),
        .I3(\u2/uk/K_r5 [25]),
        .O(\u2/u6/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__307
       (.I0(\u2/u6/X [47]),
        .I1(\u2/u6/X [46]),
        .I2(\u2/u6/X [45]),
        .I3(\u2/u6/X [44]),
        .I4(\u2/u6/X [48]),
        .I5(\u2/u6/X [43]),
        .O(\u2/out6 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__307_i_1
       (.I0(\u2/R5 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [29]),
        .I3(\u2/uk/K_r5 [9]),
        .O(\u2/u6/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__307_i_2
       (.I0(\u2/R5 [31]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [23]),
        .I3(\u2/uk/K_r5 [31]),
        .O(\u2/u6/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__307_i_3
       (.I0(\u2/R5 [30]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [35]),
        .I3(\u2/uk/K_r5 [15]),
        .O(\u2/u6/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__307_i_4
       (.I0(\u2/R5 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [38]),
        .I3(\u2/uk/K_r5 [14]),
        .O(\u2/u6/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__307_i_5
       (.I0(\u2/R5 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [50]),
        .I3(\u2/uk/K_r5 [30]),
        .O(\u2/u6/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__307_i_6
       (.I0(\u2/R5 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [7]),
        .I3(\u2/uk/K_r5 [42]),
        .O(\u2/u6/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__308
       (.I0(\u2/u6/X [23]),
        .I1(\u2/u6/X [22]),
        .I2(\u2/u6/X [21]),
        .I3(\u2/u6/X [20]),
        .I4(\u2/u6/X [24]),
        .I5(\u2/u6/X [19]),
        .O(\u2/out6 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__308_i_1
       (.I0(\u2/R5 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [3]),
        .I3(\u2/uk/K_r5 [13]),
        .O(\u2/u6/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__308_i_2
       (.I0(\u2/R5 [15]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [27]),
        .I3(\u2/uk/K_r5 [5]),
        .O(\u2/u6/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__308_i_3
       (.I0(\u2/R5 [14]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [19]),
        .I3(\u2/uk/K_r5 [54]),
        .O(\u2/u6/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__308_i_4
       (.I0(\u2/R5 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [18]),
        .I3(\u2/uk/K_r5 [53]),
        .O(\u2/u6/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__308_i_5
       (.I0(\u2/R5 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [40]),
        .I3(\u2/uk/K_r5 [18]),
        .O(\u2/u6/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__308_i_6
       (.I0(\u2/R5 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [24]),
        .I3(\u2/uk/K_r5 [34]),
        .O(\u2/u6/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__309
       (.I0(\u2/u6/X [29]),
        .I1(\u2/u6/X [28]),
        .I2(\u2/u6/X [27]),
        .I3(\u2/u6/X [26]),
        .I4(\u2/u6/X [30]),
        .I5(\u2/u6/X [25]),
        .O(\u2/out6 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__309_i_1
       (.I0(\u2/R5 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [14]),
        .I3(\u2/uk/K_r5 [49]),
        .O(\u2/u6/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__309_i_2
       (.I0(\u2/R5 [19]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [30]),
        .I3(\u2/uk/K_r5 [38]),
        .O(\u2/u6/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__309_i_3
       (.I0(\u2/R5 [18]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [43]),
        .I3(\u2/uk/K_r5 [23]),
        .O(\u2/u6/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__309_i_4
       (.I0(\u2/R5 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [49]),
        .I3(\u2/uk/K_r5 [29]),
        .O(\u2/u6/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__309_i_5
       (.I0(\u2/R5 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [15]),
        .I3(\u2/uk/K_r5 [50]),
        .O(\u2/u6/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__309_i_6
       (.I0(\u2/R5 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [31]),
        .I3(\u2/uk/K_r5 [7]),
        .O(\u2/u6/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__30_i_1
       (.I0(\u0/R2 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [48]),
        .I3(\u0/uk/K_r2 [53]),
        .O(\u0/u3/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__30_i_2
       (.I0(\u0/R2 [3]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [13]),
        .I3(\u0/uk/K_r2 [18]),
        .O(\u0/u3/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__30_i_3
       (.I0(\u0/R2 [2]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [4]),
        .I3(\u0/uk/K_r2 [41]),
        .O(\u0/u3/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__30_i_4
       (.I0(\u0/R2 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [46]),
        .I3(\u0/uk/K_r2 [26]),
        .O(\u0/u3/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__30_i_5
       (.I0(\u0/R2 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [19]),
        .I3(\u0/uk/K_r2 [24]),
        .O(\u0/u3/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__30_i_6
       (.I0(\u0/R2 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r2 [25]),
        .I3(\u0/uk/K_r2 [5]),
        .O(\u0/u3/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__31
       (.I0(\u0/u4/X [41]),
        .I1(\u0/u4/X [40]),
        .I2(\u0/u4/X [39]),
        .I3(\u0/u4/X [38]),
        .I4(\u0/u4/X [42]),
        .I5(\u0/u4/X [37]),
        .O(\u0/out4 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__310
       (.I0(\u2/u6/X [5]),
        .I1(\u2/u6/X [4]),
        .I2(\u2/u6/X [3]),
        .I3(\u2/u6/X [2]),
        .I4(\u2/u6/X [6]),
        .I5(\u2/u6/X [1]),
        .O(\u2/out6 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__310_i_1
       (.I0(\u2/R5 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [33]),
        .I3(\u2/uk/K_r5 [11]),
        .O(\u2/u6/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__310_i_2
       (.I0(\u2/R5 [3]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [55]),
        .I3(\u2/uk/K_r5 [33]),
        .O(\u2/u6/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__310_i_3
       (.I0(\u2/R5 [2]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [46]),
        .I3(\u2/uk/K_r5 [24]),
        .O(\u2/u6/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__310_i_4
       (.I0(\u2/R5 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [6]),
        .I3(\u2/uk/K_r5 [41]),
        .O(\u2/u6/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__310_i_5
       (.I0(\u2/R5 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [4]),
        .I3(\u2/uk/K_r5 [39]),
        .O(\u2/u6/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__310_i_6
       (.I0(\u2/R5 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r5 [10]),
        .I3(\u2/uk/K_r5 [20]),
        .O(\u2/u6/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__311
       (.I0(\u2/u7/X [41]),
        .I1(\u2/u7/X [40]),
        .I2(\u2/u7/X [39]),
        .I3(\u2/u7/X [38]),
        .I4(\u2/u7/X [42]),
        .I5(\u2/u7/X [37]),
        .O(\u2/out7 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__311_i_1
       (.I0(\u2/R6 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[23] ),
        .I3(\u2/uk/K_r6_reg_n_0_[30] ),
        .O(\u2/u7/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__311_i_2
       (.I0(\u2/R6 [27]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[36] ),
        .I3(\u2/uk/p_45_in ),
        .O(\u2/u7/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__311_i_3
       (.I0(\u2/R6 [26]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[31] ),
        .I3(\u2/uk/K_r6_reg_n_0_[38] ),
        .O(\u2/u7/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__311_i_4
       (.I0(\u2/R6 [25]),
        .I1(decrypt),
        .I2(\u2/uk/p_41_in ),
        .I3(\u2/uk/p_43_in ),
        .O(\u2/u7/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__311_i_5
       (.I0(\u2/R6 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[15] ),
        .I3(\u2/uk/K_r6_reg_n_0_[22] ),
        .O(\u2/u7/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__311_i_6
       (.I0(\u2/R6 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[7] ),
        .I3(\u2/uk/K_r6_reg_n_0_[14] ),
        .O(\u2/u7/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__312
       (.I0(\u2/u7/X [17]),
        .I1(\u2/u7/X [16]),
        .I2(\u2/u7/X [15]),
        .I3(\u2/u7/X [14]),
        .I4(\u2/u7/X [18]),
        .I5(\u2/u7/X [13]),
        .O(\u2/out7 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__312_i_1
       (.I0(\u2/R6 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[26] ),
        .I3(\u2/uk/K_r6_reg_n_0_[33] ),
        .O(\u2/u7/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__312_i_2
       (.I0(\u2/R6 [11]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[11] ),
        .I3(\u2/uk/K_r6_reg_n_0_[18] ),
        .O(\u2/u7/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__312_i_3
       (.I0(\u2/R6 [10]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[10] ),
        .I3(\u2/uk/K_r6_reg_n_0_[17] ),
        .O(\u2/u7/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__312_i_4
       (.I0(\u2/R6 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[34] ),
        .I3(\u2/uk/K_r6_reg_n_0_[41] ),
        .O(\u2/u7/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__312_i_5
       (.I0(\u2/R6 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[39] ),
        .I3(\u2/uk/K_r6_reg_n_0_[46] ),
        .O(\u2/u7/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__312_i_6
       (.I0(\u2/R6 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[5] ),
        .I3(\u2/uk/K_r6_reg_n_0_[12] ),
        .O(\u2/u7/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__313
       (.I0(\u2/u7/X [35]),
        .I1(\u2/u7/X [34]),
        .I2(\u2/u7/X [33]),
        .I3(\u2/u7/X [32]),
        .I4(\u2/u7/X [36]),
        .I5(\u2/u7/X [31]),
        .O(\u2/out7 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__313_i_1
       (.I0(\u2/R6 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[16] ),
        .I3(\u2/uk/K_r6_reg_n_0_[23] ),
        .O(\u2/u7/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__313_i_2
       (.I0(\u2/R6 [23]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[14] ),
        .I3(\u2/uk/K_r6_reg_n_0_[21] ),
        .O(\u2/u7/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__313_i_3
       (.I0(\u2/R6 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[1] ),
        .I3(\u2/uk/K_r6_reg_n_0_[8] ),
        .O(\u2/u7/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__313_i_4
       (.I0(\u2/R6 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[38] ),
        .I3(\u2/uk/K_r6_reg_n_0_[45] ),
        .O(\u2/u7/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__313_i_5
       (.I0(\u2/R6 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[35] ),
        .I3(\u2/uk/p_41_in ),
        .O(\u2/u7/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__313_i_6
       (.I0(\u2/R6 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[50] ),
        .I3(\u2/uk/K_r6_reg_n_0_[2] ),
        .O(\u2/u7/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__314
       (.I0(\u2/u7/X [11]),
        .I1(\u2/u7/X [10]),
        .I2(\u2/u7/X [9]),
        .I3(\u2/u7/X [8]),
        .I4(\u2/u7/X [12]),
        .I5(\u2/u7/X [7]),
        .O(\u2/out7 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__314_i_1
       (.I0(\u2/R6 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[48] ),
        .I3(\u2/uk/K_r6_reg_n_0_[55] ),
        .O(\u2/u7/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__314_i_2
       (.I0(\u2/R6 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[25] ),
        .I3(\u2/uk/K_r6_reg_n_0_[32] ),
        .O(\u2/u7/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__314_i_3
       (.I0(\u2/R6 [6]),
        .I1(decrypt),
        .I2(\u2/uk/p_53_in ),
        .I3(\u2/uk/p_52_in ),
        .O(\u2/u7/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__314_i_4
       (.I0(\u2/R6 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[40] ),
        .I3(\u2/uk/K_r6_reg_n_0_[47] ),
        .O(\u2/u7/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__314_i_5
       (.I0(\u2/R6 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[53] ),
        .I3(\u2/uk/K_r6_reg_n_0_[3] ),
        .O(\u2/u7/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__314_i_6
       (.I0(\u2/R6 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[4] ),
        .I3(\u2/uk/K_r6_reg_n_0_[11] ),
        .O(\u2/u7/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__315
       (.I0(\u2/u7/X [47]),
        .I1(\u2/u7/X [46]),
        .I2(\u2/u7/X [45]),
        .I3(\u2/u7/X [44]),
        .I4(\u2/u7/X [48]),
        .I5(\u2/u7/X [43]),
        .O(\u2/out7 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__315_i_1
       (.I0(\u2/R6 [32]),
        .I1(decrypt),
        .I2(\u2/uk/p_45_in ),
        .I3(\u2/uk/K_r6_reg_n_0_[50] ),
        .O(\u2/u7/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__315_i_2
       (.I0(\u2/R6 [31]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[37] ),
        .I3(\u2/uk/K_r6_reg_n_0_[44] ),
        .O(\u2/u7/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__315_i_3
       (.I0(\u2/R6 [30]),
        .I1(decrypt),
        .I2(\u2/uk/p_43_in ),
        .I3(\u2/uk/K_r6_reg_n_0_[1] ),
        .O(\u2/u7/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__315_i_4
       (.I0(\u2/R6 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[52] ),
        .I3(\u2/uk/K_r6_reg_n_0_ ),
        .O(\u2/u7/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__315_i_5
       (.I0(\u2/R6 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[9] ),
        .I3(\u2/uk/K_r6_reg_n_0_[16] ),
        .O(\u2/u7/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__315_i_6
       (.I0(\u2/R6 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[21] ),
        .I3(\u2/uk/K_r6_reg_n_0_[28] ),
        .O(\u2/u7/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__316
       (.I0(\u2/u7/X [23]),
        .I1(\u2/u7/X [22]),
        .I2(\u2/u7/X [21]),
        .I3(\u2/u7/X [20]),
        .I4(\u2/u7/X [24]),
        .I5(\u2/u7/X [19]),
        .O(\u2/out7 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__316_i_1
       (.I0(\u2/R6 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[17] ),
        .I3(\u2/uk/K_r6_reg_n_0_[24] ),
        .O(\u2/u7/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__316_i_2
       (.I0(\u2/R6 [15]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[41] ),
        .I3(\u2/uk/K_r6_reg_n_0_[48] ),
        .O(\u2/u7/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__316_i_3
       (.I0(\u2/R6 [14]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[33] ),
        .I3(\u2/uk/K_r6_reg_n_0_[40] ),
        .O(\u2/u7/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__316_i_4
       (.I0(\u2/R6 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[32] ),
        .I3(\u2/uk/K_r6_reg_n_0_[39] ),
        .O(\u2/u7/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__316_i_5
       (.I0(\u2/R6 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[54] ),
        .I3(\u2/uk/K_r6_reg_n_0_[4] ),
        .O(\u2/u7/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__316_i_6
       (.I0(\u2/R6 [12]),
        .I1(decrypt),
        .I2(\u2/uk/p_52_in ),
        .I3(\u2/uk/K_r6_reg_n_0_[20] ),
        .O(\u2/u7/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__317
       (.I0(\u2/u7/X [29]),
        .I1(\u2/u7/X [28]),
        .I2(\u2/u7/X [27]),
        .I3(\u2/u7/X [26]),
        .I4(\u2/u7/X [30]),
        .I5(\u2/u7/X [25]),
        .O(\u2/out7 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__317_i_1
       (.I0(\u2/R6 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[28] ),
        .I3(\u2/uk/K_r6_reg_n_0_[35] ),
        .O(\u2/u7/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__317_i_2
       (.I0(\u2/R6 [19]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[44] ),
        .I3(\u2/uk/K_r6_reg_n_0_[51] ),
        .O(\u2/u7/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__317_i_3
       (.I0(\u2/R6 [18]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[2] ),
        .I3(\u2/uk/K_r6_reg_n_0_[9] ),
        .O(\u2/u7/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__317_i_4
       (.I0(\u2/R6 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[8] ),
        .I3(\u2/uk/K_r6_reg_n_0_[15] ),
        .O(\u2/u7/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__317_i_5
       (.I0(\u2/R6 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[29] ),
        .I3(\u2/uk/K_r6_reg_n_0_[36] ),
        .O(\u2/u7/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__317_i_6
       (.I0(\u2/R6 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[45] ),
        .I3(\u2/uk/K_r6_reg_n_0_[52] ),
        .O(\u2/u7/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__318
       (.I0(\u2/u7/X [5]),
        .I1(\u2/u7/X [4]),
        .I2(\u2/u7/X [3]),
        .I3(\u2/u7/X [2]),
        .I4(\u2/u7/X [6]),
        .I5(\u2/u7/X [1]),
        .O(\u2/out7 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__318_i_1
       (.I0(\u2/R6 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[47] ),
        .I3(\u2/uk/K_r6_reg_n_0_[54] ),
        .O(\u2/u7/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__318_i_2
       (.I0(\u2/R6 [3]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[12] ),
        .I3(\u2/uk/K_r6_reg_n_0_[19] ),
        .O(\u2/u7/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__318_i_3
       (.I0(\u2/R6 [2]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[3] ),
        .I3(\u2/uk/K_r6_reg_n_0_[10] ),
        .O(\u2/u7/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__318_i_4
       (.I0(\u2/R6 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[20] ),
        .I3(\u2/uk/K_r6_reg_n_0_[27] ),
        .O(\u2/u7/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__318_i_5
       (.I0(\u2/R6 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[18] ),
        .I3(\u2/uk/K_r6_reg_n_0_[25] ),
        .O(\u2/u7/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__318_i_6
       (.I0(\u2/R6 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r6_reg_n_0_[24] ),
        .I3(\u2/uk/p_53_in ),
        .O(\u2/u7/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__319
       (.I0(\u2/u8/X [41]),
        .I1(\u2/u8/X [40]),
        .I2(\u2/u8/X [39]),
        .I3(\u2/u8/X [38]),
        .I4(\u2/u8/X [42]),
        .I5(\u2/u8/X [37]),
        .O(\u2/out8 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__319_i_1
       (.I0(\u2/R7 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[30] ),
        .I3(\u2/uk/K_r7_reg_n_0_[23] ),
        .O(\u2/u8/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__319_i_2
       (.I0(\u2/R7 [27]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[43] ),
        .I3(\u2/uk/K_r7_reg_n_0_[36] ),
        .O(\u2/u8/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__319_i_3
       (.I0(\u2/R7 [26]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[38] ),
        .I3(\u2/uk/K_r7_reg_n_0_[31] ),
        .O(\u2/u8/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__319_i_4
       (.I0(\u2/R7 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[49] ),
        .I3(\u2/uk/K_r7_reg_n_0_[42] ),
        .O(\u2/u8/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__319_i_5
       (.I0(\u2/R7 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[22] ),
        .I3(\u2/uk/K_r7_reg_n_0_[15] ),
        .O(\u2/u8/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__319_i_6
       (.I0(\u2/R7 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[14] ),
        .I3(\u2/uk/K_r7_reg_n_0_[7] ),
        .O(\u2/u8/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__31_i_1
       (.I0(\u0/R3 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [36]),
        .I3(\u0/uk/K_r3 [45]),
        .O(\u0/u4/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__31_i_2
       (.I0(\u0/R3 [27]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [49]),
        .I3(\u0/uk/K_r3 [30]),
        .O(\u0/u4/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__31_i_3
       (.I0(\u0/R3 [26]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [16]),
        .I3(\u0/uk/K_r3 [21]),
        .O(\u0/u4/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__31_i_4
       (.I0(\u0/R3 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [0]),
        .I3(\u0/uk/K_r3 [36]),
        .O(\u0/u4/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__31_i_5
       (.I0(\u0/R3 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [28]),
        .I3(\u0/uk/K_r3 [9]),
        .O(\u0/u4/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__31_i_6
       (.I0(\u0/R3 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [51]),
        .I3(\u0/uk/K_r3 [1]),
        .O(\u0/u4/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__32
       (.I0(\u0/u4/X [17]),
        .I1(\u0/u4/X [16]),
        .I2(\u0/u4/X [15]),
        .I3(\u0/u4/X [14]),
        .I4(\u0/u4/X [18]),
        .I5(\u0/u4/X [13]),
        .O(\u0/out4 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__320
       (.I0(\u2/u8/X [17]),
        .I1(\u2/u8/X [16]),
        .I2(\u2/u8/X [15]),
        .I3(\u2/u8/X [14]),
        .I4(\u2/u8/X [18]),
        .I5(\u2/u8/X [13]),
        .O(\u2/out8 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__320_i_1
       (.I0(\u2/R7 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[33] ),
        .I3(\u2/uk/K_r7_reg_n_0_[26] ),
        .O(\u2/u8/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__320_i_2
       (.I0(\u2/R7 [11]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[18] ),
        .I3(\u2/uk/K_r7_reg_n_0_[11] ),
        .O(\u2/u8/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__320_i_3
       (.I0(\u2/R7 [10]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[17] ),
        .I3(\u2/uk/K_r7_reg_n_0_[10] ),
        .O(\u2/u8/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__320_i_4
       (.I0(\u2/R7 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[41] ),
        .I3(\u2/uk/K_r7_reg_n_0_[34] ),
        .O(\u2/u8/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__320_i_5
       (.I0(\u2/R7 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[46] ),
        .I3(\u2/uk/K_r7_reg_n_0_[39] ),
        .O(\u2/u8/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__320_i_6
       (.I0(\u2/R7 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[12] ),
        .I3(\u2/uk/K_r7_reg_n_0_[5] ),
        .O(\u2/u8/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__321
       (.I0(\u2/u8/X [35]),
        .I1(\u2/u8/X [34]),
        .I2(\u2/u8/X [33]),
        .I3(\u2/u8/X [32]),
        .I4(\u2/u8/X [36]),
        .I5(\u2/u8/X [31]),
        .O(\u2/out8 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__321_i_1
       (.I0(\u2/R7 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[23] ),
        .I3(\u2/uk/K_r7_reg_n_0_[16] ),
        .O(\u2/u8/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__321_i_2
       (.I0(\u2/R7 [23]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[21] ),
        .I3(\u2/uk/K_r7_reg_n_0_[14] ),
        .O(\u2/u8/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__321_i_3
       (.I0(\u2/R7 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[8] ),
        .I3(\u2/uk/K_r7_reg_n_0_[1] ),
        .O(\u2/u8/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__321_i_4
       (.I0(\u2/R7 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[45] ),
        .I3(\u2/uk/K_r7_reg_n_0_[38] ),
        .O(\u2/u8/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__321_i_5
       (.I0(\u2/R7 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[42] ),
        .I3(\u2/uk/K_r7_reg_n_0_[35] ),
        .O(\u2/u8/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__321_i_6
       (.I0(\u2/R7 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[2] ),
        .I3(\u2/uk/K_r7_reg_n_0_[50] ),
        .O(\u2/u8/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__322
       (.I0(\u2/u8/X [11]),
        .I1(\u2/u8/X [10]),
        .I2(\u2/u8/X [9]),
        .I3(\u2/u8/X [8]),
        .I4(\u2/u8/X [12]),
        .I5(\u2/u8/X [7]),
        .O(\u2/out8 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__322_i_1
       (.I0(\u2/R7 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[55] ),
        .I3(\u2/uk/K_r7_reg_n_0_[48] ),
        .O(\u2/u8/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__322_i_2
       (.I0(\u2/R7 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[32] ),
        .I3(\u2/uk/K_r7_reg_n_0_[25] ),
        .O(\u2/u8/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__322_i_3
       (.I0(\u2/R7 [6]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[13] ),
        .I3(\u2/uk/K_r7_reg_n_0_[6] ),
        .O(\u2/u8/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__322_i_4
       (.I0(\u2/R7 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[47] ),
        .I3(\u2/uk/K_r7_reg_n_0_[40] ),
        .O(\u2/u8/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__322_i_5
       (.I0(\u2/R7 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[3] ),
        .I3(\u2/uk/K_r7_reg_n_0_[53] ),
        .O(\u2/u8/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__322_i_6
       (.I0(\u2/R7 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[11] ),
        .I3(\u2/uk/K_r7_reg_n_0_[4] ),
        .O(\u2/u8/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__323
       (.I0(\u2/u8/X [47]),
        .I1(\u2/u8/X [46]),
        .I2(\u2/u8/X [45]),
        .I3(\u2/u8/X [44]),
        .I4(\u2/u8/X [48]),
        .I5(\u2/u8/X [43]),
        .O(\u2/out8 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__323_i_1
       (.I0(\u2/R7 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[50] ),
        .I3(\u2/uk/K_r7_reg_n_0_[43] ),
        .O(\u2/u8/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__323_i_2
       (.I0(\u2/R7 [31]),
        .I1(decrypt),
        .I2(\u2/uk/p_48_in ),
        .I3(\u2/uk/K_r7_reg_n_0_[37] ),
        .O(\u2/u8/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__323_i_3
       (.I0(\u2/R7 [30]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[1] ),
        .I3(\u2/uk/K_r7_reg_n_0_[49] ),
        .O(\u2/u8/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__323_i_4
       (.I0(\u2/R7 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_ ),
        .I3(\u2/uk/K_r7_reg_n_0_[52] ),
        .O(\u2/u8/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__323_i_5
       (.I0(\u2/R7 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[16] ),
        .I3(\u2/uk/K_r7_reg_n_0_[9] ),
        .O(\u2/u8/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__323_i_6
       (.I0(\u2/R7 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[28] ),
        .I3(\u2/uk/K_r7_reg_n_0_[21] ),
        .O(\u2/u8/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__324
       (.I0(\u2/u8/X [23]),
        .I1(\u2/u8/X [22]),
        .I2(\u2/u8/X [21]),
        .I3(\u2/u8/X [20]),
        .I4(\u2/u8/X [24]),
        .I5(\u2/u8/X [19]),
        .O(\u2/out8 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__324_i_1
       (.I0(\u2/R7 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[24] ),
        .I3(\u2/uk/K_r7_reg_n_0_[17] ),
        .O(\u2/u8/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__324_i_2
       (.I0(\u2/R7 [15]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[48] ),
        .I3(\u2/uk/K_r7_reg_n_0_[41] ),
        .O(\u2/u8/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__324_i_3
       (.I0(\u2/R7 [14]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[40] ),
        .I3(\u2/uk/K_r7_reg_n_0_[33] ),
        .O(\u2/u8/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__324_i_4
       (.I0(\u2/R7 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[39] ),
        .I3(\u2/uk/K_r7_reg_n_0_[32] ),
        .O(\u2/u8/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__324_i_5
       (.I0(\u2/R7 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[4] ),
        .I3(\u2/uk/K_r7_reg_n_0_[54] ),
        .O(\u2/u8/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__324_i_6
       (.I0(\u2/R7 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[20] ),
        .I3(\u2/uk/K_r7_reg_n_0_[13] ),
        .O(\u2/u8/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__325
       (.I0(\u2/u8/X [29]),
        .I1(\u2/u8/X [28]),
        .I2(\u2/u8/X [27]),
        .I3(\u2/u8/X [26]),
        .I4(\u2/u8/X [30]),
        .I5(\u2/u8/X [25]),
        .O(\u2/out8 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__325_i_1
       (.I0(\u2/R7 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[35] ),
        .I3(\u2/uk/K_r7_reg_n_0_[28] ),
        .O(\u2/u8/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__325_i_2
       (.I0(\u2/R7 [19]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[51] ),
        .I3(\u2/uk/p_48_in ),
        .O(\u2/u8/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__325_i_3
       (.I0(\u2/R7 [18]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[9] ),
        .I3(\u2/uk/K_r7_reg_n_0_[2] ),
        .O(\u2/u8/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__325_i_4
       (.I0(\u2/R7 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[15] ),
        .I3(\u2/uk/K_r7_reg_n_0_[8] ),
        .O(\u2/u8/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__325_i_5
       (.I0(\u2/R7 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[36] ),
        .I3(\u2/uk/K_r7_reg_n_0_[29] ),
        .O(\u2/u8/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__325_i_6
       (.I0(\u2/R7 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[52] ),
        .I3(\u2/uk/K_r7_reg_n_0_[45] ),
        .O(\u2/u8/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__326
       (.I0(\u2/u8/X [5]),
        .I1(\u2/u8/X [4]),
        .I2(\u2/u8/X [3]),
        .I3(\u2/u8/X [2]),
        .I4(\u2/u8/X [6]),
        .I5(\u2/u8/X [1]),
        .O(\u2/out8 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__326_i_1
       (.I0(\u2/R7 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[54] ),
        .I3(\u2/uk/K_r7_reg_n_0_[47] ),
        .O(\u2/u8/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__326_i_2
       (.I0(\u2/R7 [3]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[19] ),
        .I3(\u2/uk/K_r7_reg_n_0_[12] ),
        .O(\u2/u8/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__326_i_3
       (.I0(\u2/R7 [2]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[10] ),
        .I3(\u2/uk/K_r7_reg_n_0_[3] ),
        .O(\u2/u8/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__326_i_4
       (.I0(\u2/R7 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[27] ),
        .I3(\u2/uk/K_r7_reg_n_0_[20] ),
        .O(\u2/u8/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__326_i_5
       (.I0(\u2/R7 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[25] ),
        .I3(\u2/uk/K_r7_reg_n_0_[18] ),
        .O(\u2/u8/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__326_i_6
       (.I0(\u2/R7 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r7_reg_n_0_[6] ),
        .I3(\u2/uk/K_r7_reg_n_0_[24] ),
        .O(\u2/u8/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__327
       (.I0(\u2/u9/X [41]),
        .I1(\u2/u9/X [40]),
        .I2(\u2/u9/X [39]),
        .I3(\u2/u9/X [38]),
        .I4(\u2/u9/X [42]),
        .I5(\u2/u9/X [37]),
        .O(\u2/out9 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__327_i_1
       (.I0(\u2/R8 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [44]),
        .I3(\u2/uk/K_r8 [9]),
        .O(\u2/u9/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__327_i_2
       (.I0(\u2/R8 [27]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [2]),
        .I3(\u2/uk/K_r8 [22]),
        .O(\u2/u9/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__327_i_3
       (.I0(\u2/R8 [26]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [52]),
        .I3(\u2/uk/K_r8 [44]),
        .O(\u2/u9/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__327_i_4
       (.I0(\u2/R8 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [8]),
        .I3(\u2/uk/K_r8 [28]),
        .O(\u2/u9/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__327_i_5
       (.I0(\u2/R8 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [36]),
        .I3(\u2/uk/K_r8 [1]),
        .O(\u2/u9/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__327_i_6
       (.I0(\u2/R8 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [28]),
        .I3(\u2/uk/K_r8 [52]),
        .O(\u2/u9/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__328
       (.I0(\u2/u9/X [17]),
        .I1(\u2/u9/X [16]),
        .I2(\u2/u9/X [15]),
        .I3(\u2/u9/X [14]),
        .I4(\u2/u9/X [18]),
        .I5(\u2/u9/X [13]),
        .O(\u2/out9 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__328_i_1
       (.I0(\u2/R8 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [47]),
        .I3(\u2/uk/K_r8 [12]),
        .O(\u2/u9/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__328_i_2
       (.I0(\u2/R8 [11]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [32]),
        .I3(\u2/uk/K_r8 [54]),
        .O(\u2/u9/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__328_i_3
       (.I0(\u2/R8 [10]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [6]),
        .I3(\u2/uk/K_r8 [53]),
        .O(\u2/u9/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__328_i_4
       (.I0(\u2/R8 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [55]),
        .I3(\u2/uk/K_r8 [20]),
        .O(\u2/u9/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__328_i_5
       (.I0(\u2/R8 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [3]),
        .I3(\u2/uk/K_r8 [25]),
        .O(\u2/u9/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__328_i_6
       (.I0(\u2/R8 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [26]),
        .I3(\u2/uk/K_r8 [48]),
        .O(\u2/u9/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__329
       (.I0(\u2/u9/X [35]),
        .I1(\u2/u9/X [34]),
        .I2(\u2/u9/X [33]),
        .I3(\u2/u9/X [32]),
        .I4(\u2/u9/X [36]),
        .I5(\u2/u9/X [31]),
        .O(\u2/out9 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__329_i_1
       (.I0(\u2/R8 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [37]),
        .I3(\u2/uk/K_r8 [2]),
        .O(\u2/u9/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__329_i_2
       (.I0(\u2/R8 [23]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [35]),
        .I3(\u2/uk/K_r8 [0]),
        .O(\u2/u9/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__329_i_3
       (.I0(\u2/R8 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [22]),
        .I3(\u2/uk/K_r8 [42]),
        .O(\u2/u9/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__329_i_4
       (.I0(\u2/R8 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [0]),
        .I3(\u2/uk/K_r8 [51]),
        .O(\u2/u9/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__329_i_5
       (.I0(\u2/R8 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [1]),
        .I3(\u2/uk/K_r8 [21]),
        .O(\u2/u9/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__329_i_6
       (.I0(\u2/R8 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [16]),
        .I3(\u2/uk/K_r8 [36]),
        .O(\u2/u9/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__32_i_1
       (.I0(\u0/R3 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [41]),
        .I3(\u0/uk/K_r3 [18]),
        .O(\u0/u4/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__32_i_2
       (.I0(\u0/R3 [11]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [26]),
        .I3(\u0/uk/K_r3 [3]),
        .O(\u0/u4/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__32_i_3
       (.I0(\u0/R3 [10]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [25]),
        .I3(\u0/uk/K_r3 [34]),
        .O(\u0/u4/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__32_i_4
       (.I0(\u0/R3 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [17]),
        .I3(\u0/uk/K_r3 [26]),
        .O(\u0/u4/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__32_i_5
       (.I0(\u0/R3 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [54]),
        .I3(\u0/uk/K_r3 [6]),
        .O(\u0/u4/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__32_i_6
       (.I0(\u0/R3 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [20]),
        .I3(\u0/uk/K_r3 [54]),
        .O(\u0/u4/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__33
       (.I0(\u0/u4/X [35]),
        .I1(\u0/u4/X [34]),
        .I2(\u0/u4/X [33]),
        .I3(\u0/u4/X [32]),
        .I4(\u0/u4/X [36]),
        .I5(\u0/u4/X [31]),
        .O(\u0/out4 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__330
       (.I0(\u2/u9/X [11]),
        .I1(\u2/u9/X [10]),
        .I2(\u2/u9/X [9]),
        .I3(\u2/u9/X [8]),
        .I4(\u2/u9/X [12]),
        .I5(\u2/u9/X [7]),
        .O(\u2/out9 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__330_i_1
       (.I0(\u2/R8 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [12]),
        .I3(\u2/uk/K_r8 [34]),
        .O(\u2/u9/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__330_i_2
       (.I0(\u2/R8 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [46]),
        .I3(\u2/uk/K_r8 [11]),
        .O(\u2/u9/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__330_i_3
       (.I0(\u2/R8 [6]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [27]),
        .I3(\u2/uk/K_r8 [17]),
        .O(\u2/u9/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__330_i_4
       (.I0(\u2/R8 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [4]),
        .I3(\u2/uk/K_r8 [26]),
        .O(\u2/u9/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__330_i_5
       (.I0(\u2/R8 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [17]),
        .I3(\u2/uk/K_r8 [39]),
        .O(\u2/u9/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__330_i_6
       (.I0(\u2/R8 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [25]),
        .I3(\u2/uk/K_r8 [47]),
        .O(\u2/u9/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__331
       (.I0(\u2/u9/X [47]),
        .I1(\u2/u9/X [46]),
        .I2(\u2/u9/X [45]),
        .I3(\u2/u9/X [44]),
        .I4(\u2/u9/X [48]),
        .I5(\u2/u9/X [43]),
        .O(\u2/out9 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__331_i_1
       (.I0(\u2/R8 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [9]),
        .I3(\u2/uk/K_r8 [29]),
        .O(\u2/u9/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__331_i_2
       (.I0(\u2/R8 [31]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [31]),
        .I3(\u2/uk/K_r8 [23]),
        .O(\u2/u9/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__331_i_3
       (.I0(\u2/R8 [30]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [15]),
        .I3(\u2/uk/K_r8 [35]),
        .O(\u2/u9/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__331_i_4
       (.I0(\u2/R8 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [14]),
        .I3(\u2/uk/K_r8 [38]),
        .O(\u2/u9/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__331_i_5
       (.I0(\u2/R8 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [30]),
        .I3(\u2/uk/K_r8 [50]),
        .O(\u2/u9/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__331_i_6
       (.I0(\u2/R8 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [42]),
        .I3(\u2/uk/K_r8 [7]),
        .O(\u2/u9/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__332
       (.I0(\u2/u9/X [23]),
        .I1(\u2/u9/X [22]),
        .I2(\u2/u9/X [21]),
        .I3(\u2/u9/X [20]),
        .I4(\u2/u9/X [24]),
        .I5(\u2/u9/X [19]),
        .O(\u2/out9 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__332_i_1
       (.I0(\u2/R8 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [13]),
        .I3(\u2/uk/K_r8 [3]),
        .O(\u2/u9/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__332_i_2
       (.I0(\u2/R8 [15]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [5]),
        .I3(\u2/uk/K_r8 [27]),
        .O(\u2/u9/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__332_i_3
       (.I0(\u2/R8 [14]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [54]),
        .I3(\u2/uk/K_r8 [19]),
        .O(\u2/u9/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__332_i_4
       (.I0(\u2/R8 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [53]),
        .I3(\u2/uk/K_r8 [18]),
        .O(\u2/u9/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__332_i_5
       (.I0(\u2/R8 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [18]),
        .I3(\u2/uk/K_r8 [40]),
        .O(\u2/u9/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__332_i_6
       (.I0(\u2/R8 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [34]),
        .I3(\u2/uk/K_r8 [24]),
        .O(\u2/u9/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__333
       (.I0(\u2/u9/X [29]),
        .I1(\u2/u9/X [28]),
        .I2(\u2/u9/X [27]),
        .I3(\u2/u9/X [26]),
        .I4(\u2/u9/X [30]),
        .I5(\u2/u9/X [25]),
        .O(\u2/out9 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__333_i_1
       (.I0(\u2/R8 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [49]),
        .I3(\u2/uk/K_r8 [14]),
        .O(\u2/u9/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__333_i_2
       (.I0(\u2/R8 [19]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [38]),
        .I3(\u2/uk/K_r8 [30]),
        .O(\u2/u9/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__333_i_3
       (.I0(\u2/R8 [18]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [23]),
        .I3(\u2/uk/K_r8 [43]),
        .O(\u2/u9/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__333_i_4
       (.I0(\u2/R8 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [29]),
        .I3(\u2/uk/K_r8 [49]),
        .O(\u2/u9/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__333_i_5
       (.I0(\u2/R8 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [50]),
        .I3(\u2/uk/K_r8 [15]),
        .O(\u2/u9/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__333_i_6
       (.I0(\u2/R8 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [7]),
        .I3(\u2/uk/K_r8 [31]),
        .O(\u2/u9/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__334
       (.I0(\u2/u9/X [5]),
        .I1(\u2/u9/X [4]),
        .I2(\u2/u9/X [3]),
        .I3(\u2/u9/X [2]),
        .I4(\u2/u9/X [6]),
        .I5(\u2/u9/X [1]),
        .O(\u2/out9 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__334_i_1
       (.I0(\u2/R8 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [11]),
        .I3(\u2/uk/K_r8 [33]),
        .O(\u2/u9/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__334_i_2
       (.I0(\u2/R8 [3]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [33]),
        .I3(\u2/uk/K_r8 [55]),
        .O(\u2/u9/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__334_i_3
       (.I0(\u2/R8 [2]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [24]),
        .I3(\u2/uk/K_r8 [46]),
        .O(\u2/u9/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__334_i_4
       (.I0(\u2/R8 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [41]),
        .I3(\u2/uk/K_r8 [6]),
        .O(\u2/u9/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__334_i_5
       (.I0(\u2/R8 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [39]),
        .I3(\u2/uk/K_r8 [4]),
        .O(\u2/u9/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__334_i_6
       (.I0(\u2/R8 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r8 [20]),
        .I3(\u2/uk/K_r8 [10]),
        .O(\u2/u9/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__335
       (.I0(\u2/u10/X [41]),
        .I1(\u2/u10/X [40]),
        .I2(\u2/u10/X [39]),
        .I3(\u2/u10/X [38]),
        .I4(\u2/u10/X [42]),
        .I5(\u2/u10/X [37]),
        .O(\u2/out10 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__335_i_1
       (.I0(\u2/R9 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [31]),
        .I3(\u2/uk/K_r9 [50]),
        .O(\u2/u10/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__335_i_2
       (.I0(\u2/R9 [27]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [16]),
        .I3(\u2/uk/K_r9 [8]),
        .O(\u2/u10/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__335_i_3
       (.I0(\u2/R9 [26]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [7]),
        .I3(\u2/uk/K_r9 [30]),
        .O(\u2/u10/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__335_i_4
       (.I0(\u2/R9 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [22]),
        .I3(\u2/uk/K_r9 [14]),
        .O(\u2/u10/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__335_i_5
       (.I0(\u2/R9 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [50]),
        .I3(\u2/uk/K_r9 [42]),
        .O(\u2/u10/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__335_i_6
       (.I0(\u2/R9 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [42]),
        .I3(\u2/uk/K_r9 [38]),
        .O(\u2/u10/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__336
       (.I0(\u2/u10/X [17]),
        .I1(\u2/u10/X [16]),
        .I2(\u2/u10/X [15]),
        .I3(\u2/u10/X [14]),
        .I4(\u2/u10/X [18]),
        .I5(\u2/u10/X [13]),
        .O(\u2/out10 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__336_i_1
       (.I0(\u2/R9 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [4]),
        .I3(\u2/uk/K_r9 [55]),
        .O(\u2/u10/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__336_i_2
       (.I0(\u2/R9 [11]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [46]),
        .I3(\u2/uk/K_r9 [40]),
        .O(\u2/u10/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__336_i_3
       (.I0(\u2/R9 [10]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [20]),
        .I3(\u2/uk/K_r9 [39]),
        .O(\u2/u10/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__336_i_4
       (.I0(\u2/R9 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [12]),
        .I3(\u2/uk/K_r9 [6]),
        .O(\u2/u10/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__336_i_5
       (.I0(\u2/R9 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [17]),
        .I3(\u2/uk/K_r9 [11]),
        .O(\u2/u10/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__336_i_6
       (.I0(\u2/R9 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [40]),
        .I3(\u2/uk/K_r9 [34]),
        .O(\u2/u10/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__337
       (.I0(\u2/u10/X [35]),
        .I1(\u2/u10/X [34]),
        .I2(\u2/u10/X [33]),
        .I3(\u2/u10/X [32]),
        .I4(\u2/u10/X [36]),
        .I5(\u2/u10/X [31]),
        .O(\u2/out10 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__337_i_1
       (.I0(\u2/R9 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [51]),
        .I3(\u2/uk/K_r9 [43]),
        .O(\u2/u10/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__337_i_2
       (.I0(\u2/R9 [23]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [49]),
        .I3(\u2/uk/K_r9 [45]),
        .O(\u2/u10/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__337_i_3
       (.I0(\u2/R9 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [36]),
        .I3(\u2/uk/K_r9 [28]),
        .O(\u2/u10/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__337_i_4
       (.I0(\u2/R9 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [14]),
        .I3(\u2/uk/K_r9 [37]),
        .O(\u2/u10/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__337_i_5
       (.I0(\u2/R9 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [15]),
        .I3(\u2/uk/K_r9 [7]),
        .O(\u2/u10/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__337_i_6
       (.I0(\u2/R9 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [30]),
        .I3(\u2/uk/K_r9 [22]),
        .O(\u2/u10/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__338
       (.I0(\u2/u10/X [11]),
        .I1(\u2/u10/X [10]),
        .I2(\u2/u10/X [9]),
        .I3(\u2/u10/X [8]),
        .I4(\u2/u10/X [12]),
        .I5(\u2/u10/X [7]),
        .O(\u2/out10 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__338_i_1
       (.I0(\u2/R9 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [26]),
        .I3(\u2/uk/K_r9 [20]),
        .O(\u2/u10/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__338_i_2
       (.I0(\u2/R9 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [3]),
        .I3(\u2/uk/K_r9 [54]),
        .O(\u2/u10/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__338_i_3
       (.I0(\u2/R9 [6]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [41]),
        .I3(\u2/uk/K_r9 [3]),
        .O(\u2/u10/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__338_i_4
       (.I0(\u2/R9 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [18]),
        .I3(\u2/uk/K_r9 [12]),
        .O(\u2/u10/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__338_i_5
       (.I0(\u2/R9 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [6]),
        .I3(\u2/uk/K_r9 [25]),
        .O(\u2/u10/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__338_i_6
       (.I0(\u2/R9 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [39]),
        .I3(\u2/uk/K_r9 [33]),
        .O(\u2/u10/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__339
       (.I0(\u2/u10/X [47]),
        .I1(\u2/u10/X [46]),
        .I2(\u2/u10/X [45]),
        .I3(\u2/u10/X [44]),
        .I4(\u2/u10/X [48]),
        .I5(\u2/u10/X [43]),
        .O(\u2/out10 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__339_i_1
       (.I0(\u2/R9 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [23]),
        .I3(\u2/uk/K_r9 [15]),
        .O(\u2/u10/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__339_i_2
       (.I0(\u2/R9 [31]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [45]),
        .I3(\u2/uk/K_r9 [9]),
        .O(\u2/u10/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__339_i_3
       (.I0(\u2/R9 [30]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [29]),
        .I3(\u2/uk/K_r9 [21]),
        .O(\u2/u10/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__339_i_4
       (.I0(\u2/R9 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [28]),
        .I3(\u2/uk/K_r9 [51]),
        .O(\u2/u10/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__339_i_5
       (.I0(\u2/R9 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [44]),
        .I3(\u2/uk/K_r9 [36]),
        .O(\u2/u10/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__339_i_6
       (.I0(\u2/R9 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [1]),
        .I3(\u2/uk/K_r9 [52]),
        .O(\u2/u10/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__33_i_1
       (.I0(\u0/R3 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [29]),
        .I3(\u0/uk/K_r3 [38]),
        .O(\u0/u4/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__33_i_2
       (.I0(\u0/R3 [23]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [31]),
        .I3(\u0/uk/K_r3 [8]),
        .O(\u0/u4/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__33_i_3
       (.I0(\u0/R3 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [14]),
        .I3(\u0/uk/K_r3 [50]),
        .O(\u0/u4/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__33_i_4
       (.I0(\u0/R3 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [23]),
        .I3(\u0/uk/K_r3 [28]),
        .O(\u0/u4/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__33_i_5
       (.I0(\u0/R3 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [52]),
        .I3(\u0/uk/K_r3 [29]),
        .O(\u0/u4/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__33_i_6
       (.I0(\u0/R3 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [8]),
        .I3(\u0/uk/K_r3 [44]),
        .O(\u0/u4/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__34
       (.I0(\u0/u4/X [11]),
        .I1(\u0/u4/X [10]),
        .I2(\u0/u4/X [9]),
        .I3(\u0/u4/X [8]),
        .I4(\u0/u4/X [12]),
        .I5(\u0/u4/X [7]),
        .O(\u0/out4 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__340
       (.I0(\u2/u10/X [23]),
        .I1(\u2/u10/X [22]),
        .I2(\u2/u10/X [21]),
        .I3(\u2/u10/X [20]),
        .I4(\u2/u10/X [24]),
        .I5(\u2/u10/X [19]),
        .O(\u2/out10 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__340_i_1
       (.I0(\u2/R9 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [27]),
        .I3(\u2/uk/K_r9 [46]),
        .O(\u2/u10/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__340_i_2
       (.I0(\u2/R9 [15]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [19]),
        .I3(\u2/uk/K_r9 [13]),
        .O(\u2/u10/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__340_i_3
       (.I0(\u2/R9 [14]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [11]),
        .I3(\u2/uk/K_r9 [5]),
        .O(\u2/u10/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__340_i_4
       (.I0(\u2/R9 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [10]),
        .I3(\u2/uk/K_r9 [4]),
        .O(\u2/u10/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__340_i_5
       (.I0(\u2/R9 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [32]),
        .I3(\u2/uk/K_r9 [26]),
        .O(\u2/u10/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__340_i_6
       (.I0(\u2/R9 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [48]),
        .I3(\u2/uk/K_r9 [10]),
        .O(\u2/u10/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__341
       (.I0(\u2/u10/X [29]),
        .I1(\u2/u10/X [28]),
        .I2(\u2/u10/X [27]),
        .I3(\u2/u10/X [26]),
        .I4(\u2/u10/X [30]),
        .I5(\u2/u10/X [25]),
        .O(\u2/out10 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__341_i_1
       (.I0(\u2/R9 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [8]),
        .I3(\u2/uk/K_r9 [0]),
        .O(\u2/u10/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__341_i_2
       (.I0(\u2/R9 [19]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [52]),
        .I3(\u2/uk/K_r9 [16]),
        .O(\u2/u10/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__341_i_3
       (.I0(\u2/R9 [18]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [37]),
        .I3(\u2/uk/K_r9 [29]),
        .O(\u2/u10/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__341_i_4
       (.I0(\u2/R9 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [43]),
        .I3(\u2/uk/K_r9 [35]),
        .O(\u2/u10/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__341_i_5
       (.I0(\u2/R9 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [9]),
        .I3(\u2/uk/K_r9 [1]),
        .O(\u2/u10/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__341_i_6
       (.I0(\u2/R9 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [21]),
        .I3(\u2/uk/K_r9 [44]),
        .O(\u2/u10/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__342
       (.I0(\u2/u10/X [5]),
        .I1(\u2/u10/X [4]),
        .I2(\u2/u10/X [3]),
        .I3(\u2/u10/X [2]),
        .I4(\u2/u10/X [6]),
        .I5(\u2/u10/X [1]),
        .O(\u2/out10 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__342_i_1
       (.I0(\u2/R9 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [25]),
        .I3(\u2/uk/K_r9 [19]),
        .O(\u2/u10/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__342_i_2
       (.I0(\u2/R9 [3]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [47]),
        .I3(\u2/uk/K_r9 [41]),
        .O(\u2/u10/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__342_i_3
       (.I0(\u2/R9 [2]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [13]),
        .I3(\u2/uk/K_r9 [32]),
        .O(\u2/u10/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__342_i_4
       (.I0(\u2/R9 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [55]),
        .I3(\u2/uk/K_r9 [17]),
        .O(\u2/u10/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__342_i_5
       (.I0(\u2/R9 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [53]),
        .I3(\u2/uk/K_r9 [47]),
        .O(\u2/u10/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__342_i_6
       (.I0(\u2/R9 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r9 [34]),
        .I3(\u2/uk/K_r9 [53]),
        .O(\u2/u10/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__343
       (.I0(\u2/u11/X [41]),
        .I1(\u2/u11/X [40]),
        .I2(\u2/u11/X [39]),
        .I3(\u2/u11/X [38]),
        .I4(\u2/u11/X [42]),
        .I5(\u2/u11/X [37]),
        .O(\u2/out11 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__343_i_1
       (.I0(\u2/R10_reg_n_0_[28] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [45]),
        .I3(\u2/uk/K_r10 [36]),
        .O(\u2/u11/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__343_i_2
       (.I0(\u2/R10_reg_n_0_[27] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [30]),
        .I3(\u2/uk/K_r10 [49]),
        .O(\u2/u11/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__343_i_3
       (.I0(\u2/R10_reg_n_0_[26] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [21]),
        .I3(\u2/uk/K_r10 [16]),
        .O(\u2/u11/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__343_i_4
       (.I0(\u2/R10_reg_n_0_[25] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [36]),
        .I3(\u2/uk/K_r10 [0]),
        .O(\u2/u11/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__343_i_5
       (.I0(\u2/R10_reg_n_0_[29] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [9]),
        .I3(\u2/uk/K_r10 [28]),
        .O(\u2/u11/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__343_i_6
       (.I0(\u2/R10_reg_n_0_[24] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [1]),
        .I3(\u2/uk/K_r10 [51]),
        .O(\u2/u11/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__344
       (.I0(\u2/u11/X [17]),
        .I1(\u2/u11/X [16]),
        .I2(\u2/u11/X [15]),
        .I3(\u2/u11/X [14]),
        .I4(\u2/u11/X [18]),
        .I5(\u2/u11/X [13]),
        .O(\u2/out11 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__344_i_1
       (.I0(\u2/R10_reg_n_0_[12] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [18]),
        .I3(\u2/uk/K_r10 [41]),
        .O(\u2/u11/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__344_i_2
       (.I0(\u2/R10_reg_n_0_[11] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [3]),
        .I3(\u2/uk/K_r10 [26]),
        .O(\u2/u11/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__344_i_3
       (.I0(\u2/R10_reg_n_0_ ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [34]),
        .I3(\u2/uk/K_r10 [25]),
        .O(\u2/u11/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__344_i_4
       (.I0(\u2/R10_reg_n_0_[9] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [26]),
        .I3(\u2/uk/K_r10 [17]),
        .O(\u2/u11/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__344_i_5
       (.I0(\u2/R10_reg_n_0_[13] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [6]),
        .I3(\u2/uk/K_r10 [54]),
        .O(\u2/u11/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__344_i_6
       (.I0(\u2/R10_reg_n_0_[8] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [54]),
        .I3(\u2/uk/K_r10 [20]),
        .O(\u2/u11/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__345
       (.I0(\u2/u11/X [35]),
        .I1(\u2/u11/X [34]),
        .I2(\u2/u11/X [33]),
        .I3(\u2/u11/X [32]),
        .I4(\u2/u11/X [36]),
        .I5(\u2/u11/X [31]),
        .O(\u2/out11 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__345_i_1
       (.I0(\u2/R10_reg_n_0_[24] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [38]),
        .I3(\u2/uk/K_r10 [29]),
        .O(\u2/u11/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__345_i_2
       (.I0(\u2/R10_reg_n_0_[23] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [8]),
        .I3(\u2/uk/K_r10 [31]),
        .O(\u2/u11/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__345_i_3
       (.I0(\u2/R10_reg_n_0_[22] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [50]),
        .I3(\u2/uk/K_r10 [14]),
        .O(\u2/u11/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__345_i_4
       (.I0(\u2/R10_reg_n_0_[21] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [28]),
        .I3(\u2/uk/K_r10 [23]),
        .O(\u2/u11/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__345_i_5
       (.I0(\u2/R10_reg_n_0_[25] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [29]),
        .I3(\u2/uk/K_r10 [52]),
        .O(\u2/u11/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__345_i_6
       (.I0(\u2/R10_reg_n_0_[20] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [44]),
        .I3(\u2/uk/K_r10 [8]),
        .O(\u2/u11/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__346
       (.I0(\u2/u11/X [11]),
        .I1(\u2/u11/X [10]),
        .I2(\u2/u11/X [9]),
        .I3(\u2/u11/X [8]),
        .I4(\u2/u11/X [12]),
        .I5(\u2/u11/X [7]),
        .O(\u2/out11 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__346_i_1
       (.I0(\u2/R10_reg_n_0_[8] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [40]),
        .I3(\u2/uk/K_r10 [6]),
        .O(\u2/u11/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__346_i_2
       (.I0(\u2/R10_reg_n_0_[7] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [17]),
        .I3(\u2/uk/K_r10 [40]),
        .O(\u2/u11/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__346_i_3
       (.I0(\u2/R10_reg_n_0_[6] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [55]),
        .I3(\u2/uk/K_r10 [46]),
        .O(\u2/u11/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__346_i_4
       (.I0(\u2/R10_reg_n_0_[5] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [32]),
        .I3(\u2/uk/K_r10 [55]),
        .O(\u2/u11/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__346_i_5
       (.I0(\u2/R10_reg_n_0_[9] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [20]),
        .I3(\u2/uk/K_r10 [11]),
        .O(\u2/u11/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__346_i_6
       (.I0(\u2/R10_reg_n_0_[4] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [53]),
        .I3(\u2/uk/K_r10 [19]),
        .O(\u2/u11/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__347
       (.I0(\u2/u11/X [47]),
        .I1(\u2/u11/X [46]),
        .I2(\u2/u11/X [45]),
        .I3(\u2/u11/X [44]),
        .I4(\u2/u11/X [48]),
        .I5(\u2/u11/X [43]),
        .O(\u2/out11 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__347_i_1
       (.I0(\u2/R10_reg_n_0_[32] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [37]),
        .I3(\u2/uk/K_r10 [1]),
        .O(\u2/u11/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__347_i_2
       (.I0(\u2/R10_reg_n_0_[31] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [0]),
        .I3(\u2/uk/K_r10 [50]),
        .O(\u2/u11/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__347_i_3
       (.I0(\u2/R10_reg_n_0_[30] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [43]),
        .I3(\u2/uk/K_r10 [7]),
        .O(\u2/u11/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__347_i_4
       (.I0(\u2/R10_reg_n_0_[29] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [42]),
        .I3(\u2/uk/K_r10 [37]),
        .O(\u2/u11/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__347_i_5
       (.I0(\u2/R10_reg_n_0_[1] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [31]),
        .I3(\u2/uk/K_r10 [22]),
        .O(\u2/u11/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__347_i_6
       (.I0(\u2/R10_reg_n_0_[28] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [15]),
        .I3(\u2/uk/K_r10 [38]),
        .O(\u2/u11/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__348
       (.I0(\u2/u11/X [23]),
        .I1(\u2/u11/X [22]),
        .I2(\u2/u11/X [21]),
        .I3(\u2/u11/X [20]),
        .I4(\u2/u11/X [24]),
        .I5(\u2/u11/X [19]),
        .O(\u2/out11 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__348_i_1
       (.I0(\u2/R10_reg_n_0_[16] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [41]),
        .I3(\u2/uk/K_r10 [32]),
        .O(\u2/u11/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__348_i_2
       (.I0(\u2/R10_reg_n_0_[15] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [33]),
        .I3(\u2/uk/K_r10 [24]),
        .O(\u2/u11/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__348_i_3
       (.I0(\u2/R10_reg_n_0_[14] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [25]),
        .I3(\u2/uk/K_r10 [48]),
        .O(\u2/u11/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__348_i_4
       (.I0(\u2/R10_reg_n_0_[13] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [24]),
        .I3(\u2/uk/K_r10 [47]),
        .O(\u2/u11/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__348_i_5
       (.I0(\u2/R10_reg_n_0_[17] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [46]),
        .I3(\u2/uk/K_r10 [12]),
        .O(\u2/u11/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__348_i_6
       (.I0(\u2/R10_reg_n_0_[12] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [5]),
        .I3(\u2/uk/K_r10 [53]),
        .O(\u2/u11/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__349
       (.I0(\u2/u11/X [29]),
        .I1(\u2/u11/X [28]),
        .I2(\u2/u11/X [27]),
        .I3(\u2/u11/X [26]),
        .I4(\u2/u11/X [30]),
        .I5(\u2/u11/X [25]),
        .O(\u2/out11 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__349_i_1
       (.I0(\u2/R10_reg_n_0_[20] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [22]),
        .I3(\u2/uk/K_r10 [45]),
        .O(\u2/u11/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__349_i_2
       (.I0(\u2/R10_reg_n_0_[19] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [7]),
        .I3(\u2/uk/K_r10 [2]),
        .O(\u2/u11/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__349_i_3
       (.I0(\u2/R10_reg_n_0_[18] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [51]),
        .I3(\u2/uk/K_r10 [15]),
        .O(\u2/u11/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__349_i_4
       (.I0(\u2/R10_reg_n_0_[17] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [2]),
        .I3(\u2/uk/K_r10 [21]),
        .O(\u2/u11/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__349_i_5
       (.I0(\u2/R10_reg_n_0_[21] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [23]),
        .I3(\u2/uk/K_r10 [42]),
        .O(\u2/u11/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__349_i_6
       (.I0(\u2/R10_reg_n_0_[16] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [35]),
        .I3(\u2/uk/K_r10 [30]),
        .O(\u2/u11/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__34_i_1
       (.I0(\u0/R3 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [6]),
        .I3(\u0/uk/K_r3 [40]),
        .O(\u0/u4/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__34_i_2
       (.I0(\u0/R3 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [40]),
        .I3(\u0/uk/K_r3 [17]),
        .O(\u0/u4/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__34_i_3
       (.I0(\u0/R3 [6]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [46]),
        .I3(\u0/uk/K_r3 [55]),
        .O(\u0/u4/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__34_i_4
       (.I0(\u0/R3 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [55]),
        .I3(\u0/uk/K_r3 [32]),
        .O(\u0/u4/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__34_i_5
       (.I0(\u0/R3 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [11]),
        .I3(\u0/uk/K_r3 [20]),
        .O(\u0/u4/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__34_i_6
       (.I0(\u0/R3 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [19]),
        .I3(\u0/uk/K_r3 [53]),
        .O(\u0/u4/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__35
       (.I0(\u0/u4/X [47]),
        .I1(\u0/u4/X [46]),
        .I2(\u0/u4/X [45]),
        .I3(\u0/u4/X [44]),
        .I4(\u0/u4/X [48]),
        .I5(\u0/u4/X [43]),
        .O(\u0/out4 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__350
       (.I0(\u2/u11/X [5]),
        .I1(\u2/u11/X [4]),
        .I2(\u2/u11/X [3]),
        .I3(\u2/u11/X [2]),
        .I4(\u2/u11/X [6]),
        .I5(\u2/u11/X [1]),
        .O(\u2/out11 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__350_i_1
       (.I0(\u2/R10_reg_n_0_[4] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [39]),
        .I3(\u2/uk/K_r10 [5]),
        .O(\u2/u11/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__350_i_2
       (.I0(\u2/R10_reg_n_0_[3] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [4]),
        .I3(\u2/uk/K_r10 [27]),
        .O(\u2/u11/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__350_i_3
       (.I0(\u2/R10_reg_n_0_[2] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [27]),
        .I3(\u2/uk/K_r10 [18]),
        .O(\u2/u11/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__350_i_4
       (.I0(\u2/R10_reg_n_0_[1] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [12]),
        .I3(\u2/uk/K_r10 [3]),
        .O(\u2/u11/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__350_i_5
       (.I0(\u2/R10_reg_n_0_[5] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [10]),
        .I3(\u2/uk/K_r10 [33]),
        .O(\u2/u11/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__350_i_6
       (.I0(\u2/R10_reg_n_0_[32] ),
        .I1(decrypt),
        .I2(\u2/uk/K_r10 [48]),
        .I3(\u2/uk/K_r10 [39]),
        .O(\u2/u11/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__351
       (.I0(\u2/u12/X [41]),
        .I1(\u2/u12/X [40]),
        .I2(\u2/u12/X [39]),
        .I3(\u2/u12/X [38]),
        .I4(\u2/u12/X [42]),
        .I5(\u2/u12/X [37]),
        .O(\u2/out12 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__351_i_1
       (.I0(\u2/R11 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [0]),
        .I3(\u2/uk/K_r11 [22]),
        .O(\u2/u12/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__351_i_2
       (.I0(\u2/R11 [27]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [44]),
        .I3(\u2/uk/K_r11 [35]),
        .O(\u2/u12/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__351_i_3
       (.I0(\u2/R11 [26]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [35]),
        .I3(\u2/uk/K_r11 [2]),
        .O(\u2/u12/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__351_i_4
       (.I0(\u2/R11 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [50]),
        .I3(\u2/uk/K_r11 [45]),
        .O(\u2/u12/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__351_i_5
       (.I0(\u2/R11 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [23]),
        .I3(\u2/uk/K_r11 [14]),
        .O(\u2/u12/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__351_i_6
       (.I0(\u2/R11 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [15]),
        .I3(\u2/uk/K_r11 [37]),
        .O(\u2/u12/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__352
       (.I0(\u2/u12/X [17]),
        .I1(\u2/u12/X [16]),
        .I2(\u2/u12/X [15]),
        .I3(\u2/u12/X [14]),
        .I4(\u2/u12/X [18]),
        .I5(\u2/u12/X [13]),
        .O(\u2/out12 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__352_i_1
       (.I0(\u2/R11 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [32]),
        .I3(\u2/uk/K_r11 [27]),
        .O(\u2/u12/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__352_i_2
       (.I0(\u2/R11 [11]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [17]),
        .I3(\u2/uk/K_r11 [12]),
        .O(\u2/u12/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__352_i_3
       (.I0(\u2/R11 [10]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [48]),
        .I3(\u2/uk/K_r11 [11]),
        .O(\u2/u12/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__352_i_4
       (.I0(\u2/R11 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [40]),
        .I3(\u2/uk/K_r11 [3]),
        .O(\u2/u12/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__352_i_5
       (.I0(\u2/R11 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [20]),
        .I3(\u2/uk/K_r11 [40]),
        .O(\u2/u12/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__352_i_6
       (.I0(\u2/R11 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [11]),
        .I3(\u2/uk/K_r11 [6]),
        .O(\u2/u12/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__353
       (.I0(\u2/u12/X [35]),
        .I1(\u2/u12/X [34]),
        .I2(\u2/u12/X [33]),
        .I3(\u2/u12/X [32]),
        .I4(\u2/u12/X [36]),
        .I5(\u2/u12/X [31]),
        .O(\u2/out12 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__353_i_1
       (.I0(\u2/R11 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [52]),
        .I3(\u2/uk/K_r11 [15]),
        .O(\u2/u12/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__353_i_2
       (.I0(\u2/R11 [23]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [22]),
        .I3(\u2/uk/K_r11 [44]),
        .O(\u2/u12/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__353_i_3
       (.I0(\u2/R11 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [9]),
        .I3(\u2/uk/K_r11 [0]),
        .O(\u2/u12/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__353_i_4
       (.I0(\u2/R11 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [42]),
        .I3(\u2/uk/K_r11 [9]),
        .O(\u2/u12/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__353_i_5
       (.I0(\u2/R11 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [43]),
        .I3(\u2/uk/K_r11 [38]),
        .O(\u2/u12/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__353_i_6
       (.I0(\u2/R11 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [31]),
        .I3(\u2/uk/K_r11 [49]),
        .O(\u2/u12/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__354
       (.I0(\u2/u12/X [11]),
        .I1(\u2/u12/X [10]),
        .I2(\u2/u12/X [9]),
        .I3(\u2/u12/X [8]),
        .I4(\u2/u12/X [12]),
        .I5(\u2/u12/X [7]),
        .O(\u2/out12 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__354_i_1
       (.I0(\u2/R11 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [54]),
        .I3(\u2/uk/K_r11 [17]),
        .O(\u2/u12/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__354_i_2
       (.I0(\u2/R11 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [6]),
        .I3(\u2/uk/K_r11 [26]),
        .O(\u2/u12/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__354_i_3
       (.I0(\u2/R11 [6]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [12]),
        .I3(\u2/uk/K_r11 [32]),
        .O(\u2/u12/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__354_i_4
       (.I0(\u2/R11 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [46]),
        .I3(\u2/uk/K_r11 [41]),
        .O(\u2/u12/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__354_i_5
       (.I0(\u2/R11 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [34]),
        .I3(\u2/uk/K_r11 [54]),
        .O(\u2/u12/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__354_i_6
       (.I0(\u2/R11 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [10]),
        .I3(\u2/uk/K_r11 [5]),
        .O(\u2/u12/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__355
       (.I0(\u2/u12/X [47]),
        .I1(\u2/u12/X [46]),
        .I2(\u2/u12/X [45]),
        .I3(\u2/u12/X [44]),
        .I4(\u2/u12/X [48]),
        .I5(\u2/u12/X [43]),
        .O(\u2/out12 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__355_i_1
       (.I0(\u2/R11 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [51]),
        .I3(\u2/uk/K_r11 [42]),
        .O(\u2/u12/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__355_i_2
       (.I0(\u2/R11 [31]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [14]),
        .I3(\u2/uk/K_r11 [36]),
        .O(\u2/u12/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__355_i_3
       (.I0(\u2/R11 [30]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [2]),
        .I3(\u2/uk/K_r11 [52]),
        .O(\u2/u12/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__355_i_4
       (.I0(\u2/R11 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [1]),
        .I3(\u2/uk/K_r11 [23]),
        .O(\u2/u12/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__355_i_5
       (.I0(\u2/R11 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [45]),
        .I3(\u2/uk/K_r11 [8]),
        .O(\u2/u12/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__355_i_6
       (.I0(\u2/R11 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [29]),
        .I3(\u2/uk/K_r11 [51]),
        .O(\u2/u12/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__356
       (.I0(\u2/u12/X [23]),
        .I1(\u2/u12/X [22]),
        .I2(\u2/u12/X [21]),
        .I3(\u2/u12/X [20]),
        .I4(\u2/u12/X [24]),
        .I5(\u2/u12/X [19]),
        .O(\u2/out12 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__356_i_1
       (.I0(\u2/R11 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [55]),
        .I3(\u2/uk/K_r11 [18]),
        .O(\u2/u12/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__356_i_2
       (.I0(\u2/R11 [15]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [47]),
        .I3(\u2/uk/K_r11 [10]),
        .O(\u2/u12/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__356_i_3
       (.I0(\u2/R11 [14]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [39]),
        .I3(\u2/uk/K_r11 [34]),
        .O(\u2/u12/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__356_i_4
       (.I0(\u2/R11 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [13]),
        .I3(\u2/uk/K_r11 [33]),
        .O(\u2/u12/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__356_i_5
       (.I0(\u2/R11 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [3]),
        .I3(\u2/uk/K_r11 [55]),
        .O(\u2/u12/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__356_i_6
       (.I0(\u2/R11 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [19]),
        .I3(\u2/uk/K_r11 [39]),
        .O(\u2/u12/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__357
       (.I0(\u2/u12/X [29]),
        .I1(\u2/u12/X [28]),
        .I2(\u2/u12/X [27]),
        .I3(\u2/u12/X [26]),
        .I4(\u2/u12/X [30]),
        .I5(\u2/u12/X [25]),
        .O(\u2/out12 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__357_i_1
       (.I0(\u2/R11 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [36]),
        .I3(\u2/uk/K_r11 [31]),
        .O(\u2/u12/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__357_i_2
       (.I0(\u2/R11 [19]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [21]),
        .I3(\u2/uk/K_r11 [43]),
        .O(\u2/u12/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__357_i_3
       (.I0(\u2/R11 [18]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [38]),
        .I3(\u2/uk/K_r11 [1]),
        .O(\u2/u12/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__357_i_4
       (.I0(\u2/R11 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [16]),
        .I3(\u2/uk/K_r11 [7]),
        .O(\u2/u12/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__357_i_5
       (.I0(\u2/R11 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [37]),
        .I3(\u2/uk/K_r11 [28]),
        .O(\u2/u12/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__357_i_6
       (.I0(\u2/R11 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [49]),
        .I3(\u2/uk/K_r11 [16]),
        .O(\u2/u12/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__358
       (.I0(\u2/u12/X [5]),
        .I1(\u2/u12/X [4]),
        .I2(\u2/u12/X [3]),
        .I3(\u2/u12/X [2]),
        .I4(\u2/u12/X [6]),
        .I5(\u2/u12/X [1]),
        .O(\u2/out12 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__358_i_1
       (.I0(\u2/R11 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [53]),
        .I3(\u2/uk/K_r11 [48]),
        .O(\u2/u12/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__358_i_2
       (.I0(\u2/R11 [3]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [18]),
        .I3(\u2/uk/K_r11 [13]),
        .O(\u2/u12/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__358_i_3
       (.I0(\u2/R11 [2]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [41]),
        .I3(\u2/uk/K_r11 [4]),
        .O(\u2/u12/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__358_i_4
       (.I0(\u2/R11 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [26]),
        .I3(\u2/uk/K_r11 [46]),
        .O(\u2/u12/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__358_i_5
       (.I0(\u2/R11 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [24]),
        .I3(\u2/uk/K_r11 [19]),
        .O(\u2/u12/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__358_i_6
       (.I0(\u2/R11 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r11 [5]),
        .I3(\u2/uk/K_r11 [25]),
        .O(\u2/u12/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__359
       (.I0(\u2/u13/X [41]),
        .I1(\u2/u13/X [40]),
        .I2(\u2/u13/X [39]),
        .I3(\u2/u13/X [38]),
        .I4(\u2/u13/X [42]),
        .I5(\u2/u13/X [37]),
        .O(\u2/out13 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__359_i_1
       (.I0(\u2/R12 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [14]),
        .I3(\u2/uk/K_r12 [8]),
        .O(\u2/u13/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__359_i_2
       (.I0(\u2/R12 [27]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [31]),
        .I3(\u2/uk/K_r12 [21]),
        .O(\u2/u13/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__359_i_3
       (.I0(\u2/R12 [26]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [49]),
        .I3(\u2/uk/K_r12 [43]),
        .O(\u2/u13/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__359_i_4
       (.I0(\u2/R12 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [9]),
        .I3(\u2/uk/K_r12 [31]),
        .O(\u2/u13/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__359_i_5
       (.I0(\u2/R12 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [37]),
        .I3(\u2/uk/K_r12 [0]),
        .O(\u2/u13/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__359_i_6
       (.I0(\u2/R12 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [29]),
        .I3(\u2/uk/K_r12 [23]),
        .O(\u2/u13/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__35_i_1
       (.I0(\u0/R3 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [1]),
        .I3(\u0/uk/K_r3 [37]),
        .O(\u0/u4/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__35_i_2
       (.I0(\u0/R3 [31]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [50]),
        .I3(\u0/uk/K_r3 [0]),
        .O(\u0/u4/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__35_i_3
       (.I0(\u0/R3 [30]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [7]),
        .I3(\u0/uk/K_r3 [43]),
        .O(\u0/u4/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__35_i_4
       (.I0(\u0/R3 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [37]),
        .I3(\u0/uk/K_r3 [42]),
        .O(\u0/u4/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__35_i_5
       (.I0(\u0/R3 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [22]),
        .I3(\u0/uk/K_r3 [31]),
        .O(\u0/u4/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__35_i_6
       (.I0(\u0/R3 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [38]),
        .I3(\u0/uk/K_r3 [15]),
        .O(\u0/u4/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__36
       (.I0(\u0/u4/X [23]),
        .I1(\u0/u4/X [22]),
        .I2(\u0/u4/X [21]),
        .I3(\u0/u4/X [20]),
        .I4(\u0/u4/X [24]),
        .I5(\u0/u4/X [19]),
        .O(\u0/out4 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__360
       (.I0(\u2/u13/X [17]),
        .I1(\u2/u13/X [16]),
        .I2(\u2/u13/X [15]),
        .I3(\u2/u13/X [14]),
        .I4(\u2/u13/X [18]),
        .I5(\u2/u13/X [13]),
        .O(\u2/out13 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__360_i_1
       (.I0(\u2/R12 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [46]),
        .I3(\u2/uk/K_r12 [13]),
        .O(\u2/u13/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__360_i_2
       (.I0(\u2/R12 [11]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [6]),
        .I3(\u2/uk/K_r12 [55]),
        .O(\u2/u13/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__360_i_3
       (.I0(\u2/R12 [10]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [5]),
        .I3(\u2/uk/K_r12 [54]),
        .O(\u2/u13/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__360_i_4
       (.I0(\u2/R12 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [54]),
        .I3(\u2/uk/K_r12 [46]),
        .O(\u2/u13/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__360_i_5
       (.I0(\u2/R12 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [34]),
        .I3(\u2/uk/K_r12 [26]),
        .O(\u2/u13/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__360_i_6
       (.I0(\u2/R12 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [25]),
        .I3(\u2/uk/K_r12 [17]),
        .O(\u2/u13/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__361
       (.I0(\u2/u13/X [35]),
        .I1(\u2/u13/X [34]),
        .I2(\u2/u13/X [33]),
        .I3(\u2/u13/X [32]),
        .I4(\u2/u13/X [36]),
        .I5(\u2/u13/X [31]),
        .O(\u2/out13 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__361_i_1
       (.I0(\u2/R12 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [7]),
        .I3(\u2/uk/K_r12 [1]),
        .O(\u2/u13/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__361_i_2
       (.I0(\u2/R12 [23]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [36]),
        .I3(\u2/uk/K_r12 [30]),
        .O(\u2/u13/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__361_i_3
       (.I0(\u2/R12 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [23]),
        .I3(\u2/uk/K_r12 [45]),
        .O(\u2/u13/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__361_i_4
       (.I0(\u2/R12 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [1]),
        .I3(\u2/uk/K_r12 [50]),
        .O(\u2/u13/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__361_i_5
       (.I0(\u2/R12 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [2]),
        .I3(\u2/uk/K_r12 [51]),
        .O(\u2/u13/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__361_i_6
       (.I0(\u2/R12 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [45]),
        .I3(\u2/uk/K_r12 [35]),
        .O(\u2/u13/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__362
       (.I0(\u2/u13/X [11]),
        .I1(\u2/u13/X [10]),
        .I2(\u2/u13/X [9]),
        .I3(\u2/u13/X [8]),
        .I4(\u2/u13/X [12]),
        .I5(\u2/u13/X [7]),
        .O(\u2/out13 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__362_i_1
       (.I0(\u2/R12 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [11]),
        .I3(\u2/uk/K_r12 [3]),
        .O(\u2/u13/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__362_i_2
       (.I0(\u2/R12 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [20]),
        .I3(\u2/uk/K_r12 [12]),
        .O(\u2/u13/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__362_i_3
       (.I0(\u2/R12 [6]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [26]),
        .I3(\u2/uk/K_r12 [18]),
        .O(\u2/u13/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__362_i_4
       (.I0(\u2/R12 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [3]),
        .I3(\u2/uk/K_r12 [27]),
        .O(\u2/u13/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__362_i_5
       (.I0(\u2/R12 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [48]),
        .I3(\u2/uk/K_r12 [40]),
        .O(\u2/u13/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__362_i_6
       (.I0(\u2/R12 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [24]),
        .I3(\u2/uk/K_r12 [48]),
        .O(\u2/u13/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__363
       (.I0(\u2/u13/X [47]),
        .I1(\u2/u13/X [46]),
        .I2(\u2/u13/X [45]),
        .I3(\u2/u13/X [44]),
        .I4(\u2/u13/X [48]),
        .I5(\u2/u13/X [43]),
        .O(\u2/out13 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__363_i_1
       (.I0(\u2/R12 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [38]),
        .I3(\u2/uk/K_r12 [28]),
        .O(\u2/u13/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__363_i_2
       (.I0(\u2/R12 [31]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [28]),
        .I3(\u2/uk/K_r12 [22]),
        .O(\u2/u13/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__363_i_3
       (.I0(\u2/R12 [30]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [16]),
        .I3(\u2/uk/K_r12 [38]),
        .O(\u2/u13/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__363_i_4
       (.I0(\u2/R12 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [15]),
        .I3(\u2/uk/K_r12 [9]),
        .O(\u2/u13/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__363_i_5
       (.I0(\u2/R12 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [0]),
        .I3(\u2/uk/K_r12 [49]),
        .O(\u2/u13/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__363_i_6
       (.I0(\u2/R12 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [43]),
        .I3(\u2/uk/K_r12 [37]),
        .O(\u2/u13/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__364
       (.I0(\u2/u13/X [23]),
        .I1(\u2/u13/X [22]),
        .I2(\u2/u13/X [21]),
        .I3(\u2/u13/X [20]),
        .I4(\u2/u13/X [24]),
        .I5(\u2/u13/X [19]),
        .O(\u2/out13 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__364_i_1
       (.I0(\u2/R12 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [12]),
        .I3(\u2/uk/K_r12 [4]),
        .O(\u2/u13/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__364_i_2
       (.I0(\u2/R12 [15]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [4]),
        .I3(\u2/uk/K_r12 [53]),
        .O(\u2/u13/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__364_i_3
       (.I0(\u2/R12 [14]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [53]),
        .I3(\u2/uk/K_r12 [20]),
        .O(\u2/u13/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__364_i_4
       (.I0(\u2/R12 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [27]),
        .I3(\u2/uk/K_r12 [19]),
        .O(\u2/u13/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__364_i_5
       (.I0(\u2/R12 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [17]),
        .I3(\u2/uk/K_r12 [41]),
        .O(\u2/u13/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__364_i_6
       (.I0(\u2/R12 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [33]),
        .I3(\u2/uk/K_r12 [25]),
        .O(\u2/u13/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__365
       (.I0(\u2/u13/X [29]),
        .I1(\u2/u13/X [28]),
        .I2(\u2/u13/X [27]),
        .I3(\u2/u13/X [26]),
        .I4(\u2/u13/X [30]),
        .I5(\u2/u13/X [25]),
        .O(\u2/out13 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__365_i_1
       (.I0(\u2/R12 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [50]),
        .I3(\u2/uk/K_r12 [44]),
        .O(\u2/u13/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__365_i_2
       (.I0(\u2/R12 [19]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [35]),
        .I3(\u2/uk/K_r12 [29]),
        .O(\u2/u13/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__365_i_3
       (.I0(\u2/R12 [18]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [52]),
        .I3(\u2/uk/K_r12 [42]),
        .O(\u2/u13/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__365_i_4
       (.I0(\u2/R12 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [30]),
        .I3(\u2/uk/K_r12 [52]),
        .O(\u2/u13/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__365_i_5
       (.I0(\u2/R12 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [51]),
        .I3(\u2/uk/K_r12 [14]),
        .O(\u2/u13/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__365_i_6
       (.I0(\u2/R12 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [8]),
        .I3(\u2/uk/K_r12 [2]),
        .O(\u2/u13/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__366
       (.I0(\u2/u13/X [5]),
        .I1(\u2/u13/X [4]),
        .I2(\u2/u13/X [3]),
        .I3(\u2/u13/X [2]),
        .I4(\u2/u13/X [6]),
        .I5(\u2/u13/X [1]),
        .O(\u2/out13 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__366_i_1
       (.I0(\u2/R12 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [10]),
        .I3(\u2/uk/K_r12 [34]),
        .O(\u2/u13/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__366_i_2
       (.I0(\u2/R12 [3]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [32]),
        .I3(\u2/uk/K_r12 [24]),
        .O(\u2/u13/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__366_i_3
       (.I0(\u2/R12 [2]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [55]),
        .I3(\u2/uk/K_r12 [47]),
        .O(\u2/u13/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__366_i_4
       (.I0(\u2/R12 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [40]),
        .I3(\u2/uk/K_r12 [32]),
        .O(\u2/u13/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__366_i_5
       (.I0(\u2/R12 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [13]),
        .I3(\u2/uk/K_r12 [5]),
        .O(\u2/u13/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__366_i_6
       (.I0(\u2/R12 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r12 [19]),
        .I3(\u2/uk/K_r12 [11]),
        .O(\u2/u13/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__367
       (.I0(\u2/u14/X [41]),
        .I1(\u2/u14/X [40]),
        .I2(\u2/u14/X [39]),
        .I3(\u2/u14/X [38]),
        .I4(\u2/u14/X [42]),
        .I5(\u2/u14/X [37]),
        .O(\u2/out14 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__367_i_1
       (.I0(\u2/R13 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [28]),
        .I3(\u2/uk/K_r13 [49]),
        .O(\u2/u14/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__367_i_2
       (.I0(\u2/R13 [27]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [45]),
        .I3(\u2/uk/K_r13 [7]),
        .O(\u2/u14/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__367_i_3
       (.I0(\u2/R13 [26]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [8]),
        .I3(\u2/uk/K_r13 [29]),
        .O(\u2/u14/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__367_i_4
       (.I0(\u2/R13 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [23]),
        .I3(\u2/uk/K_r13 [44]),
        .O(\u2/u14/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__367_i_5
       (.I0(\u2/R13 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [51]),
        .I3(\u2/uk/K_r13 [45]),
        .O(\u2/u14/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__367_i_6
       (.I0(\u2/R13 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [43]),
        .I3(\u2/uk/K_r13 [9]),
        .O(\u2/u14/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__368
       (.I0(\u2/u14/X [17]),
        .I1(\u2/u14/X [16]),
        .I2(\u2/u14/X [15]),
        .I3(\u2/u14/X [14]),
        .I4(\u2/u14/X [18]),
        .I5(\u2/u14/X [13]),
        .O(\u2/out14 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__368_i_1
       (.I0(\u2/R13 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [3]),
        .I3(\u2/uk/K_r13 [24]),
        .O(\u2/u14/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__368_i_2
       (.I0(\u2/R13 [11]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [20]),
        .I3(\u2/uk/K_r13 [41]),
        .O(\u2/u14/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__368_i_3
       (.I0(\u2/R13 [10]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [19]),
        .I3(\u2/uk/K_r13 [40]),
        .O(\u2/u14/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__368_i_4
       (.I0(\u2/R13 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [11]),
        .I3(\u2/uk/K_r13 [32]),
        .O(\u2/u14/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__368_i_5
       (.I0(\u2/R13 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [48]),
        .I3(\u2/uk/K_r13 [12]),
        .O(\u2/u14/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__368_i_6
       (.I0(\u2/R13 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [39]),
        .I3(\u2/uk/K_r13 [3]),
        .O(\u2/u14/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__369
       (.I0(\u2/u14/X [35]),
        .I1(\u2/u14/X [34]),
        .I2(\u2/u14/X [33]),
        .I3(\u2/u14/X [32]),
        .I4(\u2/u14/X [36]),
        .I5(\u2/u14/X [31]),
        .O(\u2/out14 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__369_i_1
       (.I0(\u2/R13 [24]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [21]),
        .I3(\u2/uk/K_r13 [42]),
        .O(\u2/u14/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__369_i_2
       (.I0(\u2/R13 [23]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [50]),
        .I3(\u2/uk/K_r13 [16]),
        .O(\u2/u14/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__369_i_3
       (.I0(\u2/R13 [22]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [37]),
        .I3(\u2/uk/K_r13 [31]),
        .O(\u2/u14/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__369_i_4
       (.I0(\u2/R13 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [15]),
        .I3(\u2/uk/K_r13 [36]),
        .O(\u2/u14/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__369_i_5
       (.I0(\u2/R13 [25]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [16]),
        .I3(\u2/uk/K_r13 [37]),
        .O(\u2/u14/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__369_i_6
       (.I0(\u2/R13 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [0]),
        .I3(\u2/uk/K_r13 [21]),
        .O(\u2/u14/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__36_i_1
       (.I0(\u0/R3 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [32]),
        .I3(\u0/uk/K_r3 [41]),
        .O(\u0/u4/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__36_i_2
       (.I0(\u0/R3 [15]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [24]),
        .I3(\u0/uk/K_r3 [33]),
        .O(\u0/u4/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__36_i_3
       (.I0(\u0/R3 [14]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [48]),
        .I3(\u0/uk/K_r3 [25]),
        .O(\u0/u4/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__36_i_4
       (.I0(\u0/R3 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [47]),
        .I3(\u0/uk/K_r3 [24]),
        .O(\u0/u4/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__36_i_5
       (.I0(\u0/R3 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [12]),
        .I3(\u0/uk/K_r3 [46]),
        .O(\u0/u4/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__36_i_6
       (.I0(\u0/R3 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [53]),
        .I3(\u0/uk/K_r3 [5]),
        .O(\u0/u4/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__37
       (.I0(\u0/u4/X [29]),
        .I1(\u0/u4/X [28]),
        .I2(\u0/u4/X [27]),
        .I3(\u0/u4/X [26]),
        .I4(\u0/u4/X [30]),
        .I5(\u0/u4/X [25]),
        .O(\u0/out4 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__370
       (.I0(\u2/u14/X [11]),
        .I1(\u2/u14/X [10]),
        .I2(\u2/u14/X [9]),
        .I3(\u2/u14/X [8]),
        .I4(\u2/u14/X [12]),
        .I5(\u2/u14/X [7]),
        .O(\u2/out14 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__370_i_1
       (.I0(\u2/R13 [8]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [25]),
        .I3(\u2/uk/K_r13 [46]),
        .O(\u2/u14/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__370_i_2
       (.I0(\u2/R13 [7]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [34]),
        .I3(\u2/uk/K_r13 [55]),
        .O(\u2/u14/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__370_i_3
       (.I0(\u2/R13 [6]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [40]),
        .I3(\u2/uk/K_r13 [4]),
        .O(\u2/u14/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__370_i_4
       (.I0(\u2/R13 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [17]),
        .I3(\u2/uk/K_r13 [13]),
        .O(\u2/u14/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__370_i_5
       (.I0(\u2/R13 [9]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [5]),
        .I3(\u2/uk/K_r13 [26]),
        .O(\u2/u14/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__370_i_6
       (.I0(\u2/R13 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [13]),
        .I3(\u2/uk/K_r13 [34]),
        .O(\u2/u14/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__371
       (.I0(\u2/u14/X [47]),
        .I1(\u2/u14/X [46]),
        .I2(\u2/u14/X [45]),
        .I3(\u2/u14/X [44]),
        .I4(\u2/u14/X [48]),
        .I5(\u2/u14/X [43]),
        .O(\u2/out14 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__371_i_1
       (.I0(\u2/R13 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [52]),
        .I3(\u2/uk/K_r13 [14]),
        .O(\u2/u14/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__371_i_2
       (.I0(\u2/R13 [31]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [42]),
        .I3(\u2/uk/K_r13 [8]),
        .O(\u2/u14/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__371_i_3
       (.I0(\u2/R13 [30]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [30]),
        .I3(\u2/uk/K_r13 [51]),
        .O(\u2/u14/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__371_i_4
       (.I0(\u2/R13 [29]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [29]),
        .I3(\u2/uk/K_r13 [50]),
        .O(\u2/u14/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__371_i_5
       (.I0(\u2/R13 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [14]),
        .I3(\u2/uk/K_r13 [35]),
        .O(\u2/u14/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__371_i_6
       (.I0(\u2/R13 [28]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [2]),
        .I3(\u2/uk/K_r13 [23]),
        .O(\u2/u14/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__372
       (.I0(\u2/u14/X [23]),
        .I1(\u2/u14/X [22]),
        .I2(\u2/u14/X [21]),
        .I3(\u2/u14/X [20]),
        .I4(\u2/u14/X [24]),
        .I5(\u2/u14/X [19]),
        .O(\u2/out14 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__372_i_1
       (.I0(\u2/R13 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [26]),
        .I3(\u2/uk/K_r13 [47]),
        .O(\u2/u14/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__372_i_2
       (.I0(\u2/R13 [15]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [18]),
        .I3(\u2/uk/K_r13 [39]),
        .O(\u2/u14/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__372_i_3
       (.I0(\u2/R13 [14]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [10]),
        .I3(\u2/uk/K_r13 [6]),
        .O(\u2/u14/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__372_i_4
       (.I0(\u2/R13 [13]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [41]),
        .I3(\u2/uk/K_r13 [5]),
        .O(\u2/u14/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__372_i_5
       (.I0(\u2/R13 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [6]),
        .I3(\u2/uk/K_r13 [27]),
        .O(\u2/u14/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__372_i_6
       (.I0(\u2/R13 [12]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [47]),
        .I3(\u2/uk/K_r13 [11]),
        .O(\u2/u14/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__373
       (.I0(\u2/u14/X [29]),
        .I1(\u2/u14/X [28]),
        .I2(\u2/u14/X [27]),
        .I3(\u2/u14/X [26]),
        .I4(\u2/u14/X [30]),
        .I5(\u2/u14/X [25]),
        .O(\u2/out14 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__373_i_1
       (.I0(\u2/R13 [20]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [9]),
        .I3(\u2/uk/K_r13 [30]),
        .O(\u2/u14/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__373_i_2
       (.I0(\u2/R13 [19]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [49]),
        .I3(\u2/uk/K_r13 [15]),
        .O(\u2/u14/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__373_i_3
       (.I0(\u2/R13 [18]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [7]),
        .I3(\u2/uk/K_r13 [28]),
        .O(\u2/u14/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__373_i_4
       (.I0(\u2/R13 [17]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [44]),
        .I3(\u2/uk/K_r13 [38]),
        .O(\u2/u14/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__373_i_5
       (.I0(\u2/R13 [21]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [38]),
        .I3(\u2/uk/K_r13 [0]),
        .O(\u2/u14/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__373_i_6
       (.I0(\u2/R13 [16]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [22]),
        .I3(\u2/uk/K_r13 [43]),
        .O(\u2/u14/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__374
       (.I0(\u2/u14/X [5]),
        .I1(\u2/u14/X [4]),
        .I2(\u2/u14/X [3]),
        .I3(\u2/u14/X [2]),
        .I4(\u2/u14/X [6]),
        .I5(\u2/u14/X [1]),
        .O(\u2/out14 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__374_i_1
       (.I0(\u2/R13 [4]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [24]),
        .I3(\u2/uk/K_r13 [20]),
        .O(\u2/u14/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__374_i_2
       (.I0(\u2/R13 [3]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [46]),
        .I3(\u2/uk/K_r13 [10]),
        .O(\u2/u14/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__374_i_3
       (.I0(\u2/R13 [2]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [12]),
        .I3(\u2/uk/K_r13 [33]),
        .O(\u2/u14/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__374_i_4
       (.I0(\u2/R13 [1]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [54]),
        .I3(\u2/uk/K_r13 [18]),
        .O(\u2/u14/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__374_i_5
       (.I0(\u2/R13 [5]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [27]),
        .I3(\u2/uk/K_r13 [48]),
        .O(\u2/u14/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__374_i_6
       (.I0(\u2/R13 [32]),
        .I1(decrypt),
        .I2(\u2/uk/K_r13 [33]),
        .I3(\u2/uk/K_r13 [54]),
        .O(\u2/u14/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__375
       (.I0(\u2/u15/X [41]),
        .I1(\u2/u15/X [40]),
        .I2(\u2/u15/X [39]),
        .I3(\u2/u15/X [38]),
        .I4(\u2/u15/X [42]),
        .I5(\u2/u15/X [37]),
        .O(\u2/out15 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__375_i_1
       (.I0(\u2/FP [60]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[35] ),
        .I3(\u2/uk/K_r14_reg_n_0_[42] ),
        .O(\u2/u15/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__375_i_2
       (.I0(\u2/FP [59]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[52] ),
        .I3(\u2/uk/K_r14_reg_n_0_ ),
        .O(\u2/u15/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__375_i_3
       (.I0(\u2/FP [58]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[15] ),
        .I3(\u2/uk/K_r14_reg_n_0_[22] ),
        .O(\u2/u15/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__375_i_4
       (.I0(\u2/FP [57]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[30] ),
        .I3(\u2/uk/K_r14_reg_n_0_[37] ),
        .O(\u2/u15/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__375_i_5
       (.I0(\u2/FP [61]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[31] ),
        .I3(\u2/uk/K_r14_reg_n_0_[38] ),
        .O(\u2/u15/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__375_i_6
       (.I0(\u2/FP [56]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[50] ),
        .I3(\u2/uk/K_r14_reg_n_0_[2] ),
        .O(\u2/u15/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__376
       (.I0(\u2/u15/X [17]),
        .I1(\u2/u15/X [16]),
        .I2(\u2/u15/X [15]),
        .I3(\u2/u15/X [14]),
        .I4(\u2/u15/X [18]),
        .I5(\u2/u15/X [13]),
        .O(\u2/out15 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__376_i_1
       (.I0(\u2/FP [44]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[10] ),
        .I3(\u2/uk/K_r14_reg_n_0_[17] ),
        .O(\u2/u15/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__376_i_2
       (.I0(\u2/FP [43]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[27] ),
        .I3(\u2/uk/K_r14_reg_n_0_[34] ),
        .O(\u2/u15/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__376_i_3
       (.I0(\u2/FP [42]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[26] ),
        .I3(\u2/uk/K_r14_reg_n_0_[33] ),
        .O(\u2/u15/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__376_i_4
       (.I0(\u2/FP [41]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[18] ),
        .I3(\u2/uk/K_r14_reg_n_0_[25] ),
        .O(\u2/u15/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__376_i_5
       (.I0(\u2/FP [45]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[55] ),
        .I3(\u2/uk/K_r14_reg_n_0_[5] ),
        .O(\u2/u15/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__376_i_6
       (.I0(\u2/FP [40]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[46] ),
        .I3(\u2/uk/K_r14_reg_n_0_[53] ),
        .O(\u2/u15/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__377
       (.I0(\u2/u15/X [35]),
        .I1(\u2/u15/X [34]),
        .I2(\u2/u15/X [33]),
        .I3(\u2/u15/X [32]),
        .I4(\u2/u15/X [36]),
        .I5(\u2/u15/X [31]),
        .O(\u2/out15 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__377_i_1
       (.I0(\u2/FP [56]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[28] ),
        .I3(\u2/uk/K_r14_reg_n_0_[35] ),
        .O(\u2/u15/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__377_i_2
       (.I0(\u2/FP [55]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[2] ),
        .I3(\u2/uk/K_r14_reg_n_0_[9] ),
        .O(\u2/u15/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__377_i_3
       (.I0(\u2/FP [54]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[44] ),
        .I3(\u2/uk/K_r14_reg_n_0_[51] ),
        .O(\u2/u15/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__377_i_4
       (.I0(\u2/FP [53]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[22] ),
        .I3(\u2/uk/K_r14_reg_n_0_[29] ),
        .O(\u2/u15/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__377_i_5
       (.I0(\u2/FP [57]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[23] ),
        .I3(\u2/uk/K_r14_reg_n_0_[30] ),
        .O(\u2/u15/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__377_i_6
       (.I0(\u2/FP [52]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[7] ),
        .I3(\u2/uk/K_r14_reg_n_0_[14] ),
        .O(\u2/u15/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__378
       (.I0(\u2/u15/X [11]),
        .I1(\u2/u15/X [10]),
        .I2(\u2/u15/X [9]),
        .I3(\u2/u15/X [8]),
        .I4(\u2/u15/X [12]),
        .I5(\u2/u15/X [7]),
        .O(\u2/out15 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__378_i_1
       (.I0(\u2/FP [40]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[32] ),
        .I3(\u2/uk/K_r14_reg_n_0_[39] ),
        .O(\u2/u15/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__378_i_2
       (.I0(\u2/FP [39]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[41] ),
        .I3(\u2/uk/K_r14_reg_n_0_[48] ),
        .O(\u2/u15/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__378_i_3
       (.I0(\u2/FP [38]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[47] ),
        .I3(\u2/uk/K_r14_reg_n_0_[54] ),
        .O(\u2/u15/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__378_i_4
       (.I0(\u2/FP [37]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[24] ),
        .I3(\u2/uk/K_r14_reg_n_0_[6] ),
        .O(\u2/u15/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__378_i_5
       (.I0(\u2/FP [41]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[12] ),
        .I3(\u2/uk/K_r14_reg_n_0_[19] ),
        .O(\u2/u15/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__378_i_6
       (.I0(\u2/FP [36]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[20] ),
        .I3(\u2/uk/K_r14_reg_n_0_[27] ),
        .O(\u2/u15/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__379
       (.I0(\u2/u15/X [47]),
        .I1(\u2/u15/X [46]),
        .I2(\u2/u15/X [45]),
        .I3(\u2/u15/X [44]),
        .I4(\u2/u15/X [48]),
        .I5(\u2/u15/X [43]),
        .O(\u2/out15 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__379_i_1
       (.I0(\u2/FP [64]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_ ),
        .I3(\u2/uk/K_r14_reg_n_0_[7] ),
        .O(\u2/u15/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__379_i_2
       (.I0(\u2/FP [63]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[49] ),
        .I3(\u2/uk/K_r14_reg_n_0_[1] ),
        .O(\u2/u15/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__379_i_3
       (.I0(\u2/FP [62]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[37] ),
        .I3(\u2/uk/K_r14_reg_n_0_[44] ),
        .O(\u2/u15/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__379_i_4
       (.I0(\u2/FP [61]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[36] ),
        .I3(\u2/uk/K_r14_reg_n_0_[43] ),
        .O(\u2/u15/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__379_i_5
       (.I0(\u2/FP [33]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[21] ),
        .I3(\u2/uk/K_r14_reg_n_0_[28] ),
        .O(\u2/u15/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__379_i_6
       (.I0(\u2/FP [60]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[9] ),
        .I3(\u2/uk/K_r14_reg_n_0_[16] ),
        .O(\u2/u15/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__37_i_1
       (.I0(\u0/R3 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [45]),
        .I3(\u0/uk/K_r3 [22]),
        .O(\u0/u4/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__37_i_2
       (.I0(\u0/R3 [19]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [2]),
        .I3(\u0/uk/K_r3 [7]),
        .O(\u0/u4/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__37_i_3
       (.I0(\u0/R3 [18]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [15]),
        .I3(\u0/uk/K_r3 [51]),
        .O(\u0/u4/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__37_i_4
       (.I0(\u0/R3 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [21]),
        .I3(\u0/uk/K_r3 [2]),
        .O(\u0/u4/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__37_i_5
       (.I0(\u0/R3 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [42]),
        .I3(\u0/uk/K_r3 [23]),
        .O(\u0/u4/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__37_i_6
       (.I0(\u0/R3 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [30]),
        .I3(\u0/uk/K_r3 [35]),
        .O(\u0/u4/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__38
       (.I0(\u0/u4/X [5]),
        .I1(\u0/u4/X [4]),
        .I2(\u0/u4/X [3]),
        .I3(\u0/u4/X [2]),
        .I4(\u0/u4/X [6]),
        .I5(\u0/u4/X [1]),
        .O(\u0/out4 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__380
       (.I0(\u2/u15/X [23]),
        .I1(\u2/u15/X [22]),
        .I2(\u2/u15/X [21]),
        .I3(\u2/u15/X [20]),
        .I4(\u2/u15/X [24]),
        .I5(\u2/u15/X [19]),
        .O(\u2/out15 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__380_i_1
       (.I0(\u2/FP [48]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[33] ),
        .I3(\u2/uk/K_r14_reg_n_0_[40] ),
        .O(\u2/u15/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__380_i_2
       (.I0(\u2/FP [47]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[25] ),
        .I3(\u2/uk/K_r14_reg_n_0_[32] ),
        .O(\u2/u15/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__380_i_3
       (.I0(\u2/FP [46]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[17] ),
        .I3(\u2/uk/K_r14_reg_n_0_[24] ),
        .O(\u2/u15/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__380_i_4
       (.I0(\u2/FP [45]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[48] ),
        .I3(\u2/uk/K_r14_reg_n_0_[55] ),
        .O(\u2/u15/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__380_i_5
       (.I0(\u2/FP [49]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[13] ),
        .I3(\u2/uk/K_r14_reg_n_0_[20] ),
        .O(\u2/u15/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__380_i_6
       (.I0(\u2/FP [44]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[54] ),
        .I3(\u2/uk/K_r14_reg_n_0_[4] ),
        .O(\u2/u15/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__381
       (.I0(\u2/u15/X [29]),
        .I1(\u2/u15/X [28]),
        .I2(\u2/u15/X [27]),
        .I3(\u2/u15/X [26]),
        .I4(\u2/u15/X [30]),
        .I5(\u2/u15/X [25]),
        .O(\u2/out15 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__381_i_1
       (.I0(\u2/FP [52]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[16] ),
        .I3(\u2/uk/K_r14_reg_n_0_[23] ),
        .O(\u2/u15/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__381_i_2
       (.I0(\u2/FP [51]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[1] ),
        .I3(\u2/uk/K_r14_reg_n_0_[8] ),
        .O(\u2/u15/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__381_i_3
       (.I0(\u2/FP [50]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[14] ),
        .I3(\u2/uk/K_r14_reg_n_0_[21] ),
        .O(\u2/u15/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__381_i_4
       (.I0(\u2/FP [49]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[51] ),
        .I3(\u2/uk/K_r14_reg_n_0_[31] ),
        .O(\u2/u15/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__381_i_5
       (.I0(\u2/FP [53]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[45] ),
        .I3(\u2/uk/K_r14_reg_n_0_[52] ),
        .O(\u2/u15/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__381_i_6
       (.I0(\u2/FP [48]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[29] ),
        .I3(\u2/uk/K_r14_reg_n_0_[36] ),
        .O(\u2/u15/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__382
       (.I0(\u2/u15/X [5]),
        .I1(\u2/u15/X [4]),
        .I2(\u2/u15/X [3]),
        .I3(\u2/u15/X [2]),
        .I4(\u2/u15/X [6]),
        .I5(\u2/u15/X [1]),
        .O(\u2/out15 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__382_i_1
       (.I0(\u2/FP [36]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[6] ),
        .I3(\u2/uk/K_r14_reg_n_0_[13] ),
        .O(\u2/u15/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__382_i_2
       (.I0(\u2/FP [35]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[53] ),
        .I3(\u2/uk/K_r14_reg_n_0_[3] ),
        .O(\u2/u15/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__382_i_3
       (.I0(\u2/FP [34]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[19] ),
        .I3(\u2/uk/K_r14_reg_n_0_[26] ),
        .O(\u2/u15/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__382_i_4
       (.I0(\u2/FP [33]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[4] ),
        .I3(\u2/uk/K_r14_reg_n_0_[11] ),
        .O(\u2/u15/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__382_i_5
       (.I0(\u2/FP [37]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[34] ),
        .I3(\u2/uk/K_r14_reg_n_0_[41] ),
        .O(\u2/u15/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__382_i_6
       (.I0(\u2/FP [64]),
        .I1(decrypt),
        .I2(\u2/uk/K_r14_reg_n_0_[40] ),
        .I3(\u2/uk/K_r14_reg_n_0_[47] ),
        .O(\u2/u15/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__38_i_1
       (.I0(\u0/R3 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [5]),
        .I3(\u0/uk/K_r3 [39]),
        .O(\u0/u4/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__38_i_2
       (.I0(\u0/R3 [3]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [27]),
        .I3(\u0/uk/K_r3 [4]),
        .O(\u0/u4/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__38_i_3
       (.I0(\u0/R3 [2]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [18]),
        .I3(\u0/uk/K_r3 [27]),
        .O(\u0/u4/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__38_i_4
       (.I0(\u0/R3 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [3]),
        .I3(\u0/uk/K_r3 [12]),
        .O(\u0/u4/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__38_i_5
       (.I0(\u0/R3 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [33]),
        .I3(\u0/uk/K_r3 [10]),
        .O(\u0/u4/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__38_i_6
       (.I0(\u0/R3 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r3 [39]),
        .I3(\u0/uk/K_r3 [48]),
        .O(\u0/u4/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__39
       (.I0(\u0/u5/X [41]),
        .I1(\u0/u5/X [40]),
        .I2(\u0/u5/X [39]),
        .I3(\u0/u5/X [38]),
        .I4(\u0/u5/X [42]),
        .I5(\u0/u5/X [37]),
        .O(\u0/out5 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__39_i_1
       (.I0(\u0/R4 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[50] ),
        .I3(\u0/uk/K_r4_reg_n_0_[31] ),
        .O(\u0/u5/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__39_i_2
       (.I0(\u0/R4 [27]),
        .I1(decrypt),
        .I2(\u0/uk/p_42_in ),
        .I3(\u0/uk/K_r4_reg_n_0_[16] ),
        .O(\u0/u5/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__39_i_3
       (.I0(\u0/R4 [26]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[30] ),
        .I3(\u0/uk/K_r4_reg_n_0_[7] ),
        .O(\u0/u5/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__39_i_4
       (.I0(\u0/R4 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[14] ),
        .I3(\u0/uk/K_r4_reg_n_0_[22] ),
        .O(\u0/u5/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__39_i_5
       (.I0(\u0/R4 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[42] ),
        .I3(\u0/uk/K_r4_reg_n_0_[50] ),
        .O(\u0/u5/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__39_i_6
       (.I0(\u0/R4 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[38] ),
        .I3(\u0/uk/K_r4_reg_n_0_[42] ),
        .O(\u0/u5/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__3_i_1
       (.I0(\u0/IP [64]),
        .I1(decrypt),
        .I2(\u0/key_r [7]),
        .I3(\u0/key_r [0]),
        .O(\u0/u0/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__3_i_2
       (.I0(\u0/IP [63]),
        .I1(decrypt),
        .I2(\u0/key_r [1]),
        .I3(\u0/key_r [49]),
        .O(\u0/u0/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__3_i_3
       (.I0(\u0/IP [62]),
        .I1(decrypt),
        .I2(\u0/key_r [44]),
        .I3(\u0/key_r [37]),
        .O(\u0/u0/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__3_i_4
       (.I0(\u0/IP [61]),
        .I1(decrypt),
        .I2(\u0/key_r [43]),
        .I3(\u0/key_r [36]),
        .O(\u0/u0/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__3_i_5
       (.I0(\u0/IP [33]),
        .I1(decrypt),
        .I2(\u0/key_r [28]),
        .I3(\u0/key_r [21]),
        .O(\u0/u0/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__3_i_6
       (.I0(\u0/IP [60]),
        .I1(decrypt),
        .I2(\u0/key_r [16]),
        .I3(\u0/key_r [9]),
        .O(\u0/u0/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__4
       (.I0(\u0/u0/X [23]),
        .I1(\u0/u0/X [22]),
        .I2(\u0/u0/X [21]),
        .I3(\u0/u0/X [20]),
        .I4(\u0/u0/X [24]),
        .I5(\u0/u0/X [19]),
        .O(\u0/out0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__40
       (.I0(\u0/u5/X [17]),
        .I1(\u0/u5/X [16]),
        .I2(\u0/u5/X [15]),
        .I3(\u0/u5/X [14]),
        .I4(\u0/u5/X [18]),
        .I5(\u0/u5/X [13]),
        .O(\u0/out5 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__40_i_1
       (.I0(\u0/R4 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[55] ),
        .I3(\u0/uk/K_r4_reg_n_0_[4] ),
        .O(\u0/u5/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__40_i_2
       (.I0(\u0/R4 [11]),
        .I1(decrypt),
        .I2(\u0/uk/p_49_in ),
        .I3(\u0/uk/p_47_in ),
        .O(\u0/u5/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__40_i_3
       (.I0(\u0/R4 [10]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[39] ),
        .I3(\u0/uk/K_r4_reg_n_0_[20] ),
        .O(\u0/u5/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__40_i_4
       (.I0(\u0/R4 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[6] ),
        .I3(\u0/uk/K_r4_reg_n_0_[12] ),
        .O(\u0/u5/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__40_i_5
       (.I0(\u0/R4 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[11] ),
        .I3(\u0/uk/K_r4_reg_n_0_[17] ),
        .O(\u0/u5/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__40_i_6
       (.I0(\u0/R4 [8]),
        .I1(decrypt),
        .I2(\u0/uk/p_50_in ),
        .I3(\u0/uk/p_49_in ),
        .O(\u0/u5/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__41
       (.I0(\u0/u5/X [35]),
        .I1(\u0/u5/X [34]),
        .I2(\u0/u5/X [33]),
        .I3(\u0/u5/X [32]),
        .I4(\u0/u5/X [36]),
        .I5(\u0/u5/X [31]),
        .O(\u0/out5 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__41_i_1
       (.I0(\u0/R4 [24]),
        .I1(decrypt),
        .I2(\u0/uk/p_44_in ),
        .I3(\u0/uk/K_r4_reg_n_0_[51] ),
        .O(\u0/u5/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__41_i_2
       (.I0(\u0/R4 [23]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[45] ),
        .I3(\u0/uk/K_r4_reg_n_0_[49] ),
        .O(\u0/u5/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__41_i_3
       (.I0(\u0/R4 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[28] ),
        .I3(\u0/uk/K_r4_reg_n_0_[36] ),
        .O(\u0/u5/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__41_i_4
       (.I0(\u0/R4 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[37] ),
        .I3(\u0/uk/K_r4_reg_n_0_[14] ),
        .O(\u0/u5/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__41_i_5
       (.I0(\u0/R4 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[7] ),
        .I3(\u0/uk/K_r4_reg_n_0_[15] ),
        .O(\u0/u5/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__41_i_6
       (.I0(\u0/R4 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[22] ),
        .I3(\u0/uk/K_r4_reg_n_0_[30] ),
        .O(\u0/u5/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__42
       (.I0(\u0/u5/X [11]),
        .I1(\u0/u5/X [10]),
        .I2(\u0/u5/X [9]),
        .I3(\u0/u5/X [8]),
        .I4(\u0/u5/X [12]),
        .I5(\u0/u5/X [7]),
        .O(\u0/out5 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__42_i_1
       (.I0(\u0/R4 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[20] ),
        .I3(\u0/uk/K_r4_reg_n_0_[26] ),
        .O(\u0/u5/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__42_i_2
       (.I0(\u0/R4 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[54] ),
        .I3(\u0/uk/K_r4_reg_n_0_[3] ),
        .O(\u0/u5/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__42_i_3
       (.I0(\u0/R4 [6]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[3] ),
        .I3(\u0/uk/K_r4_reg_n_0_[41] ),
        .O(\u0/u5/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__42_i_4
       (.I0(\u0/R4 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[12] ),
        .I3(\u0/uk/K_r4_reg_n_0_[18] ),
        .O(\u0/u5/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__42_i_5
       (.I0(\u0/R4 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[25] ),
        .I3(\u0/uk/K_r4_reg_n_0_[6] ),
        .O(\u0/u5/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__42_i_6
       (.I0(\u0/R4 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[33] ),
        .I3(\u0/uk/K_r4_reg_n_0_[39] ),
        .O(\u0/u5/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__43
       (.I0(\u0/u5/X [47]),
        .I1(\u0/u5/X [46]),
        .I2(\u0/u5/X [45]),
        .I3(\u0/u5/X [44]),
        .I4(\u0/u5/X [48]),
        .I5(\u0/u5/X [43]),
        .O(\u0/out5 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__43_i_1
       (.I0(\u0/R4 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[15] ),
        .I3(\u0/uk/K_r4_reg_n_0_[23] ),
        .O(\u0/u5/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__43_i_2
       (.I0(\u0/R4 [31]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[9] ),
        .I3(\u0/uk/K_r4_reg_n_0_[45] ),
        .O(\u0/u5/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__43_i_3
       (.I0(\u0/R4 [30]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[21] ),
        .I3(\u0/uk/K_r4_reg_n_0_[29] ),
        .O(\u0/u5/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__43_i_4
       (.I0(\u0/R4 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[51] ),
        .I3(\u0/uk/K_r4_reg_n_0_[28] ),
        .O(\u0/u5/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__43_i_5
       (.I0(\u0/R4 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[36] ),
        .I3(\u0/uk/K_r4_reg_n_0_[44] ),
        .O(\u0/u5/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__43_i_6
       (.I0(\u0/R4 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[52] ),
        .I3(\u0/uk/K_r4_reg_n_0_[1] ),
        .O(\u0/u5/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__44
       (.I0(\u0/u5/X [23]),
        .I1(\u0/u5/X [22]),
        .I2(\u0/u5/X [21]),
        .I3(\u0/u5/X [20]),
        .I4(\u0/u5/X [24]),
        .I5(\u0/u5/X [19]),
        .O(\u0/out5 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__44_i_1
       (.I0(\u0/R4 [16]),
        .I1(decrypt),
        .I2(\u0/uk/p_47_in ),
        .I3(\u0/uk/K_r4_reg_n_0_[27] ),
        .O(\u0/u5/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__44_i_2
       (.I0(\u0/R4 [15]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[13] ),
        .I3(\u0/uk/K_r4_reg_n_0_[19] ),
        .O(\u0/u5/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__44_i_3
       (.I0(\u0/R4 [14]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[5] ),
        .I3(\u0/uk/K_r4_reg_n_0_[11] ),
        .O(\u0/u5/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__44_i_4
       (.I0(\u0/R4 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[4] ),
        .I3(\u0/uk/K_r4_reg_n_0_[10] ),
        .O(\u0/u5/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__44_i_5
       (.I0(\u0/R4 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[26] ),
        .I3(\u0/uk/K_r4_reg_n_0_[32] ),
        .O(\u0/u5/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__44_i_6
       (.I0(\u0/R4 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[10] ),
        .I3(\u0/uk/K_r4_reg_n_0_[48] ),
        .O(\u0/u5/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__45
       (.I0(\u0/u5/X [29]),
        .I1(\u0/u5/X [28]),
        .I2(\u0/u5/X [27]),
        .I3(\u0/u5/X [26]),
        .I4(\u0/u5/X [30]),
        .I5(\u0/u5/X [25]),
        .O(\u0/out5 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__45_i_1
       (.I0(\u0/R4 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_ ),
        .I3(\u0/uk/p_42_in ),
        .O(\u0/u5/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__45_i_2
       (.I0(\u0/R4 [19]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[16] ),
        .I3(\u0/uk/K_r4_reg_n_0_[52] ),
        .O(\u0/u5/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__45_i_3
       (.I0(\u0/R4 [18]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[29] ),
        .I3(\u0/uk/K_r4_reg_n_0_[37] ),
        .O(\u0/u5/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__45_i_4
       (.I0(\u0/R4 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[35] ),
        .I3(\u0/uk/p_44_in ),
        .O(\u0/u5/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__45_i_5
       (.I0(\u0/R4 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[1] ),
        .I3(\u0/uk/K_r4_reg_n_0_[9] ),
        .O(\u0/u5/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__45_i_6
       (.I0(\u0/R4 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[44] ),
        .I3(\u0/uk/K_r4_reg_n_0_[21] ),
        .O(\u0/u5/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__46
       (.I0(\u0/u5/X [5]),
        .I1(\u0/u5/X [4]),
        .I2(\u0/u5/X [3]),
        .I3(\u0/u5/X [2]),
        .I4(\u0/u5/X [6]),
        .I5(\u0/u5/X [1]),
        .O(\u0/out5 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__46_i_1
       (.I0(\u0/R4 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[19] ),
        .I3(\u0/uk/K_r4_reg_n_0_[25] ),
        .O(\u0/u5/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__46_i_2
       (.I0(\u0/R4 [3]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[41] ),
        .I3(\u0/uk/K_r4_reg_n_0_[47] ),
        .O(\u0/u5/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__46_i_3
       (.I0(\u0/R4 [2]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[32] ),
        .I3(\u0/uk/K_r4_reg_n_0_[13] ),
        .O(\u0/u5/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__46_i_4
       (.I0(\u0/R4 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[17] ),
        .I3(\u0/uk/K_r4_reg_n_0_[55] ),
        .O(\u0/u5/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__46_i_5
       (.I0(\u0/R4 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r4_reg_n_0_[47] ),
        .I3(\u0/uk/p_51_in ),
        .O(\u0/u5/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__46_i_6
       (.I0(\u0/R4 [32]),
        .I1(decrypt),
        .I2(\u0/uk/p_51_in ),
        .I3(\u0/uk/p_50_in ),
        .O(\u0/u5/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__47
       (.I0(\u0/u6/X [41]),
        .I1(\u0/u6/X [40]),
        .I2(\u0/u6/X [39]),
        .I3(\u0/u6/X [38]),
        .I4(\u0/u6/X [42]),
        .I5(\u0/u6/X [37]),
        .O(\u0/out6 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__47_i_1
       (.I0(\u0/R5 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [9]),
        .I3(\u0/uk/K_r5 [44]),
        .O(\u0/u6/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__47_i_2
       (.I0(\u0/R5 [27]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [22]),
        .I3(\u0/uk/K_r5 [2]),
        .O(\u0/u6/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__47_i_3
       (.I0(\u0/R5 [26]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [44]),
        .I3(\u0/uk/K_r5 [52]),
        .O(\u0/u6/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__47_i_4
       (.I0(\u0/R5 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [28]),
        .I3(\u0/uk/K_r5 [8]),
        .O(\u0/u6/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__47_i_5
       (.I0(\u0/R5 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [1]),
        .I3(\u0/uk/K_r5 [36]),
        .O(\u0/u6/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__47_i_6
       (.I0(\u0/R5 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [52]),
        .I3(\u0/uk/K_r5 [28]),
        .O(\u0/u6/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__48
       (.I0(\u0/u6/X [17]),
        .I1(\u0/u6/X [16]),
        .I2(\u0/u6/X [15]),
        .I3(\u0/u6/X [14]),
        .I4(\u0/u6/X [18]),
        .I5(\u0/u6/X [13]),
        .O(\u0/out6 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__48_i_1
       (.I0(\u0/R5 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [12]),
        .I3(\u0/uk/K_r5 [47]),
        .O(\u0/u6/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__48_i_2
       (.I0(\u0/R5 [11]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [54]),
        .I3(\u0/uk/K_r5 [32]),
        .O(\u0/u6/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__48_i_3
       (.I0(\u0/R5 [10]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [53]),
        .I3(\u0/uk/K_r5 [6]),
        .O(\u0/u6/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__48_i_4
       (.I0(\u0/R5 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [20]),
        .I3(\u0/uk/K_r5 [55]),
        .O(\u0/u6/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__48_i_5
       (.I0(\u0/R5 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [25]),
        .I3(\u0/uk/K_r5 [3]),
        .O(\u0/u6/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__48_i_6
       (.I0(\u0/R5 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [48]),
        .I3(\u0/uk/K_r5 [26]),
        .O(\u0/u6/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__49
       (.I0(\u0/u6/X [35]),
        .I1(\u0/u6/X [34]),
        .I2(\u0/u6/X [33]),
        .I3(\u0/u6/X [32]),
        .I4(\u0/u6/X [36]),
        .I5(\u0/u6/X [31]),
        .O(\u0/out6 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__49_i_1
       (.I0(\u0/R5 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [2]),
        .I3(\u0/uk/K_r5 [37]),
        .O(\u0/u6/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__49_i_2
       (.I0(\u0/R5 [23]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [0]),
        .I3(\u0/uk/K_r5 [35]),
        .O(\u0/u6/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__49_i_3
       (.I0(\u0/R5 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [42]),
        .I3(\u0/uk/K_r5 [22]),
        .O(\u0/u6/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__49_i_4
       (.I0(\u0/R5 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [51]),
        .I3(\u0/uk/K_r5 [0]),
        .O(\u0/u6/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__49_i_5
       (.I0(\u0/R5 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [21]),
        .I3(\u0/uk/K_r5 [1]),
        .O(\u0/u6/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__49_i_6
       (.I0(\u0/R5 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [36]),
        .I3(\u0/uk/K_r5 [16]),
        .O(\u0/u6/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__4_i_1
       (.I0(\u0/IP [48]),
        .I1(decrypt),
        .I2(\u0/key_r [40]),
        .I3(\u0/key_r [33]),
        .O(\u0/u0/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__4_i_2
       (.I0(\u0/IP [47]),
        .I1(decrypt),
        .I2(\u0/key_r [32]),
        .I3(\u0/key_r [25]),
        .O(\u0/u0/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__4_i_3
       (.I0(\u0/IP [46]),
        .I1(decrypt),
        .I2(\u0/key_r [24]),
        .I3(\u0/key_r [17]),
        .O(\u0/u0/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__4_i_4
       (.I0(\u0/IP [45]),
        .I1(decrypt),
        .I2(\u0/key_r [55]),
        .I3(\u0/key_r [48]),
        .O(\u0/u0/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__4_i_5
       (.I0(\u0/IP [49]),
        .I1(decrypt),
        .I2(\u0/key_r [20]),
        .I3(\u0/key_r [13]),
        .O(\u0/u0/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__4_i_6
       (.I0(\u0/IP [44]),
        .I1(decrypt),
        .I2(\u0/key_r [4]),
        .I3(\u0/key_r [54]),
        .O(\u0/u0/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__5
       (.I0(\u0/u0/X [29]),
        .I1(\u0/u0/X [28]),
        .I2(\u0/u0/X [27]),
        .I3(\u0/u0/X [26]),
        .I4(\u0/u0/X [30]),
        .I5(\u0/u0/X [25]),
        .O(\u0/out0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__50
       (.I0(\u0/u6/X [11]),
        .I1(\u0/u6/X [10]),
        .I2(\u0/u6/X [9]),
        .I3(\u0/u6/X [8]),
        .I4(\u0/u6/X [12]),
        .I5(\u0/u6/X [7]),
        .O(\u0/out6 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__50_i_1
       (.I0(\u0/R5 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [34]),
        .I3(\u0/uk/K_r5 [12]),
        .O(\u0/u6/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__50_i_2
       (.I0(\u0/R5 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [11]),
        .I3(\u0/uk/K_r5 [46]),
        .O(\u0/u6/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__50_i_3
       (.I0(\u0/R5 [6]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [17]),
        .I3(\u0/uk/K_r5 [27]),
        .O(\u0/u6/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__50_i_4
       (.I0(\u0/R5 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [26]),
        .I3(\u0/uk/K_r5 [4]),
        .O(\u0/u6/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__50_i_5
       (.I0(\u0/R5 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [39]),
        .I3(\u0/uk/K_r5 [17]),
        .O(\u0/u6/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__50_i_6
       (.I0(\u0/R5 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [47]),
        .I3(\u0/uk/K_r5 [25]),
        .O(\u0/u6/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__51
       (.I0(\u0/u6/X [47]),
        .I1(\u0/u6/X [46]),
        .I2(\u0/u6/X [45]),
        .I3(\u0/u6/X [44]),
        .I4(\u0/u6/X [48]),
        .I5(\u0/u6/X [43]),
        .O(\u0/out6 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__51_i_1
       (.I0(\u0/R5 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [29]),
        .I3(\u0/uk/K_r5 [9]),
        .O(\u0/u6/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__51_i_2
       (.I0(\u0/R5 [31]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [23]),
        .I3(\u0/uk/K_r5 [31]),
        .O(\u0/u6/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__51_i_3
       (.I0(\u0/R5 [30]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [35]),
        .I3(\u0/uk/K_r5 [15]),
        .O(\u0/u6/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__51_i_4
       (.I0(\u0/R5 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [38]),
        .I3(\u0/uk/K_r5 [14]),
        .O(\u0/u6/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__51_i_5
       (.I0(\u0/R5 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [50]),
        .I3(\u0/uk/K_r5 [30]),
        .O(\u0/u6/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__51_i_6
       (.I0(\u0/R5 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [7]),
        .I3(\u0/uk/K_r5 [42]),
        .O(\u0/u6/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__52
       (.I0(\u0/u6/X [23]),
        .I1(\u0/u6/X [22]),
        .I2(\u0/u6/X [21]),
        .I3(\u0/u6/X [20]),
        .I4(\u0/u6/X [24]),
        .I5(\u0/u6/X [19]),
        .O(\u0/out6 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__52_i_1
       (.I0(\u0/R5 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [3]),
        .I3(\u0/uk/K_r5 [13]),
        .O(\u0/u6/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__52_i_2
       (.I0(\u0/R5 [15]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [27]),
        .I3(\u0/uk/K_r5 [5]),
        .O(\u0/u6/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__52_i_3
       (.I0(\u0/R5 [14]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [19]),
        .I3(\u0/uk/K_r5 [54]),
        .O(\u0/u6/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__52_i_4
       (.I0(\u0/R5 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [18]),
        .I3(\u0/uk/K_r5 [53]),
        .O(\u0/u6/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__52_i_5
       (.I0(\u0/R5 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [40]),
        .I3(\u0/uk/K_r5 [18]),
        .O(\u0/u6/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__52_i_6
       (.I0(\u0/R5 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [24]),
        .I3(\u0/uk/K_r5 [34]),
        .O(\u0/u6/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__53
       (.I0(\u0/u6/X [29]),
        .I1(\u0/u6/X [28]),
        .I2(\u0/u6/X [27]),
        .I3(\u0/u6/X [26]),
        .I4(\u0/u6/X [30]),
        .I5(\u0/u6/X [25]),
        .O(\u0/out6 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__53_i_1
       (.I0(\u0/R5 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [14]),
        .I3(\u0/uk/K_r5 [49]),
        .O(\u0/u6/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__53_i_2
       (.I0(\u0/R5 [19]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [30]),
        .I3(\u0/uk/K_r5 [38]),
        .O(\u0/u6/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__53_i_3
       (.I0(\u0/R5 [18]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [43]),
        .I3(\u0/uk/K_r5 [23]),
        .O(\u0/u6/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__53_i_4
       (.I0(\u0/R5 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [49]),
        .I3(\u0/uk/K_r5 [29]),
        .O(\u0/u6/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__53_i_5
       (.I0(\u0/R5 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [15]),
        .I3(\u0/uk/K_r5 [50]),
        .O(\u0/u6/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__53_i_6
       (.I0(\u0/R5 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [31]),
        .I3(\u0/uk/K_r5 [7]),
        .O(\u0/u6/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__54
       (.I0(\u0/u6/X [5]),
        .I1(\u0/u6/X [4]),
        .I2(\u0/u6/X [3]),
        .I3(\u0/u6/X [2]),
        .I4(\u0/u6/X [6]),
        .I5(\u0/u6/X [1]),
        .O(\u0/out6 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__54_i_1
       (.I0(\u0/R5 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [33]),
        .I3(\u0/uk/K_r5 [11]),
        .O(\u0/u6/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__54_i_2
       (.I0(\u0/R5 [3]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [55]),
        .I3(\u0/uk/K_r5 [33]),
        .O(\u0/u6/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__54_i_3
       (.I0(\u0/R5 [2]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [46]),
        .I3(\u0/uk/K_r5 [24]),
        .O(\u0/u6/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__54_i_4
       (.I0(\u0/R5 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [6]),
        .I3(\u0/uk/K_r5 [41]),
        .O(\u0/u6/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__54_i_5
       (.I0(\u0/R5 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [4]),
        .I3(\u0/uk/K_r5 [39]),
        .O(\u0/u6/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__54_i_6
       (.I0(\u0/R5 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r5 [10]),
        .I3(\u0/uk/K_r5 [20]),
        .O(\u0/u6/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__55
       (.I0(\u0/u7/X [41]),
        .I1(\u0/u7/X [40]),
        .I2(\u0/u7/X [39]),
        .I3(\u0/u7/X [38]),
        .I4(\u0/u7/X [42]),
        .I5(\u0/u7/X [37]),
        .O(\u0/out7 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__55_i_1
       (.I0(\u0/R6 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[23] ),
        .I3(\u0/uk/K_r6_reg_n_0_[30] ),
        .O(\u0/u7/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__55_i_2
       (.I0(\u0/R6 [27]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[36] ),
        .I3(\u0/uk/p_45_in ),
        .O(\u0/u7/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__55_i_3
       (.I0(\u0/R6 [26]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[31] ),
        .I3(\u0/uk/K_r6_reg_n_0_[38] ),
        .O(\u0/u7/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__55_i_4
       (.I0(\u0/R6 [25]),
        .I1(decrypt),
        .I2(\u0/uk/p_41_in ),
        .I3(\u0/uk/p_43_in ),
        .O(\u0/u7/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__55_i_5
       (.I0(\u0/R6 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[15] ),
        .I3(\u0/uk/K_r6_reg_n_0_[22] ),
        .O(\u0/u7/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__55_i_6
       (.I0(\u0/R6 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[7] ),
        .I3(\u0/uk/K_r6_reg_n_0_[14] ),
        .O(\u0/u7/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__56
       (.I0(\u0/u7/X [17]),
        .I1(\u0/u7/X [16]),
        .I2(\u0/u7/X [15]),
        .I3(\u0/u7/X [14]),
        .I4(\u0/u7/X [18]),
        .I5(\u0/u7/X [13]),
        .O(\u0/out7 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__56_i_1
       (.I0(\u0/R6 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[26] ),
        .I3(\u0/uk/K_r6_reg_n_0_[33] ),
        .O(\u0/u7/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__56_i_2
       (.I0(\u0/R6 [11]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[11] ),
        .I3(\u0/uk/K_r6_reg_n_0_[18] ),
        .O(\u0/u7/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__56_i_3
       (.I0(\u0/R6 [10]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[10] ),
        .I3(\u0/uk/K_r6_reg_n_0_[17] ),
        .O(\u0/u7/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__56_i_4
       (.I0(\u0/R6 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[34] ),
        .I3(\u0/uk/K_r6_reg_n_0_[41] ),
        .O(\u0/u7/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__56_i_5
       (.I0(\u0/R6 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[39] ),
        .I3(\u0/uk/K_r6_reg_n_0_[46] ),
        .O(\u0/u7/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__56_i_6
       (.I0(\u0/R6 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[5] ),
        .I3(\u0/uk/K_r6_reg_n_0_[12] ),
        .O(\u0/u7/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__57
       (.I0(\u0/u7/X [35]),
        .I1(\u0/u7/X [34]),
        .I2(\u0/u7/X [33]),
        .I3(\u0/u7/X [32]),
        .I4(\u0/u7/X [36]),
        .I5(\u0/u7/X [31]),
        .O(\u0/out7 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__57_i_1
       (.I0(\u0/R6 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[16] ),
        .I3(\u0/uk/K_r6_reg_n_0_[23] ),
        .O(\u0/u7/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__57_i_2
       (.I0(\u0/R6 [23]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[14] ),
        .I3(\u0/uk/K_r6_reg_n_0_[21] ),
        .O(\u0/u7/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__57_i_3
       (.I0(\u0/R6 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[1] ),
        .I3(\u0/uk/K_r6_reg_n_0_[8] ),
        .O(\u0/u7/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__57_i_4
       (.I0(\u0/R6 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[38] ),
        .I3(\u0/uk/K_r6_reg_n_0_[45] ),
        .O(\u0/u7/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__57_i_5
       (.I0(\u0/R6 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[35] ),
        .I3(\u0/uk/p_41_in ),
        .O(\u0/u7/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__57_i_6
       (.I0(\u0/R6 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[50] ),
        .I3(\u0/uk/K_r6_reg_n_0_[2] ),
        .O(\u0/u7/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__58
       (.I0(\u0/u7/X [11]),
        .I1(\u0/u7/X [10]),
        .I2(\u0/u7/X [9]),
        .I3(\u0/u7/X [8]),
        .I4(\u0/u7/X [12]),
        .I5(\u0/u7/X [7]),
        .O(\u0/out7 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__58_i_1
       (.I0(\u0/R6 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[48] ),
        .I3(\u0/uk/K_r6_reg_n_0_[55] ),
        .O(\u0/u7/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__58_i_2
       (.I0(\u0/R6 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[25] ),
        .I3(\u0/uk/K_r6_reg_n_0_[32] ),
        .O(\u0/u7/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__58_i_3
       (.I0(\u0/R6 [6]),
        .I1(decrypt),
        .I2(\u0/uk/p_53_in ),
        .I3(\u0/uk/p_52_in ),
        .O(\u0/u7/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__58_i_4
       (.I0(\u0/R6 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[40] ),
        .I3(\u0/uk/K_r6_reg_n_0_[47] ),
        .O(\u0/u7/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__58_i_5
       (.I0(\u0/R6 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[53] ),
        .I3(\u0/uk/K_r6_reg_n_0_[3] ),
        .O(\u0/u7/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__58_i_6
       (.I0(\u0/R6 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[4] ),
        .I3(\u0/uk/K_r6_reg_n_0_[11] ),
        .O(\u0/u7/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__59
       (.I0(\u0/u7/X [47]),
        .I1(\u0/u7/X [46]),
        .I2(\u0/u7/X [45]),
        .I3(\u0/u7/X [44]),
        .I4(\u0/u7/X [48]),
        .I5(\u0/u7/X [43]),
        .O(\u0/out7 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__59_i_1
       (.I0(\u0/R6 [32]),
        .I1(decrypt),
        .I2(\u0/uk/p_45_in ),
        .I3(\u0/uk/K_r6_reg_n_0_[50] ),
        .O(\u0/u7/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__59_i_2
       (.I0(\u0/R6 [31]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[37] ),
        .I3(\u0/uk/K_r6_reg_n_0_[44] ),
        .O(\u0/u7/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__59_i_3
       (.I0(\u0/R6 [30]),
        .I1(decrypt),
        .I2(\u0/uk/p_43_in ),
        .I3(\u0/uk/K_r6_reg_n_0_[1] ),
        .O(\u0/u7/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__59_i_4
       (.I0(\u0/R6 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[52] ),
        .I3(\u0/uk/K_r6_reg_n_0_ ),
        .O(\u0/u7/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__59_i_5
       (.I0(\u0/R6 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[9] ),
        .I3(\u0/uk/K_r6_reg_n_0_[16] ),
        .O(\u0/u7/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__59_i_6
       (.I0(\u0/R6 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[21] ),
        .I3(\u0/uk/K_r6_reg_n_0_[28] ),
        .O(\u0/u7/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__5_i_1
       (.I0(\u0/IP [52]),
        .I1(decrypt),
        .I2(\u0/key_r [23]),
        .I3(\u0/key_r [16]),
        .O(\u0/u0/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__5_i_2
       (.I0(\u0/IP [51]),
        .I1(decrypt),
        .I2(\u0/key_r [8]),
        .I3(\u0/key_r [1]),
        .O(\u0/u0/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__5_i_3
       (.I0(\u0/IP [50]),
        .I1(decrypt),
        .I2(\u0/key_r [21]),
        .I3(\u0/key_r [14]),
        .O(\u0/u0/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__5_i_4
       (.I0(\u0/IP [49]),
        .I1(decrypt),
        .I2(\u0/key_r [31]),
        .I3(\u0/key_r [51]),
        .O(\u0/u0/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__5_i_5
       (.I0(\u0/IP [53]),
        .I1(decrypt),
        .I2(\u0/key_r [52]),
        .I3(\u0/key_r [45]),
        .O(\u0/u0/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__5_i_6
       (.I0(\u0/IP [48]),
        .I1(decrypt),
        .I2(\u0/key_r [36]),
        .I3(\u0/key_r [29]),
        .O(\u0/u0/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__6
       (.I0(\u0/u0/X [5]),
        .I1(\u0/u0/X [4]),
        .I2(\u0/u0/X [3]),
        .I3(\u0/u0/X [2]),
        .I4(\u0/u0/X [6]),
        .I5(\u0/u0/X [1]),
        .O(\u0/out0 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__60
       (.I0(\u0/u7/X [23]),
        .I1(\u0/u7/X [22]),
        .I2(\u0/u7/X [21]),
        .I3(\u0/u7/X [20]),
        .I4(\u0/u7/X [24]),
        .I5(\u0/u7/X [19]),
        .O(\u0/out7 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__60_i_1
       (.I0(\u0/R6 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[17] ),
        .I3(\u0/uk/K_r6_reg_n_0_[24] ),
        .O(\u0/u7/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__60_i_2
       (.I0(\u0/R6 [15]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[41] ),
        .I3(\u0/uk/K_r6_reg_n_0_[48] ),
        .O(\u0/u7/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__60_i_3
       (.I0(\u0/R6 [14]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[33] ),
        .I3(\u0/uk/K_r6_reg_n_0_[40] ),
        .O(\u0/u7/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__60_i_4
       (.I0(\u0/R6 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[32] ),
        .I3(\u0/uk/K_r6_reg_n_0_[39] ),
        .O(\u0/u7/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__60_i_5
       (.I0(\u0/R6 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[54] ),
        .I3(\u0/uk/K_r6_reg_n_0_[4] ),
        .O(\u0/u7/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__60_i_6
       (.I0(\u0/R6 [12]),
        .I1(decrypt),
        .I2(\u0/uk/p_52_in ),
        .I3(\u0/uk/K_r6_reg_n_0_[20] ),
        .O(\u0/u7/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__61
       (.I0(\u0/u7/X [29]),
        .I1(\u0/u7/X [28]),
        .I2(\u0/u7/X [27]),
        .I3(\u0/u7/X [26]),
        .I4(\u0/u7/X [30]),
        .I5(\u0/u7/X [25]),
        .O(\u0/out7 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__61_i_1
       (.I0(\u0/R6 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[28] ),
        .I3(\u0/uk/K_r6_reg_n_0_[35] ),
        .O(\u0/u7/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__61_i_2
       (.I0(\u0/R6 [19]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[44] ),
        .I3(\u0/uk/K_r6_reg_n_0_[51] ),
        .O(\u0/u7/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__61_i_3
       (.I0(\u0/R6 [18]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[2] ),
        .I3(\u0/uk/K_r6_reg_n_0_[9] ),
        .O(\u0/u7/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__61_i_4
       (.I0(\u0/R6 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[8] ),
        .I3(\u0/uk/K_r6_reg_n_0_[15] ),
        .O(\u0/u7/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__61_i_5
       (.I0(\u0/R6 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[29] ),
        .I3(\u0/uk/K_r6_reg_n_0_[36] ),
        .O(\u0/u7/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__61_i_6
       (.I0(\u0/R6 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[45] ),
        .I3(\u0/uk/K_r6_reg_n_0_[52] ),
        .O(\u0/u7/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__62
       (.I0(\u0/u7/X [5]),
        .I1(\u0/u7/X [4]),
        .I2(\u0/u7/X [3]),
        .I3(\u0/u7/X [2]),
        .I4(\u0/u7/X [6]),
        .I5(\u0/u7/X [1]),
        .O(\u0/out7 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__62_i_1
       (.I0(\u0/R6 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[47] ),
        .I3(\u0/uk/K_r6_reg_n_0_[54] ),
        .O(\u0/u7/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__62_i_2
       (.I0(\u0/R6 [3]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[12] ),
        .I3(\u0/uk/K_r6_reg_n_0_[19] ),
        .O(\u0/u7/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__62_i_3
       (.I0(\u0/R6 [2]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[3] ),
        .I3(\u0/uk/K_r6_reg_n_0_[10] ),
        .O(\u0/u7/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__62_i_4
       (.I0(\u0/R6 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[20] ),
        .I3(\u0/uk/K_r6_reg_n_0_[27] ),
        .O(\u0/u7/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__62_i_5
       (.I0(\u0/R6 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[18] ),
        .I3(\u0/uk/K_r6_reg_n_0_[25] ),
        .O(\u0/u7/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__62_i_6
       (.I0(\u0/R6 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r6_reg_n_0_[24] ),
        .I3(\u0/uk/p_53_in ),
        .O(\u0/u7/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__63
       (.I0(\u0/u8/X [41]),
        .I1(\u0/u8/X [40]),
        .I2(\u0/u8/X [39]),
        .I3(\u0/u8/X [38]),
        .I4(\u0/u8/X [42]),
        .I5(\u0/u8/X [37]),
        .O(\u0/out8 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__63_i_1
       (.I0(\u0/R7 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[30] ),
        .I3(\u0/uk/K_r7_reg_n_0_[23] ),
        .O(\u0/u8/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__63_i_2
       (.I0(\u0/R7 [27]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[43] ),
        .I3(\u0/uk/K_r7_reg_n_0_[36] ),
        .O(\u0/u8/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__63_i_3
       (.I0(\u0/R7 [26]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[38] ),
        .I3(\u0/uk/K_r7_reg_n_0_[31] ),
        .O(\u0/u8/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__63_i_4
       (.I0(\u0/R7 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[49] ),
        .I3(\u0/uk/K_r7_reg_n_0_[42] ),
        .O(\u0/u8/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__63_i_5
       (.I0(\u0/R7 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[22] ),
        .I3(\u0/uk/K_r7_reg_n_0_[15] ),
        .O(\u0/u8/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__63_i_6
       (.I0(\u0/R7 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[14] ),
        .I3(\u0/uk/K_r7_reg_n_0_[7] ),
        .O(\u0/u8/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__64
       (.I0(\u0/u8/X [17]),
        .I1(\u0/u8/X [16]),
        .I2(\u0/u8/X [15]),
        .I3(\u0/u8/X [14]),
        .I4(\u0/u8/X [18]),
        .I5(\u0/u8/X [13]),
        .O(\u0/out8 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__64_i_1
       (.I0(\u0/R7 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[33] ),
        .I3(\u0/uk/K_r7_reg_n_0_[26] ),
        .O(\u0/u8/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__64_i_2
       (.I0(\u0/R7 [11]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[18] ),
        .I3(\u0/uk/K_r7_reg_n_0_[11] ),
        .O(\u0/u8/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__64_i_3
       (.I0(\u0/R7 [10]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[17] ),
        .I3(\u0/uk/K_r7_reg_n_0_[10] ),
        .O(\u0/u8/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__64_i_4
       (.I0(\u0/R7 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[41] ),
        .I3(\u0/uk/K_r7_reg_n_0_[34] ),
        .O(\u0/u8/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__64_i_5
       (.I0(\u0/R7 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[46] ),
        .I3(\u0/uk/K_r7_reg_n_0_[39] ),
        .O(\u0/u8/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__64_i_6
       (.I0(\u0/R7 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[12] ),
        .I3(\u0/uk/K_r7_reg_n_0_[5] ),
        .O(\u0/u8/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__65
       (.I0(\u0/u8/X [35]),
        .I1(\u0/u8/X [34]),
        .I2(\u0/u8/X [33]),
        .I3(\u0/u8/X [32]),
        .I4(\u0/u8/X [36]),
        .I5(\u0/u8/X [31]),
        .O(\u0/out8 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__65_i_1
       (.I0(\u0/R7 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[23] ),
        .I3(\u0/uk/K_r7_reg_n_0_[16] ),
        .O(\u0/u8/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__65_i_2
       (.I0(\u0/R7 [23]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[21] ),
        .I3(\u0/uk/K_r7_reg_n_0_[14] ),
        .O(\u0/u8/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__65_i_3
       (.I0(\u0/R7 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[8] ),
        .I3(\u0/uk/K_r7_reg_n_0_[1] ),
        .O(\u0/u8/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__65_i_4
       (.I0(\u0/R7 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[45] ),
        .I3(\u0/uk/K_r7_reg_n_0_[38] ),
        .O(\u0/u8/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__65_i_5
       (.I0(\u0/R7 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[42] ),
        .I3(\u0/uk/K_r7_reg_n_0_[35] ),
        .O(\u0/u8/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__65_i_6
       (.I0(\u0/R7 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[2] ),
        .I3(\u0/uk/K_r7_reg_n_0_[50] ),
        .O(\u0/u8/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__66
       (.I0(\u0/u8/X [11]),
        .I1(\u0/u8/X [10]),
        .I2(\u0/u8/X [9]),
        .I3(\u0/u8/X [8]),
        .I4(\u0/u8/X [12]),
        .I5(\u0/u8/X [7]),
        .O(\u0/out8 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__66_i_1
       (.I0(\u0/R7 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[55] ),
        .I3(\u0/uk/K_r7_reg_n_0_[48] ),
        .O(\u0/u8/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__66_i_2
       (.I0(\u0/R7 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[32] ),
        .I3(\u0/uk/K_r7_reg_n_0_[25] ),
        .O(\u0/u8/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__66_i_3
       (.I0(\u0/R7 [6]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[13] ),
        .I3(\u0/uk/K_r7_reg_n_0_[6] ),
        .O(\u0/u8/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__66_i_4
       (.I0(\u0/R7 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[47] ),
        .I3(\u0/uk/K_r7_reg_n_0_[40] ),
        .O(\u0/u8/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__66_i_5
       (.I0(\u0/R7 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[3] ),
        .I3(\u0/uk/K_r7_reg_n_0_[53] ),
        .O(\u0/u8/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__66_i_6
       (.I0(\u0/R7 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[11] ),
        .I3(\u0/uk/K_r7_reg_n_0_[4] ),
        .O(\u0/u8/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__67
       (.I0(\u0/u8/X [47]),
        .I1(\u0/u8/X [46]),
        .I2(\u0/u8/X [45]),
        .I3(\u0/u8/X [44]),
        .I4(\u0/u8/X [48]),
        .I5(\u0/u8/X [43]),
        .O(\u0/out8 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__67_i_1
       (.I0(\u0/R7 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[50] ),
        .I3(\u0/uk/K_r7_reg_n_0_[43] ),
        .O(\u0/u8/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__67_i_2
       (.I0(\u0/R7 [31]),
        .I1(decrypt),
        .I2(\u0/uk/p_48_in ),
        .I3(\u0/uk/K_r7_reg_n_0_[37] ),
        .O(\u0/u8/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__67_i_3
       (.I0(\u0/R7 [30]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[1] ),
        .I3(\u0/uk/K_r7_reg_n_0_[49] ),
        .O(\u0/u8/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__67_i_4
       (.I0(\u0/R7 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_ ),
        .I3(\u0/uk/K_r7_reg_n_0_[52] ),
        .O(\u0/u8/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__67_i_5
       (.I0(\u0/R7 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[16] ),
        .I3(\u0/uk/K_r7_reg_n_0_[9] ),
        .O(\u0/u8/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__67_i_6
       (.I0(\u0/R7 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[28] ),
        .I3(\u0/uk/K_r7_reg_n_0_[21] ),
        .O(\u0/u8/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__68
       (.I0(\u0/u8/X [23]),
        .I1(\u0/u8/X [22]),
        .I2(\u0/u8/X [21]),
        .I3(\u0/u8/X [20]),
        .I4(\u0/u8/X [24]),
        .I5(\u0/u8/X [19]),
        .O(\u0/out8 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__68_i_1
       (.I0(\u0/R7 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[24] ),
        .I3(\u0/uk/K_r7_reg_n_0_[17] ),
        .O(\u0/u8/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__68_i_2
       (.I0(\u0/R7 [15]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[48] ),
        .I3(\u0/uk/K_r7_reg_n_0_[41] ),
        .O(\u0/u8/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__68_i_3
       (.I0(\u0/R7 [14]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[40] ),
        .I3(\u0/uk/K_r7_reg_n_0_[33] ),
        .O(\u0/u8/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__68_i_4
       (.I0(\u0/R7 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[39] ),
        .I3(\u0/uk/K_r7_reg_n_0_[32] ),
        .O(\u0/u8/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__68_i_5
       (.I0(\u0/R7 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[4] ),
        .I3(\u0/uk/K_r7_reg_n_0_[54] ),
        .O(\u0/u8/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__68_i_6
       (.I0(\u0/R7 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[20] ),
        .I3(\u0/uk/K_r7_reg_n_0_[13] ),
        .O(\u0/u8/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__69
       (.I0(\u0/u8/X [29]),
        .I1(\u0/u8/X [28]),
        .I2(\u0/u8/X [27]),
        .I3(\u0/u8/X [26]),
        .I4(\u0/u8/X [30]),
        .I5(\u0/u8/X [25]),
        .O(\u0/out8 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__69_i_1
       (.I0(\u0/R7 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[35] ),
        .I3(\u0/uk/K_r7_reg_n_0_[28] ),
        .O(\u0/u8/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__69_i_2
       (.I0(\u0/R7 [19]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[51] ),
        .I3(\u0/uk/p_48_in ),
        .O(\u0/u8/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__69_i_3
       (.I0(\u0/R7 [18]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[9] ),
        .I3(\u0/uk/K_r7_reg_n_0_[2] ),
        .O(\u0/u8/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__69_i_4
       (.I0(\u0/R7 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[15] ),
        .I3(\u0/uk/K_r7_reg_n_0_[8] ),
        .O(\u0/u8/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__69_i_5
       (.I0(\u0/R7 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[36] ),
        .I3(\u0/uk/K_r7_reg_n_0_[29] ),
        .O(\u0/u8/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__69_i_6
       (.I0(\u0/R7 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[52] ),
        .I3(\u0/uk/K_r7_reg_n_0_[45] ),
        .O(\u0/u8/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__6_i_1
       (.I0(\u0/IP [36]),
        .I1(decrypt),
        .I2(\u0/key_r [13]),
        .I3(\u0/key_r [6]),
        .O(\u0/u0/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__6_i_2
       (.I0(\u0/IP [35]),
        .I1(decrypt),
        .I2(\u0/key_r [3]),
        .I3(\u0/key_r [53]),
        .O(\u0/u0/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__6_i_3
       (.I0(\u0/IP [34]),
        .I1(decrypt),
        .I2(\u0/key_r [26]),
        .I3(\u0/key_r [19]),
        .O(\u0/u0/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__6_i_4
       (.I0(\u0/IP [33]),
        .I1(decrypt),
        .I2(\u0/key_r [11]),
        .I3(\u0/key_r [4]),
        .O(\u0/u0/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__6_i_5
       (.I0(\u0/IP [37]),
        .I1(decrypt),
        .I2(\u0/key_r [41]),
        .I3(\u0/key_r [34]),
        .O(\u0/u0/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__6_i_6
       (.I0(\u0/IP [64]),
        .I1(decrypt),
        .I2(\u0/key_r [47]),
        .I3(\u0/key_r [40]),
        .O(\u0/u0/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__7
       (.I0(\u0/u1/X [41]),
        .I1(\u0/u1/X [40]),
        .I2(\u0/u1/X [39]),
        .I3(\u0/u1/X [38]),
        .I4(\u0/u1/X [42]),
        .I5(\u0/u1/X [37]),
        .O(\u0/out1 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__70
       (.I0(\u0/u8/X [5]),
        .I1(\u0/u8/X [4]),
        .I2(\u0/u8/X [3]),
        .I3(\u0/u8/X [2]),
        .I4(\u0/u8/X [6]),
        .I5(\u0/u8/X [1]),
        .O(\u0/out8 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__70_i_1
       (.I0(\u0/R7 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[54] ),
        .I3(\u0/uk/K_r7_reg_n_0_[47] ),
        .O(\u0/u8/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__70_i_2
       (.I0(\u0/R7 [3]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[19] ),
        .I3(\u0/uk/K_r7_reg_n_0_[12] ),
        .O(\u0/u8/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__70_i_3
       (.I0(\u0/R7 [2]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[10] ),
        .I3(\u0/uk/K_r7_reg_n_0_[3] ),
        .O(\u0/u8/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__70_i_4
       (.I0(\u0/R7 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[27] ),
        .I3(\u0/uk/K_r7_reg_n_0_[20] ),
        .O(\u0/u8/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__70_i_5
       (.I0(\u0/R7 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[25] ),
        .I3(\u0/uk/K_r7_reg_n_0_[18] ),
        .O(\u0/u8/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__70_i_6
       (.I0(\u0/R7 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r7_reg_n_0_[6] ),
        .I3(\u0/uk/K_r7_reg_n_0_[24] ),
        .O(\u0/u8/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__71
       (.I0(\u0/u9/X [41]),
        .I1(\u0/u9/X [40]),
        .I2(\u0/u9/X [39]),
        .I3(\u0/u9/X [38]),
        .I4(\u0/u9/X [42]),
        .I5(\u0/u9/X [37]),
        .O(\u0/out9 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__71_i_1
       (.I0(\u0/R8 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [44]),
        .I3(\u0/uk/K_r8 [9]),
        .O(\u0/u9/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__71_i_2
       (.I0(\u0/R8 [27]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [2]),
        .I3(\u0/uk/K_r8 [22]),
        .O(\u0/u9/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__71_i_3
       (.I0(\u0/R8 [26]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [52]),
        .I3(\u0/uk/K_r8 [44]),
        .O(\u0/u9/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__71_i_4
       (.I0(\u0/R8 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [8]),
        .I3(\u0/uk/K_r8 [28]),
        .O(\u0/u9/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__71_i_5
       (.I0(\u0/R8 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [36]),
        .I3(\u0/uk/K_r8 [1]),
        .O(\u0/u9/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__71_i_6
       (.I0(\u0/R8 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [28]),
        .I3(\u0/uk/K_r8 [52]),
        .O(\u0/u9/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__72
       (.I0(\u0/u9/X [17]),
        .I1(\u0/u9/X [16]),
        .I2(\u0/u9/X [15]),
        .I3(\u0/u9/X [14]),
        .I4(\u0/u9/X [18]),
        .I5(\u0/u9/X [13]),
        .O(\u0/out9 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__72_i_1
       (.I0(\u0/R8 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [47]),
        .I3(\u0/uk/K_r8 [12]),
        .O(\u0/u9/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__72_i_2
       (.I0(\u0/R8 [11]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [32]),
        .I3(\u0/uk/K_r8 [54]),
        .O(\u0/u9/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__72_i_3
       (.I0(\u0/R8 [10]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [6]),
        .I3(\u0/uk/K_r8 [53]),
        .O(\u0/u9/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__72_i_4
       (.I0(\u0/R8 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [55]),
        .I3(\u0/uk/K_r8 [20]),
        .O(\u0/u9/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__72_i_5
       (.I0(\u0/R8 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [3]),
        .I3(\u0/uk/K_r8 [25]),
        .O(\u0/u9/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__72_i_6
       (.I0(\u0/R8 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [26]),
        .I3(\u0/uk/K_r8 [48]),
        .O(\u0/u9/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__73
       (.I0(\u0/u9/X [35]),
        .I1(\u0/u9/X [34]),
        .I2(\u0/u9/X [33]),
        .I3(\u0/u9/X [32]),
        .I4(\u0/u9/X [36]),
        .I5(\u0/u9/X [31]),
        .O(\u0/out9 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__73_i_1
       (.I0(\u0/R8 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [37]),
        .I3(\u0/uk/K_r8 [2]),
        .O(\u0/u9/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__73_i_2
       (.I0(\u0/R8 [23]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [35]),
        .I3(\u0/uk/K_r8 [0]),
        .O(\u0/u9/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__73_i_3
       (.I0(\u0/R8 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [22]),
        .I3(\u0/uk/K_r8 [42]),
        .O(\u0/u9/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__73_i_4
       (.I0(\u0/R8 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [0]),
        .I3(\u0/uk/K_r8 [51]),
        .O(\u0/u9/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__73_i_5
       (.I0(\u0/R8 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [1]),
        .I3(\u0/uk/K_r8 [21]),
        .O(\u0/u9/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__73_i_6
       (.I0(\u0/R8 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [16]),
        .I3(\u0/uk/K_r8 [36]),
        .O(\u0/u9/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__74
       (.I0(\u0/u9/X [11]),
        .I1(\u0/u9/X [10]),
        .I2(\u0/u9/X [9]),
        .I3(\u0/u9/X [8]),
        .I4(\u0/u9/X [12]),
        .I5(\u0/u9/X [7]),
        .O(\u0/out9 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__74_i_1
       (.I0(\u0/R8 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [12]),
        .I3(\u0/uk/K_r8 [34]),
        .O(\u0/u9/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__74_i_2
       (.I0(\u0/R8 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [46]),
        .I3(\u0/uk/K_r8 [11]),
        .O(\u0/u9/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__74_i_3
       (.I0(\u0/R8 [6]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [27]),
        .I3(\u0/uk/K_r8 [17]),
        .O(\u0/u9/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__74_i_4
       (.I0(\u0/R8 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [4]),
        .I3(\u0/uk/K_r8 [26]),
        .O(\u0/u9/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__74_i_5
       (.I0(\u0/R8 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [17]),
        .I3(\u0/uk/K_r8 [39]),
        .O(\u0/u9/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__74_i_6
       (.I0(\u0/R8 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [25]),
        .I3(\u0/uk/K_r8 [47]),
        .O(\u0/u9/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__75
       (.I0(\u0/u9/X [47]),
        .I1(\u0/u9/X [46]),
        .I2(\u0/u9/X [45]),
        .I3(\u0/u9/X [44]),
        .I4(\u0/u9/X [48]),
        .I5(\u0/u9/X [43]),
        .O(\u0/out9 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__75_i_1
       (.I0(\u0/R8 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [9]),
        .I3(\u0/uk/K_r8 [29]),
        .O(\u0/u9/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__75_i_2
       (.I0(\u0/R8 [31]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [31]),
        .I3(\u0/uk/K_r8 [23]),
        .O(\u0/u9/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__75_i_3
       (.I0(\u0/R8 [30]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [15]),
        .I3(\u0/uk/K_r8 [35]),
        .O(\u0/u9/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__75_i_4
       (.I0(\u0/R8 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [14]),
        .I3(\u0/uk/K_r8 [38]),
        .O(\u0/u9/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__75_i_5
       (.I0(\u0/R8 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [30]),
        .I3(\u0/uk/K_r8 [50]),
        .O(\u0/u9/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__75_i_6
       (.I0(\u0/R8 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [42]),
        .I3(\u0/uk/K_r8 [7]),
        .O(\u0/u9/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__76
       (.I0(\u0/u9/X [23]),
        .I1(\u0/u9/X [22]),
        .I2(\u0/u9/X [21]),
        .I3(\u0/u9/X [20]),
        .I4(\u0/u9/X [24]),
        .I5(\u0/u9/X [19]),
        .O(\u0/out9 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__76_i_1
       (.I0(\u0/R8 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [13]),
        .I3(\u0/uk/K_r8 [3]),
        .O(\u0/u9/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__76_i_2
       (.I0(\u0/R8 [15]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [5]),
        .I3(\u0/uk/K_r8 [27]),
        .O(\u0/u9/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__76_i_3
       (.I0(\u0/R8 [14]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [54]),
        .I3(\u0/uk/K_r8 [19]),
        .O(\u0/u9/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__76_i_4
       (.I0(\u0/R8 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [53]),
        .I3(\u0/uk/K_r8 [18]),
        .O(\u0/u9/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__76_i_5
       (.I0(\u0/R8 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [18]),
        .I3(\u0/uk/K_r8 [40]),
        .O(\u0/u9/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__76_i_6
       (.I0(\u0/R8 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [34]),
        .I3(\u0/uk/K_r8 [24]),
        .O(\u0/u9/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__77
       (.I0(\u0/u9/X [29]),
        .I1(\u0/u9/X [28]),
        .I2(\u0/u9/X [27]),
        .I3(\u0/u9/X [26]),
        .I4(\u0/u9/X [30]),
        .I5(\u0/u9/X [25]),
        .O(\u0/out9 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__77_i_1
       (.I0(\u0/R8 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [49]),
        .I3(\u0/uk/K_r8 [14]),
        .O(\u0/u9/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__77_i_2
       (.I0(\u0/R8 [19]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [38]),
        .I3(\u0/uk/K_r8 [30]),
        .O(\u0/u9/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__77_i_3
       (.I0(\u0/R8 [18]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [23]),
        .I3(\u0/uk/K_r8 [43]),
        .O(\u0/u9/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__77_i_4
       (.I0(\u0/R8 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [29]),
        .I3(\u0/uk/K_r8 [49]),
        .O(\u0/u9/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__77_i_5
       (.I0(\u0/R8 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [50]),
        .I3(\u0/uk/K_r8 [15]),
        .O(\u0/u9/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__77_i_6
       (.I0(\u0/R8 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [7]),
        .I3(\u0/uk/K_r8 [31]),
        .O(\u0/u9/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__78
       (.I0(\u0/u9/X [5]),
        .I1(\u0/u9/X [4]),
        .I2(\u0/u9/X [3]),
        .I3(\u0/u9/X [2]),
        .I4(\u0/u9/X [6]),
        .I5(\u0/u9/X [1]),
        .O(\u0/out9 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__78_i_1
       (.I0(\u0/R8 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [11]),
        .I3(\u0/uk/K_r8 [33]),
        .O(\u0/u9/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__78_i_2
       (.I0(\u0/R8 [3]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [33]),
        .I3(\u0/uk/K_r8 [55]),
        .O(\u0/u9/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__78_i_3
       (.I0(\u0/R8 [2]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [24]),
        .I3(\u0/uk/K_r8 [46]),
        .O(\u0/u9/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__78_i_4
       (.I0(\u0/R8 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [41]),
        .I3(\u0/uk/K_r8 [6]),
        .O(\u0/u9/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__78_i_5
       (.I0(\u0/R8 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [39]),
        .I3(\u0/uk/K_r8 [4]),
        .O(\u0/u9/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__78_i_6
       (.I0(\u0/R8 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r8 [20]),
        .I3(\u0/uk/K_r8 [10]),
        .O(\u0/u9/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__79
       (.I0(\u0/u10/X [41]),
        .I1(\u0/u10/X [40]),
        .I2(\u0/u10/X [39]),
        .I3(\u0/u10/X [38]),
        .I4(\u0/u10/X [42]),
        .I5(\u0/u10/X [37]),
        .O(\u0/out10 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__79_i_1
       (.I0(\u0/R9 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [31]),
        .I3(\u0/uk/K_r9 [50]),
        .O(\u0/u10/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__79_i_2
       (.I0(\u0/R9 [27]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [16]),
        .I3(\u0/uk/K_r9 [8]),
        .O(\u0/u10/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__79_i_3
       (.I0(\u0/R9 [26]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [7]),
        .I3(\u0/uk/K_r9 [30]),
        .O(\u0/u10/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__79_i_4
       (.I0(\u0/R9 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [22]),
        .I3(\u0/uk/K_r9 [14]),
        .O(\u0/u10/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__79_i_5
       (.I0(\u0/R9 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [50]),
        .I3(\u0/uk/K_r9 [42]),
        .O(\u0/u10/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__79_i_6
       (.I0(\u0/R9 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [42]),
        .I3(\u0/uk/K_r9 [38]),
        .O(\u0/u10/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__7_i_1
       (.I0(\u0/R0 [28]),
        .I1(decrypt),
        .I2(\u0/uk/p_34_in ),
        .I3(\u0/uk/p_20_in ),
        .O(\u0/u1/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__7_i_2
       (.I0(\u0/R0 [27]),
        .I1(decrypt),
        .I2(\u0/uk/p_21_in ),
        .I3(\u0/uk/p_33_in ),
        .O(\u0/u1/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__7_i_3
       (.I0(\u0/R0 [26]),
        .I1(decrypt),
        .I2(\u0/uk/p_31_in ),
        .I3(\u0/uk/p_32_in ),
        .O(\u0/u1/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__7_i_4
       (.I0(\u0/R0 [25]),
        .I1(decrypt),
        .I2(\u0/uk/p_19_in ),
        .I3(\u0/uk/p_30_in ),
        .O(\u0/u1/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__7_i_5
       (.I0(\u0/R0 [29]),
        .I1(decrypt),
        .I2(\u0/uk/p_33_in ),
        .I3(\u0/uk/p_35_in ),
        .O(\u0/u1/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__7_i_6
       (.I0(\u0/R0 [24]),
        .I1(decrypt),
        .I2(\u0/uk/p_23_in ),
        .I3(\u0/uk/p_17_in ),
        .O(\u0/u1/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__8
       (.I0(\u0/u1/X [17]),
        .I1(\u0/u1/X [16]),
        .I2(\u0/u1/X [15]),
        .I3(\u0/u1/X [14]),
        .I4(\u0/u1/X [18]),
        .I5(\u0/u1/X [13]),
        .O(\u0/out1 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__80
       (.I0(\u0/u10/X [17]),
        .I1(\u0/u10/X [16]),
        .I2(\u0/u10/X [15]),
        .I3(\u0/u10/X [14]),
        .I4(\u0/u10/X [18]),
        .I5(\u0/u10/X [13]),
        .O(\u0/out10 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__80_i_1
       (.I0(\u0/R9 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [4]),
        .I3(\u0/uk/K_r9 [55]),
        .O(\u0/u10/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__80_i_2
       (.I0(\u0/R9 [11]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [46]),
        .I3(\u0/uk/K_r9 [40]),
        .O(\u0/u10/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__80_i_3
       (.I0(\u0/R9 [10]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [20]),
        .I3(\u0/uk/K_r9 [39]),
        .O(\u0/u10/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__80_i_4
       (.I0(\u0/R9 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [12]),
        .I3(\u0/uk/K_r9 [6]),
        .O(\u0/u10/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__80_i_5
       (.I0(\u0/R9 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [17]),
        .I3(\u0/uk/K_r9 [11]),
        .O(\u0/u10/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__80_i_6
       (.I0(\u0/R9 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [40]),
        .I3(\u0/uk/K_r9 [34]),
        .O(\u0/u10/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__81
       (.I0(\u0/u10/X [35]),
        .I1(\u0/u10/X [34]),
        .I2(\u0/u10/X [33]),
        .I3(\u0/u10/X [32]),
        .I4(\u0/u10/X [36]),
        .I5(\u0/u10/X [31]),
        .O(\u0/out10 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__81_i_1
       (.I0(\u0/R9 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [51]),
        .I3(\u0/uk/K_r9 [43]),
        .O(\u0/u10/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__81_i_2
       (.I0(\u0/R9 [23]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [49]),
        .I3(\u0/uk/K_r9 [45]),
        .O(\u0/u10/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__81_i_3
       (.I0(\u0/R9 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [36]),
        .I3(\u0/uk/K_r9 [28]),
        .O(\u0/u10/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__81_i_4
       (.I0(\u0/R9 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [14]),
        .I3(\u0/uk/K_r9 [37]),
        .O(\u0/u10/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__81_i_5
       (.I0(\u0/R9 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [15]),
        .I3(\u0/uk/K_r9 [7]),
        .O(\u0/u10/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__81_i_6
       (.I0(\u0/R9 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [30]),
        .I3(\u0/uk/K_r9 [22]),
        .O(\u0/u10/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__82
       (.I0(\u0/u10/X [11]),
        .I1(\u0/u10/X [10]),
        .I2(\u0/u10/X [9]),
        .I3(\u0/u10/X [8]),
        .I4(\u0/u10/X [12]),
        .I5(\u0/u10/X [7]),
        .O(\u0/out10 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__82_i_1
       (.I0(\u0/R9 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [26]),
        .I3(\u0/uk/K_r9 [20]),
        .O(\u0/u10/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__82_i_2
       (.I0(\u0/R9 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [3]),
        .I3(\u0/uk/K_r9 [54]),
        .O(\u0/u10/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__82_i_3
       (.I0(\u0/R9 [6]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [41]),
        .I3(\u0/uk/K_r9 [3]),
        .O(\u0/u10/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__82_i_4
       (.I0(\u0/R9 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [18]),
        .I3(\u0/uk/K_r9 [12]),
        .O(\u0/u10/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__82_i_5
       (.I0(\u0/R9 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [6]),
        .I3(\u0/uk/K_r9 [25]),
        .O(\u0/u10/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__82_i_6
       (.I0(\u0/R9 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [39]),
        .I3(\u0/uk/K_r9 [33]),
        .O(\u0/u10/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__83
       (.I0(\u0/u10/X [47]),
        .I1(\u0/u10/X [46]),
        .I2(\u0/u10/X [45]),
        .I3(\u0/u10/X [44]),
        .I4(\u0/u10/X [48]),
        .I5(\u0/u10/X [43]),
        .O(\u0/out10 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__83_i_1
       (.I0(\u0/R9 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [23]),
        .I3(\u0/uk/K_r9 [15]),
        .O(\u0/u10/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__83_i_2
       (.I0(\u0/R9 [31]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [45]),
        .I3(\u0/uk/K_r9 [9]),
        .O(\u0/u10/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__83_i_3
       (.I0(\u0/R9 [30]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [29]),
        .I3(\u0/uk/K_r9 [21]),
        .O(\u0/u10/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__83_i_4
       (.I0(\u0/R9 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [28]),
        .I3(\u0/uk/K_r9 [51]),
        .O(\u0/u10/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__83_i_5
       (.I0(\u0/R9 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [44]),
        .I3(\u0/uk/K_r9 [36]),
        .O(\u0/u10/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__83_i_6
       (.I0(\u0/R9 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [1]),
        .I3(\u0/uk/K_r9 [52]),
        .O(\u0/u10/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__84
       (.I0(\u0/u10/X [23]),
        .I1(\u0/u10/X [22]),
        .I2(\u0/u10/X [21]),
        .I3(\u0/u10/X [20]),
        .I4(\u0/u10/X [24]),
        .I5(\u0/u10/X [19]),
        .O(\u0/out10 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__84_i_1
       (.I0(\u0/R9 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [27]),
        .I3(\u0/uk/K_r9 [46]),
        .O(\u0/u10/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__84_i_2
       (.I0(\u0/R9 [15]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [19]),
        .I3(\u0/uk/K_r9 [13]),
        .O(\u0/u10/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__84_i_3
       (.I0(\u0/R9 [14]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [11]),
        .I3(\u0/uk/K_r9 [5]),
        .O(\u0/u10/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__84_i_4
       (.I0(\u0/R9 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [10]),
        .I3(\u0/uk/K_r9 [4]),
        .O(\u0/u10/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__84_i_5
       (.I0(\u0/R9 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [32]),
        .I3(\u0/uk/K_r9 [26]),
        .O(\u0/u10/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__84_i_6
       (.I0(\u0/R9 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [48]),
        .I3(\u0/uk/K_r9 [10]),
        .O(\u0/u10/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__85
       (.I0(\u0/u10/X [29]),
        .I1(\u0/u10/X [28]),
        .I2(\u0/u10/X [27]),
        .I3(\u0/u10/X [26]),
        .I4(\u0/u10/X [30]),
        .I5(\u0/u10/X [25]),
        .O(\u0/out10 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__85_i_1
       (.I0(\u0/R9 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [8]),
        .I3(\u0/uk/K_r9 [0]),
        .O(\u0/u10/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__85_i_2
       (.I0(\u0/R9 [19]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [52]),
        .I3(\u0/uk/K_r9 [16]),
        .O(\u0/u10/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__85_i_3
       (.I0(\u0/R9 [18]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [37]),
        .I3(\u0/uk/K_r9 [29]),
        .O(\u0/u10/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__85_i_4
       (.I0(\u0/R9 [17]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [43]),
        .I3(\u0/uk/K_r9 [35]),
        .O(\u0/u10/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__85_i_5
       (.I0(\u0/R9 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [9]),
        .I3(\u0/uk/K_r9 [1]),
        .O(\u0/u10/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__85_i_6
       (.I0(\u0/R9 [16]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [21]),
        .I3(\u0/uk/K_r9 [44]),
        .O(\u0/u10/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__86
       (.I0(\u0/u10/X [5]),
        .I1(\u0/u10/X [4]),
        .I2(\u0/u10/X [3]),
        .I3(\u0/u10/X [2]),
        .I4(\u0/u10/X [6]),
        .I5(\u0/u10/X [1]),
        .O(\u0/out10 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__86_i_1
       (.I0(\u0/R9 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [25]),
        .I3(\u0/uk/K_r9 [19]),
        .O(\u0/u10/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__86_i_2
       (.I0(\u0/R9 [3]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [47]),
        .I3(\u0/uk/K_r9 [41]),
        .O(\u0/u10/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__86_i_3
       (.I0(\u0/R9 [2]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [13]),
        .I3(\u0/uk/K_r9 [32]),
        .O(\u0/u10/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__86_i_4
       (.I0(\u0/R9 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [55]),
        .I3(\u0/uk/K_r9 [17]),
        .O(\u0/u10/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__86_i_5
       (.I0(\u0/R9 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [53]),
        .I3(\u0/uk/K_r9 [47]),
        .O(\u0/u10/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__86_i_6
       (.I0(\u0/R9 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r9 [34]),
        .I3(\u0/uk/K_r9 [53]),
        .O(\u0/u10/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__87
       (.I0(\u0/u11/X [41]),
        .I1(\u0/u11/X [40]),
        .I2(\u0/u11/X [39]),
        .I3(\u0/u11/X [38]),
        .I4(\u0/u11/X [42]),
        .I5(\u0/u11/X [37]),
        .O(\u0/out11 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__87_i_1
       (.I0(\u0/R10_reg_n_0_[28] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [45]),
        .I3(\u0/uk/K_r10 [36]),
        .O(\u0/u11/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__87_i_2
       (.I0(\u0/R10_reg_n_0_[27] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [30]),
        .I3(\u0/uk/K_r10 [49]),
        .O(\u0/u11/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__87_i_3
       (.I0(\u0/R10_reg_n_0_[26] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [21]),
        .I3(\u0/uk/K_r10 [16]),
        .O(\u0/u11/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__87_i_4
       (.I0(\u0/R10_reg_n_0_[25] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [36]),
        .I3(\u0/uk/K_r10 [0]),
        .O(\u0/u11/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__87_i_5
       (.I0(\u0/R10_reg_n_0_[29] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [9]),
        .I3(\u0/uk/K_r10 [28]),
        .O(\u0/u11/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__87_i_6
       (.I0(\u0/R10_reg_n_0_[24] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [1]),
        .I3(\u0/uk/K_r10 [51]),
        .O(\u0/u11/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__88
       (.I0(\u0/u11/X [17]),
        .I1(\u0/u11/X [16]),
        .I2(\u0/u11/X [15]),
        .I3(\u0/u11/X [14]),
        .I4(\u0/u11/X [18]),
        .I5(\u0/u11/X [13]),
        .O(\u0/out11 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__88_i_1
       (.I0(\u0/R10_reg_n_0_[12] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [18]),
        .I3(\u0/uk/K_r10 [41]),
        .O(\u0/u11/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__88_i_2
       (.I0(\u0/R10_reg_n_0_[11] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [3]),
        .I3(\u0/uk/K_r10 [26]),
        .O(\u0/u11/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__88_i_3
       (.I0(\u0/R10_reg_n_0_ ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [34]),
        .I3(\u0/uk/K_r10 [25]),
        .O(\u0/u11/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__88_i_4
       (.I0(\u0/R10_reg_n_0_[9] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [26]),
        .I3(\u0/uk/K_r10 [17]),
        .O(\u0/u11/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__88_i_5
       (.I0(\u0/R10_reg_n_0_[13] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [6]),
        .I3(\u0/uk/K_r10 [54]),
        .O(\u0/u11/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__88_i_6
       (.I0(\u0/R10_reg_n_0_[8] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [54]),
        .I3(\u0/uk/K_r10 [20]),
        .O(\u0/u11/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__89
       (.I0(\u0/u11/X [35]),
        .I1(\u0/u11/X [34]),
        .I2(\u0/u11/X [33]),
        .I3(\u0/u11/X [32]),
        .I4(\u0/u11/X [36]),
        .I5(\u0/u11/X [31]),
        .O(\u0/out11 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__89_i_1
       (.I0(\u0/R10_reg_n_0_[24] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [38]),
        .I3(\u0/uk/K_r10 [29]),
        .O(\u0/u11/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__89_i_2
       (.I0(\u0/R10_reg_n_0_[23] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [8]),
        .I3(\u0/uk/K_r10 [31]),
        .O(\u0/u11/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__89_i_3
       (.I0(\u0/R10_reg_n_0_[22] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [50]),
        .I3(\u0/uk/K_r10 [14]),
        .O(\u0/u11/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__89_i_4
       (.I0(\u0/R10_reg_n_0_[21] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [28]),
        .I3(\u0/uk/K_r10 [23]),
        .O(\u0/u11/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__89_i_5
       (.I0(\u0/R10_reg_n_0_[25] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [29]),
        .I3(\u0/uk/K_r10 [52]),
        .O(\u0/u11/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__89_i_6
       (.I0(\u0/R10_reg_n_0_[20] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [44]),
        .I3(\u0/uk/K_r10 [8]),
        .O(\u0/u11/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__8_i_1
       (.I0(\u0/R0 [12]),
        .I1(decrypt),
        .I2(\u0/uk/p_3_in ),
        .I3(\u0/uk/p_11_in ),
        .O(\u0/u1/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__8_i_2
       (.I0(\u0/R0 [11]),
        .I1(decrypt),
        .I2(\u0/uk/p_13_in ),
        .I3(\u0/uk/p_2_in ),
        .O(\u0/u1/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__8_i_3
       (.I0(\u0/R0 [10]),
        .I1(decrypt),
        .I2(\u0/uk/p_8_in ),
        .I3(\u0/uk/K_r0_reg_n_0_[19] ),
        .O(\u0/u1/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__8_i_4
       (.I0(\u0/R0 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r0_reg_n_0_[32] ),
        .I3(\u0/uk/p_14_in ),
        .O(\u0/u1/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__8_i_5
       (.I0(\u0/R0 [13]),
        .I1(decrypt),
        .I2(\u0/uk/p_38_in ),
        .I3(\u0/uk/p_4_in ),
        .O(\u0/u1/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__8_i_6
       (.I0(\u0/R0 [8]),
        .I1(decrypt),
        .I2(\u0/uk/p_11_in ),
        .I3(\u0/uk/p_12_in ),
        .O(\u0/u1/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__9
       (.I0(\u0/u1/X [35]),
        .I1(\u0/u1/X [34]),
        .I2(\u0/u1/X [33]),
        .I3(\u0/u1/X [32]),
        .I4(\u0/u1/X [36]),
        .I5(\u0/u1/X [31]),
        .O(\u0/out1 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__90
       (.I0(\u0/u11/X [11]),
        .I1(\u0/u11/X [10]),
        .I2(\u0/u11/X [9]),
        .I3(\u0/u11/X [8]),
        .I4(\u0/u11/X [12]),
        .I5(\u0/u11/X [7]),
        .O(\u0/out11 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__90_i_1
       (.I0(\u0/R10_reg_n_0_[8] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [40]),
        .I3(\u0/uk/K_r10 [6]),
        .O(\u0/u11/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__90_i_2
       (.I0(\u0/R10_reg_n_0_[7] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [17]),
        .I3(\u0/uk/K_r10 [40]),
        .O(\u0/u11/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__90_i_3
       (.I0(\u0/R10_reg_n_0_[6] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [55]),
        .I3(\u0/uk/K_r10 [46]),
        .O(\u0/u11/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__90_i_4
       (.I0(\u0/R10_reg_n_0_[5] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [32]),
        .I3(\u0/uk/K_r10 [55]),
        .O(\u0/u11/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__90_i_5
       (.I0(\u0/R10_reg_n_0_[9] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [20]),
        .I3(\u0/uk/K_r10 [11]),
        .O(\u0/u11/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__90_i_6
       (.I0(\u0/R10_reg_n_0_[4] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [53]),
        .I3(\u0/uk/K_r10 [19]),
        .O(\u0/u11/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__91
       (.I0(\u0/u11/X [47]),
        .I1(\u0/u11/X [46]),
        .I2(\u0/u11/X [45]),
        .I3(\u0/u11/X [44]),
        .I4(\u0/u11/X [48]),
        .I5(\u0/u11/X [43]),
        .O(\u0/out11 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__91_i_1
       (.I0(\u0/R10_reg_n_0_[32] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [37]),
        .I3(\u0/uk/K_r10 [1]),
        .O(\u0/u11/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__91_i_2
       (.I0(\u0/R10_reg_n_0_[31] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [0]),
        .I3(\u0/uk/K_r10 [50]),
        .O(\u0/u11/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__91_i_3
       (.I0(\u0/R10_reg_n_0_[30] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [43]),
        .I3(\u0/uk/K_r10 [7]),
        .O(\u0/u11/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__91_i_4
       (.I0(\u0/R10_reg_n_0_[29] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [42]),
        .I3(\u0/uk/K_r10 [37]),
        .O(\u0/u11/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__91_i_5
       (.I0(\u0/R10_reg_n_0_[1] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [31]),
        .I3(\u0/uk/K_r10 [22]),
        .O(\u0/u11/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__91_i_6
       (.I0(\u0/R10_reg_n_0_[28] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [15]),
        .I3(\u0/uk/K_r10 [38]),
        .O(\u0/u11/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2D6317E492AD994B)) 
    g0_b0__92
       (.I0(\u0/u11/X [23]),
        .I1(\u0/u11/X [22]),
        .I2(\u0/u11/X [21]),
        .I3(\u0/u11/X [20]),
        .I4(\u0/u11/X [24]),
        .I5(\u0/u11/X [19]),
        .O(\u0/out11 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__92_i_1
       (.I0(\u0/R10_reg_n_0_[16] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [41]),
        .I3(\u0/uk/K_r10 [32]),
        .O(\u0/u11/X [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__92_i_2
       (.I0(\u0/R10_reg_n_0_[15] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [33]),
        .I3(\u0/uk/K_r10 [24]),
        .O(\u0/u11/X [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__92_i_3
       (.I0(\u0/R10_reg_n_0_[14] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [25]),
        .I3(\u0/uk/K_r10 [48]),
        .O(\u0/u11/X [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__92_i_4
       (.I0(\u0/R10_reg_n_0_[13] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [24]),
        .I3(\u0/uk/K_r10 [47]),
        .O(\u0/u11/X [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__92_i_5
       (.I0(\u0/R10_reg_n_0_[17] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [46]),
        .I3(\u0/uk/K_r10 [12]),
        .O(\u0/u11/X [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__92_i_6
       (.I0(\u0/R10_reg_n_0_[12] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [5]),
        .I3(\u0/uk/K_r10 [53]),
        .O(\u0/u11/X [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCA992B6C35E29E58)) 
    g0_b0__93
       (.I0(\u0/u11/X [29]),
        .I1(\u0/u11/X [28]),
        .I2(\u0/u11/X [27]),
        .I3(\u0/u11/X [26]),
        .I4(\u0/u11/X [30]),
        .I5(\u0/u11/X [25]),
        .O(\u0/out11 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__93_i_1
       (.I0(\u0/R10_reg_n_0_[20] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [22]),
        .I3(\u0/uk/K_r10 [45]),
        .O(\u0/u11/X [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__93_i_2
       (.I0(\u0/R10_reg_n_0_[19] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [7]),
        .I3(\u0/uk/K_r10 [2]),
        .O(\u0/u11/X [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__93_i_3
       (.I0(\u0/R10_reg_n_0_[18] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [51]),
        .I3(\u0/uk/K_r10 [15]),
        .O(\u0/u11/X [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__93_i_4
       (.I0(\u0/R10_reg_n_0_[17] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [2]),
        .I3(\u0/uk/K_r10 [21]),
        .O(\u0/u11/X [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__93_i_5
       (.I0(\u0/R10_reg_n_0_[21] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [23]),
        .I3(\u0/uk/K_r10 [42]),
        .O(\u0/u11/X [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__93_i_6
       (.I0(\u0/R10_reg_n_0_[16] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [35]),
        .I3(\u0/uk/K_r10 [30]),
        .O(\u0/u11/X [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E15D9278C6B16C)) 
    g0_b0__94
       (.I0(\u0/u11/X [5]),
        .I1(\u0/u11/X [4]),
        .I2(\u0/u11/X [3]),
        .I3(\u0/u11/X [2]),
        .I4(\u0/u11/X [6]),
        .I5(\u0/u11/X [1]),
        .O(\u0/out11 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__94_i_1
       (.I0(\u0/R10_reg_n_0_[4] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [39]),
        .I3(\u0/uk/K_r10 [5]),
        .O(\u0/u11/X [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__94_i_2
       (.I0(\u0/R10_reg_n_0_[3] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [4]),
        .I3(\u0/uk/K_r10 [27]),
        .O(\u0/u11/X [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__94_i_3
       (.I0(\u0/R10_reg_n_0_[2] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [27]),
        .I3(\u0/uk/K_r10 [18]),
        .O(\u0/u11/X [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__94_i_4
       (.I0(\u0/R10_reg_n_0_[1] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [12]),
        .I3(\u0/uk/K_r10 [3]),
        .O(\u0/u11/X [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__94_i_5
       (.I0(\u0/R10_reg_n_0_[5] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [10]),
        .I3(\u0/uk/K_r10 [33]),
        .O(\u0/u11/X [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__94_i_6
       (.I0(\u0/R10_reg_n_0_[32] ),
        .I1(decrypt),
        .I2(\u0/uk/K_r10 [48]),
        .I3(\u0/uk/K_r10 [39]),
        .O(\u0/u11/X [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B96626D266D9D92)) 
    g0_b0__95
       (.I0(\u0/u12/X [41]),
        .I1(\u0/u12/X [40]),
        .I2(\u0/u12/X [39]),
        .I3(\u0/u12/X [38]),
        .I4(\u0/u12/X [42]),
        .I5(\u0/u12/X [37]),
        .O(\u0/out12 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__95_i_1
       (.I0(\u0/R11 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [0]),
        .I3(\u0/uk/K_r11 [22]),
        .O(\u0/u12/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__95_i_2
       (.I0(\u0/R11 [27]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [44]),
        .I3(\u0/uk/K_r11 [35]),
        .O(\u0/u12/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__95_i_3
       (.I0(\u0/R11 [26]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [35]),
        .I3(\u0/uk/K_r11 [2]),
        .O(\u0/u12/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__95_i_4
       (.I0(\u0/R11 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [50]),
        .I3(\u0/uk/K_r11 [45]),
        .O(\u0/u12/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__95_i_5
       (.I0(\u0/R11 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [23]),
        .I3(\u0/uk/K_r11 [14]),
        .O(\u0/u12/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__95_i_6
       (.I0(\u0/R11 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [15]),
        .I3(\u0/uk/K_r11 [37]),
        .O(\u0/u12/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3AA59369E41B1BE4)) 
    g0_b0__96
       (.I0(\u0/u12/X [17]),
        .I1(\u0/u12/X [16]),
        .I2(\u0/u12/X [15]),
        .I3(\u0/u12/X [14]),
        .I4(\u0/u12/X [18]),
        .I5(\u0/u12/X [13]),
        .O(\u0/out12 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__96_i_1
       (.I0(\u0/R11 [12]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [32]),
        .I3(\u0/uk/K_r11 [27]),
        .O(\u0/u12/X [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__96_i_2
       (.I0(\u0/R11 [11]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [17]),
        .I3(\u0/uk/K_r11 [12]),
        .O(\u0/u12/X [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__96_i_3
       (.I0(\u0/R11 [10]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [48]),
        .I3(\u0/uk/K_r11 [11]),
        .O(\u0/u12/X [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__96_i_4
       (.I0(\u0/R11 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [40]),
        .I3(\u0/uk/K_r11 [3]),
        .O(\u0/u12/X [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__96_i_5
       (.I0(\u0/R11 [13]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [20]),
        .I3(\u0/uk/K_r11 [40]),
        .O(\u0/u12/X [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__96_i_6
       (.I0(\u0/R11 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [11]),
        .I3(\u0/uk/K_r11 [6]),
        .O(\u0/u12/X [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8D72718D66D2E61A)) 
    g0_b0__97
       (.I0(\u0/u12/X [35]),
        .I1(\u0/u12/X [34]),
        .I2(\u0/u12/X [33]),
        .I3(\u0/u12/X [32]),
        .I4(\u0/u12/X [36]),
        .I5(\u0/u12/X [31]),
        .O(\u0/out12 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__97_i_1
       (.I0(\u0/R11 [24]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [52]),
        .I3(\u0/uk/K_r11 [15]),
        .O(\u0/u12/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__97_i_2
       (.I0(\u0/R11 [23]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [22]),
        .I3(\u0/uk/K_r11 [44]),
        .O(\u0/u12/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__97_i_3
       (.I0(\u0/R11 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [9]),
        .I3(\u0/uk/K_r11 [0]),
        .O(\u0/u12/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__97_i_4
       (.I0(\u0/R11 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [42]),
        .I3(\u0/uk/K_r11 [9]),
        .O(\u0/u12/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__97_i_5
       (.I0(\u0/R11 [25]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [43]),
        .I3(\u0/uk/K_r11 [38]),
        .O(\u0/u12/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__97_i_6
       (.I0(\u0/R11 [20]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [31]),
        .I3(\u0/uk/K_r11 [49]),
        .O(\u0/u12/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA539B1CCE41B4B63)) 
    g0_b0__98
       (.I0(\u0/u12/X [11]),
        .I1(\u0/u12/X [10]),
        .I2(\u0/u12/X [9]),
        .I3(\u0/u12/X [8]),
        .I4(\u0/u12/X [12]),
        .I5(\u0/u12/X [7]),
        .O(\u0/out12 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__98_i_1
       (.I0(\u0/R11 [8]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [54]),
        .I3(\u0/uk/K_r11 [17]),
        .O(\u0/u12/X [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__98_i_2
       (.I0(\u0/R11 [7]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [6]),
        .I3(\u0/uk/K_r11 [26]),
        .O(\u0/u12/X [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__98_i_3
       (.I0(\u0/R11 [6]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [12]),
        .I3(\u0/uk/K_r11 [32]),
        .O(\u0/u12/X [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__98_i_4
       (.I0(\u0/R11 [5]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [46]),
        .I3(\u0/uk/K_r11 [41]),
        .O(\u0/u12/X [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__98_i_5
       (.I0(\u0/R11 [9]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [34]),
        .I3(\u0/uk/K_r11 [54]),
        .O(\u0/u12/X [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__98_i_6
       (.I0(\u0/R11 [4]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [10]),
        .I3(\u0/uk/K_r11 [5]),
        .O(\u0/u12/X [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB58A781B4A6796E1)) 
    g0_b0__99
       (.I0(\u0/u12/X [47]),
        .I1(\u0/u12/X [46]),
        .I2(\u0/u12/X [45]),
        .I3(\u0/u12/X [44]),
        .I4(\u0/u12/X [48]),
        .I5(\u0/u12/X [43]),
        .O(\u0/out12 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__99_i_1
       (.I0(\u0/R11 [32]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [51]),
        .I3(\u0/uk/K_r11 [42]),
        .O(\u0/u12/X [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__99_i_2
       (.I0(\u0/R11 [31]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [14]),
        .I3(\u0/uk/K_r11 [36]),
        .O(\u0/u12/X [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__99_i_3
       (.I0(\u0/R11 [30]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [2]),
        .I3(\u0/uk/K_r11 [52]),
        .O(\u0/u12/X [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__99_i_4
       (.I0(\u0/R11 [29]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [1]),
        .I3(\u0/uk/K_r11 [23]),
        .O(\u0/u12/X [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__99_i_5
       (.I0(\u0/R11 [1]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [45]),
        .I3(\u0/uk/K_r11 [8]),
        .O(\u0/u12/X [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__99_i_6
       (.I0(\u0/R11 [28]),
        .I1(decrypt),
        .I2(\u0/uk/K_r11 [29]),
        .I3(\u0/uk/K_r11 [51]),
        .O(\u0/u12/X [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__9_i_1
       (.I0(\u0/R0 [24]),
        .I1(decrypt),
        .I2(\u0/uk/p_29_in ),
        .I3(\u0/uk/p_24_in ),
        .O(\u0/u1/X [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__9_i_2
       (.I0(\u0/R0 [23]),
        .I1(decrypt),
        .I2(\u0/uk/p_27_in ),
        .I3(\u0/uk/p_28_in ),
        .O(\u0/u1/X [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__9_i_3
       (.I0(\u0/R0 [22]),
        .I1(decrypt),
        .I2(\u0/uk/K_r0_reg_n_0_[31] ),
        .I3(\u0/uk/p_26_in ),
        .O(\u0/u1/X [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__9_i_4
       (.I0(\u0/R0 [21]),
        .I1(decrypt),
        .I2(\u0/uk/K_r0_reg_n_0_[36] ),
        .I3(\u0/uk/p_25_in ),
        .O(\u0/u1/X [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__9_i_5
       (.I0(\u0/R0 [25]),
        .I1(decrypt),
        .I2(\u0/uk/p_26_in ),
        .I3(\u0/uk/p_27_in ),
        .O(\u0/u1/X [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0__9_i_6
       (.I0(\u0/R0 [20]),
        .I1(decrypt),
        .I2(\u0/uk/p_24_in ),
        .I3(\u0/uk/K_r0_reg_n_0_ ),
        .O(\u0/u1/X [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0_i_1
       (.I0(\u0/IP [60]),
        .I1(decrypt),
        .I2(\u0/key_r [42]),
        .I3(\u0/key_r [35]),
        .O(\u0/u0/X [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0_i_2
       (.I0(\u0/IP [59]),
        .I1(decrypt),
        .I2(\u0/key_r [0]),
        .I3(\u0/key_r [52]),
        .O(\u0/u0/X [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0_i_3
       (.I0(\u0/IP [58]),
        .I1(decrypt),
        .I2(\u0/key_r [22]),
        .I3(\u0/key_r [15]),
        .O(\u0/u0/X [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0_i_4
       (.I0(\u0/IP [57]),
        .I1(decrypt),
        .I2(\u0/key_r [37]),
        .I3(\u0/key_r [30]),
        .O(\u0/u0/X [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0_i_5
       (.I0(\u0/IP [61]),
        .I1(decrypt),
        .I2(\u0/key_r [38]),
        .I3(\u0/key_r [31]),
        .O(\u0/u0/X [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h569A)) 
    g0_b0_i_6
       (.I0(\u0/IP [56]),
        .I1(decrypt),
        .I2(\u0/key_r [2]),
        .I3(\u0/key_r [50]),
        .O(\u0/u0/X [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1
       (.I0(\u0/u0/X [41]),
        .I1(\u0/u0/X [40]),
        .I2(\u0/u0/X [39]),
        .I3(\u0/u0/X [38]),
        .I4(\u0/u0/X [42]),
        .I5(\u0/u0/X [37]),
        .O(\u0/out0 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__0
       (.I0(\u0/u0/X [17]),
        .I1(\u0/u0/X [16]),
        .I2(\u0/u0/X [15]),
        .I3(\u0/u0/X [14]),
        .I4(\u0/u0/X [18]),
        .I5(\u0/u0/X [13]),
        .O(\u0/out0 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__1
       (.I0(\u0/u0/X [35]),
        .I1(\u0/u0/X [34]),
        .I2(\u0/u0/X [33]),
        .I3(\u0/u0/X [32]),
        .I4(\u0/u0/X [36]),
        .I5(\u0/u0/X [31]),
        .O(\u0/out0 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__10
       (.I0(\u0/u1/X [11]),
        .I1(\u0/u1/X [10]),
        .I2(\u0/u1/X [9]),
        .I3(\u0/u1/X [8]),
        .I4(\u0/u1/X [12]),
        .I5(\u0/u1/X [7]),
        .O(\u0/out1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__100
       (.I0(\u0/u12/X [23]),
        .I1(\u0/u12/X [22]),
        .I2(\u0/u12/X [21]),
        .I3(\u0/u12/X [20]),
        .I4(\u0/u12/X [24]),
        .I5(\u0/u12/X [19]),
        .O(\u0/out12 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__101
       (.I0(\u0/u12/X [29]),
        .I1(\u0/u12/X [28]),
        .I2(\u0/u12/X [27]),
        .I3(\u0/u12/X [26]),
        .I4(\u0/u12/X [30]),
        .I5(\u0/u12/X [25]),
        .O(\u0/out12 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__102
       (.I0(\u0/u12/X [5]),
        .I1(\u0/u12/X [4]),
        .I2(\u0/u12/X [3]),
        .I3(\u0/u12/X [2]),
        .I4(\u0/u12/X [6]),
        .I5(\u0/u12/X [1]),
        .O(\u0/out12 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__103
       (.I0(\u0/u13/X [41]),
        .I1(\u0/u13/X [40]),
        .I2(\u0/u13/X [39]),
        .I3(\u0/u13/X [38]),
        .I4(\u0/u13/X [42]),
        .I5(\u0/u13/X [37]),
        .O(\u0/out13 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__104
       (.I0(\u0/u13/X [17]),
        .I1(\u0/u13/X [16]),
        .I2(\u0/u13/X [15]),
        .I3(\u0/u13/X [14]),
        .I4(\u0/u13/X [18]),
        .I5(\u0/u13/X [13]),
        .O(\u0/out13 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__105
       (.I0(\u0/u13/X [35]),
        .I1(\u0/u13/X [34]),
        .I2(\u0/u13/X [33]),
        .I3(\u0/u13/X [32]),
        .I4(\u0/u13/X [36]),
        .I5(\u0/u13/X [31]),
        .O(\u0/out13 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__106
       (.I0(\u0/u13/X [11]),
        .I1(\u0/u13/X [10]),
        .I2(\u0/u13/X [9]),
        .I3(\u0/u13/X [8]),
        .I4(\u0/u13/X [12]),
        .I5(\u0/u13/X [7]),
        .O(\u0/out13 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__107
       (.I0(\u0/u13/X [47]),
        .I1(\u0/u13/X [46]),
        .I2(\u0/u13/X [45]),
        .I3(\u0/u13/X [44]),
        .I4(\u0/u13/X [48]),
        .I5(\u0/u13/X [43]),
        .O(\u0/out13 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__108
       (.I0(\u0/u13/X [23]),
        .I1(\u0/u13/X [22]),
        .I2(\u0/u13/X [21]),
        .I3(\u0/u13/X [20]),
        .I4(\u0/u13/X [24]),
        .I5(\u0/u13/X [19]),
        .O(\u0/out13 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__109
       (.I0(\u0/u13/X [29]),
        .I1(\u0/u13/X [28]),
        .I2(\u0/u13/X [27]),
        .I3(\u0/u13/X [26]),
        .I4(\u0/u13/X [30]),
        .I5(\u0/u13/X [25]),
        .O(\u0/out13 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__11
       (.I0(\u0/u1/X [47]),
        .I1(\u0/u1/X [46]),
        .I2(\u0/u1/X [45]),
        .I3(\u0/u1/X [44]),
        .I4(\u0/u1/X [48]),
        .I5(\u0/u1/X [43]),
        .O(\u0/out1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__110
       (.I0(\u0/u13/X [5]),
        .I1(\u0/u13/X [4]),
        .I2(\u0/u13/X [3]),
        .I3(\u0/u13/X [2]),
        .I4(\u0/u13/X [6]),
        .I5(\u0/u13/X [1]),
        .O(\u0/out13 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__111
       (.I0(\u0/u14/X [41]),
        .I1(\u0/u14/X [40]),
        .I2(\u0/u14/X [39]),
        .I3(\u0/u14/X [38]),
        .I4(\u0/u14/X [42]),
        .I5(\u0/u14/X [37]),
        .O(\u0/out14 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__112
       (.I0(\u0/u14/X [17]),
        .I1(\u0/u14/X [16]),
        .I2(\u0/u14/X [15]),
        .I3(\u0/u14/X [14]),
        .I4(\u0/u14/X [18]),
        .I5(\u0/u14/X [13]),
        .O(\u0/out14 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__113
       (.I0(\u0/u14/X [35]),
        .I1(\u0/u14/X [34]),
        .I2(\u0/u14/X [33]),
        .I3(\u0/u14/X [32]),
        .I4(\u0/u14/X [36]),
        .I5(\u0/u14/X [31]),
        .O(\u0/out14 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__114
       (.I0(\u0/u14/X [11]),
        .I1(\u0/u14/X [10]),
        .I2(\u0/u14/X [9]),
        .I3(\u0/u14/X [8]),
        .I4(\u0/u14/X [12]),
        .I5(\u0/u14/X [7]),
        .O(\u0/out14 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__115
       (.I0(\u0/u14/X [47]),
        .I1(\u0/u14/X [46]),
        .I2(\u0/u14/X [45]),
        .I3(\u0/u14/X [44]),
        .I4(\u0/u14/X [48]),
        .I5(\u0/u14/X [43]),
        .O(\u0/out14 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__116
       (.I0(\u0/u14/X [23]),
        .I1(\u0/u14/X [22]),
        .I2(\u0/u14/X [21]),
        .I3(\u0/u14/X [20]),
        .I4(\u0/u14/X [24]),
        .I5(\u0/u14/X [19]),
        .O(\u0/out14 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__117
       (.I0(\u0/u14/X [29]),
        .I1(\u0/u14/X [28]),
        .I2(\u0/u14/X [27]),
        .I3(\u0/u14/X [26]),
        .I4(\u0/u14/X [30]),
        .I5(\u0/u14/X [25]),
        .O(\u0/out14 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__118
       (.I0(\u0/u14/X [5]),
        .I1(\u0/u14/X [4]),
        .I2(\u0/u14/X [3]),
        .I3(\u0/u14/X [2]),
        .I4(\u0/u14/X [6]),
        .I5(\u0/u14/X [1]),
        .O(\u0/out14 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__119
       (.I0(\u0/u15/X [41]),
        .I1(\u0/u15/X [40]),
        .I2(\u0/u15/X [39]),
        .I3(\u0/u15/X [38]),
        .I4(\u0/u15/X [42]),
        .I5(\u0/u15/X [37]),
        .O(\u0/out15 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__12
       (.I0(\u0/u1/X [23]),
        .I1(\u0/u1/X [22]),
        .I2(\u0/u1/X [21]),
        .I3(\u0/u1/X [20]),
        .I4(\u0/u1/X [24]),
        .I5(\u0/u1/X [19]),
        .O(\u0/out1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__120
       (.I0(\u0/u15/X [17]),
        .I1(\u0/u15/X [16]),
        .I2(\u0/u15/X [15]),
        .I3(\u0/u15/X [14]),
        .I4(\u0/u15/X [18]),
        .I5(\u0/u15/X [13]),
        .O(\u0/out15 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__121
       (.I0(\u0/u15/X [35]),
        .I1(\u0/u15/X [34]),
        .I2(\u0/u15/X [33]),
        .I3(\u0/u15/X [32]),
        .I4(\u0/u15/X [36]),
        .I5(\u0/u15/X [31]),
        .O(\u0/out15 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__122
       (.I0(\u0/u15/X [11]),
        .I1(\u0/u15/X [10]),
        .I2(\u0/u15/X [9]),
        .I3(\u0/u15/X [8]),
        .I4(\u0/u15/X [12]),
        .I5(\u0/u15/X [7]),
        .O(\u0/out15 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__123
       (.I0(\u0/u15/X [47]),
        .I1(\u0/u15/X [46]),
        .I2(\u0/u15/X [45]),
        .I3(\u0/u15/X [44]),
        .I4(\u0/u15/X [48]),
        .I5(\u0/u15/X [43]),
        .O(\u0/out15 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__124
       (.I0(\u0/u15/X [23]),
        .I1(\u0/u15/X [22]),
        .I2(\u0/u15/X [21]),
        .I3(\u0/u15/X [20]),
        .I4(\u0/u15/X [24]),
        .I5(\u0/u15/X [19]),
        .O(\u0/out15 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__125
       (.I0(\u0/u15/X [29]),
        .I1(\u0/u15/X [28]),
        .I2(\u0/u15/X [27]),
        .I3(\u0/u15/X [26]),
        .I4(\u0/u15/X [30]),
        .I5(\u0/u15/X [25]),
        .O(\u0/out15 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__126
       (.I0(\u0/u15/X [5]),
        .I1(\u0/u15/X [4]),
        .I2(\u0/u15/X [3]),
        .I3(\u0/u15/X [2]),
        .I4(\u0/u15/X [6]),
        .I5(\u0/u15/X [1]),
        .O(\u0/out15 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__127
       (.I0(\u1/u0/X [41]),
        .I1(\u1/u0/X [40]),
        .I2(\u1/u0/X [39]),
        .I3(\u1/u0/X [38]),
        .I4(\u1/u0/X [42]),
        .I5(\u1/u0/X [37]),
        .O(\u1/out0 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__128
       (.I0(\u1/u0/X [17]),
        .I1(\u1/u0/X [16]),
        .I2(\u1/u0/X [15]),
        .I3(\u1/u0/X [14]),
        .I4(\u1/u0/X [18]),
        .I5(\u1/u0/X [13]),
        .O(\u1/out0 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__129
       (.I0(\u1/u0/X [35]),
        .I1(\u1/u0/X [34]),
        .I2(\u1/u0/X [33]),
        .I3(\u1/u0/X [32]),
        .I4(\u1/u0/X [36]),
        .I5(\u1/u0/X [31]),
        .O(\u1/out0 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__13
       (.I0(\u0/u1/X [29]),
        .I1(\u0/u1/X [28]),
        .I2(\u0/u1/X [27]),
        .I3(\u0/u1/X [26]),
        .I4(\u0/u1/X [30]),
        .I5(\u0/u1/X [25]),
        .O(\u0/out1 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__130
       (.I0(\u1/u0/X [11]),
        .I1(\u1/u0/X [10]),
        .I2(\u1/u0/X [9]),
        .I3(\u1/u0/X [8]),
        .I4(\u1/u0/X [12]),
        .I5(\u1/u0/X [7]),
        .O(\u1/out0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__131
       (.I0(\u1/u0/X [47]),
        .I1(\u1/u0/X [46]),
        .I2(\u1/u0/X [45]),
        .I3(\u1/u0/X [44]),
        .I4(\u1/u0/X [48]),
        .I5(\u1/u0/X [43]),
        .O(\u1/out0 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__132
       (.I0(\u1/u0/X [23]),
        .I1(\u1/u0/X [22]),
        .I2(\u1/u0/X [21]),
        .I3(\u1/u0/X [20]),
        .I4(\u1/u0/X [24]),
        .I5(\u1/u0/X [19]),
        .O(\u1/out0 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__133
       (.I0(\u1/u0/X [29]),
        .I1(\u1/u0/X [28]),
        .I2(\u1/u0/X [27]),
        .I3(\u1/u0/X [26]),
        .I4(\u1/u0/X [30]),
        .I5(\u1/u0/X [25]),
        .O(\u1/out0 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__134
       (.I0(\u1/u0/X [5]),
        .I1(\u1/u0/X [4]),
        .I2(\u1/u0/X [3]),
        .I3(\u1/u0/X [2]),
        .I4(\u1/u0/X [6]),
        .I5(\u1/u0/X [1]),
        .O(\u1/out0 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__135
       (.I0(\u1/u1/X [41]),
        .I1(\u1/u1/X [40]),
        .I2(\u1/u1/X [39]),
        .I3(\u1/u1/X [38]),
        .I4(\u1/u1/X [42]),
        .I5(\u1/u1/X [37]),
        .O(\u1/out1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__136
       (.I0(\u1/u1/X [17]),
        .I1(\u1/u1/X [16]),
        .I2(\u1/u1/X [15]),
        .I3(\u1/u1/X [14]),
        .I4(\u1/u1/X [18]),
        .I5(\u1/u1/X [13]),
        .O(\u1/out1 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__137
       (.I0(\u1/u1/X [35]),
        .I1(\u1/u1/X [34]),
        .I2(\u1/u1/X [33]),
        .I3(\u1/u1/X [32]),
        .I4(\u1/u1/X [36]),
        .I5(\u1/u1/X [31]),
        .O(\u1/out1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__138
       (.I0(\u1/u1/X [11]),
        .I1(\u1/u1/X [10]),
        .I2(\u1/u1/X [9]),
        .I3(\u1/u1/X [8]),
        .I4(\u1/u1/X [12]),
        .I5(\u1/u1/X [7]),
        .O(\u1/out1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__139
       (.I0(\u1/u1/X [47]),
        .I1(\u1/u1/X [46]),
        .I2(\u1/u1/X [45]),
        .I3(\u1/u1/X [44]),
        .I4(\u1/u1/X [48]),
        .I5(\u1/u1/X [43]),
        .O(\u1/out1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__14
       (.I0(\u0/u1/X [5]),
        .I1(\u0/u1/X [4]),
        .I2(\u0/u1/X [3]),
        .I3(\u0/u1/X [2]),
        .I4(\u0/u1/X [6]),
        .I5(\u0/u1/X [1]),
        .O(\u0/out1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__140
       (.I0(\u1/u1/X [23]),
        .I1(\u1/u1/X [22]),
        .I2(\u1/u1/X [21]),
        .I3(\u1/u1/X [20]),
        .I4(\u1/u1/X [24]),
        .I5(\u1/u1/X [19]),
        .O(\u1/out1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__141
       (.I0(\u1/u1/X [29]),
        .I1(\u1/u1/X [28]),
        .I2(\u1/u1/X [27]),
        .I3(\u1/u1/X [26]),
        .I4(\u1/u1/X [30]),
        .I5(\u1/u1/X [25]),
        .O(\u1/out1 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__142
       (.I0(\u1/u1/X [5]),
        .I1(\u1/u1/X [4]),
        .I2(\u1/u1/X [3]),
        .I3(\u1/u1/X [2]),
        .I4(\u1/u1/X [6]),
        .I5(\u1/u1/X [1]),
        .O(\u1/out1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__143
       (.I0(\u1/u2/X [41]),
        .I1(\u1/u2/X [40]),
        .I2(\u1/u2/X [39]),
        .I3(\u1/u2/X [38]),
        .I4(\u1/u2/X [42]),
        .I5(\u1/u2/X [37]),
        .O(\u1/out2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__144
       (.I0(\u1/u2/X [17]),
        .I1(\u1/u2/X [16]),
        .I2(\u1/u2/X [15]),
        .I3(\u1/u2/X [14]),
        .I4(\u1/u2/X [18]),
        .I5(\u1/u2/X [13]),
        .O(\u1/out2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__145
       (.I0(\u1/u2/X [35]),
        .I1(\u1/u2/X [34]),
        .I2(\u1/u2/X [33]),
        .I3(\u1/u2/X [32]),
        .I4(\u1/u2/X [36]),
        .I5(\u1/u2/X [31]),
        .O(\u1/out2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__146
       (.I0(\u1/u2/X [11]),
        .I1(\u1/u2/X [10]),
        .I2(\u1/u2/X [9]),
        .I3(\u1/u2/X [8]),
        .I4(\u1/u2/X [12]),
        .I5(\u1/u2/X [7]),
        .O(\u1/out2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__147
       (.I0(\u1/u2/X [47]),
        .I1(\u1/u2/X [46]),
        .I2(\u1/u2/X [45]),
        .I3(\u1/u2/X [44]),
        .I4(\u1/u2/X [48]),
        .I5(\u1/u2/X [43]),
        .O(\u1/out2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__148
       (.I0(\u1/u2/X [23]),
        .I1(\u1/u2/X [22]),
        .I2(\u1/u2/X [21]),
        .I3(\u1/u2/X [20]),
        .I4(\u1/u2/X [24]),
        .I5(\u1/u2/X [19]),
        .O(\u1/out2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__149
       (.I0(\u1/u2/X [29]),
        .I1(\u1/u2/X [28]),
        .I2(\u1/u2/X [27]),
        .I3(\u1/u2/X [26]),
        .I4(\u1/u2/X [30]),
        .I5(\u1/u2/X [25]),
        .O(\u1/out2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__15
       (.I0(\u0/u2/X [41]),
        .I1(\u0/u2/X [40]),
        .I2(\u0/u2/X [39]),
        .I3(\u0/u2/X [38]),
        .I4(\u0/u2/X [42]),
        .I5(\u0/u2/X [37]),
        .O(\u0/out2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__150
       (.I0(\u1/u2/X [5]),
        .I1(\u1/u2/X [4]),
        .I2(\u1/u2/X [3]),
        .I3(\u1/u2/X [2]),
        .I4(\u1/u2/X [6]),
        .I5(\u1/u2/X [1]),
        .O(\u1/out2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__151
       (.I0(\u1/u3/X [41]),
        .I1(\u1/u3/X [40]),
        .I2(\u1/u3/X [39]),
        .I3(\u1/u3/X [38]),
        .I4(\u1/u3/X [42]),
        .I5(\u1/u3/X [37]),
        .O(\u1/out3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__152
       (.I0(\u1/u3/X [17]),
        .I1(\u1/u3/X [16]),
        .I2(\u1/u3/X [15]),
        .I3(\u1/u3/X [14]),
        .I4(\u1/u3/X [18]),
        .I5(\u1/u3/X [13]),
        .O(\u1/out3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__153
       (.I0(\u1/u3/X [35]),
        .I1(\u1/u3/X [34]),
        .I2(\u1/u3/X [33]),
        .I3(\u1/u3/X [32]),
        .I4(\u1/u3/X [36]),
        .I5(\u1/u3/X [31]),
        .O(\u1/out3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__154
       (.I0(\u1/u3/X [11]),
        .I1(\u1/u3/X [10]),
        .I2(\u1/u3/X [9]),
        .I3(\u1/u3/X [8]),
        .I4(\u1/u3/X [12]),
        .I5(\u1/u3/X [7]),
        .O(\u1/out3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__155
       (.I0(\u1/u3/X [47]),
        .I1(\u1/u3/X [46]),
        .I2(\u1/u3/X [45]),
        .I3(\u1/u3/X [44]),
        .I4(\u1/u3/X [48]),
        .I5(\u1/u3/X [43]),
        .O(\u1/out3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__156
       (.I0(\u1/u3/X [23]),
        .I1(\u1/u3/X [22]),
        .I2(\u1/u3/X [21]),
        .I3(\u1/u3/X [20]),
        .I4(\u1/u3/X [24]),
        .I5(\u1/u3/X [19]),
        .O(\u1/out3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__157
       (.I0(\u1/u3/X [29]),
        .I1(\u1/u3/X [28]),
        .I2(\u1/u3/X [27]),
        .I3(\u1/u3/X [26]),
        .I4(\u1/u3/X [30]),
        .I5(\u1/u3/X [25]),
        .O(\u1/out3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__158
       (.I0(\u1/u3/X [5]),
        .I1(\u1/u3/X [4]),
        .I2(\u1/u3/X [3]),
        .I3(\u1/u3/X [2]),
        .I4(\u1/u3/X [6]),
        .I5(\u1/u3/X [1]),
        .O(\u1/out3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__159
       (.I0(\u1/u4/X [41]),
        .I1(\u1/u4/X [40]),
        .I2(\u1/u4/X [39]),
        .I3(\u1/u4/X [38]),
        .I4(\u1/u4/X [42]),
        .I5(\u1/u4/X [37]),
        .O(\u1/out4 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__16
       (.I0(\u0/u2/X [17]),
        .I1(\u0/u2/X [16]),
        .I2(\u0/u2/X [15]),
        .I3(\u0/u2/X [14]),
        .I4(\u0/u2/X [18]),
        .I5(\u0/u2/X [13]),
        .O(\u0/out2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__160
       (.I0(\u1/u4/X [17]),
        .I1(\u1/u4/X [16]),
        .I2(\u1/u4/X [15]),
        .I3(\u1/u4/X [14]),
        .I4(\u1/u4/X [18]),
        .I5(\u1/u4/X [13]),
        .O(\u1/out4 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__161
       (.I0(\u1/u4/X [35]),
        .I1(\u1/u4/X [34]),
        .I2(\u1/u4/X [33]),
        .I3(\u1/u4/X [32]),
        .I4(\u1/u4/X [36]),
        .I5(\u1/u4/X [31]),
        .O(\u1/out4 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__162
       (.I0(\u1/u4/X [11]),
        .I1(\u1/u4/X [10]),
        .I2(\u1/u4/X [9]),
        .I3(\u1/u4/X [8]),
        .I4(\u1/u4/X [12]),
        .I5(\u1/u4/X [7]),
        .O(\u1/out4 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__163
       (.I0(\u1/u4/X [47]),
        .I1(\u1/u4/X [46]),
        .I2(\u1/u4/X [45]),
        .I3(\u1/u4/X [44]),
        .I4(\u1/u4/X [48]),
        .I5(\u1/u4/X [43]),
        .O(\u1/out4 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__164
       (.I0(\u1/u4/X [23]),
        .I1(\u1/u4/X [22]),
        .I2(\u1/u4/X [21]),
        .I3(\u1/u4/X [20]),
        .I4(\u1/u4/X [24]),
        .I5(\u1/u4/X [19]),
        .O(\u1/out4 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__165
       (.I0(\u1/u4/X [29]),
        .I1(\u1/u4/X [28]),
        .I2(\u1/u4/X [27]),
        .I3(\u1/u4/X [26]),
        .I4(\u1/u4/X [30]),
        .I5(\u1/u4/X [25]),
        .O(\u1/out4 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__166
       (.I0(\u1/u4/X [5]),
        .I1(\u1/u4/X [4]),
        .I2(\u1/u4/X [3]),
        .I3(\u1/u4/X [2]),
        .I4(\u1/u4/X [6]),
        .I5(\u1/u4/X [1]),
        .O(\u1/out4 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__167
       (.I0(\u1/u5/X [41]),
        .I1(\u1/u5/X [40]),
        .I2(\u1/u5/X [39]),
        .I3(\u1/u5/X [38]),
        .I4(\u1/u5/X [42]),
        .I5(\u1/u5/X [37]),
        .O(\u1/out5 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__168
       (.I0(\u1/u5/X [17]),
        .I1(\u1/u5/X [16]),
        .I2(\u1/u5/X [15]),
        .I3(\u1/u5/X [14]),
        .I4(\u1/u5/X [18]),
        .I5(\u1/u5/X [13]),
        .O(\u1/out5 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__169
       (.I0(\u1/u5/X [35]),
        .I1(\u1/u5/X [34]),
        .I2(\u1/u5/X [33]),
        .I3(\u1/u5/X [32]),
        .I4(\u1/u5/X [36]),
        .I5(\u1/u5/X [31]),
        .O(\u1/out5 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__17
       (.I0(\u0/u2/X [35]),
        .I1(\u0/u2/X [34]),
        .I2(\u0/u2/X [33]),
        .I3(\u0/u2/X [32]),
        .I4(\u0/u2/X [36]),
        .I5(\u0/u2/X [31]),
        .O(\u0/out2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__170
       (.I0(\u1/u5/X [11]),
        .I1(\u1/u5/X [10]),
        .I2(\u1/u5/X [9]),
        .I3(\u1/u5/X [8]),
        .I4(\u1/u5/X [12]),
        .I5(\u1/u5/X [7]),
        .O(\u1/out5 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__171
       (.I0(\u1/u5/X [47]),
        .I1(\u1/u5/X [46]),
        .I2(\u1/u5/X [45]),
        .I3(\u1/u5/X [44]),
        .I4(\u1/u5/X [48]),
        .I5(\u1/u5/X [43]),
        .O(\u1/out5 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__172
       (.I0(\u1/u5/X [23]),
        .I1(\u1/u5/X [22]),
        .I2(\u1/u5/X [21]),
        .I3(\u1/u5/X [20]),
        .I4(\u1/u5/X [24]),
        .I5(\u1/u5/X [19]),
        .O(\u1/out5 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__173
       (.I0(\u1/u5/X [29]),
        .I1(\u1/u5/X [28]),
        .I2(\u1/u5/X [27]),
        .I3(\u1/u5/X [26]),
        .I4(\u1/u5/X [30]),
        .I5(\u1/u5/X [25]),
        .O(\u1/out5 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__174
       (.I0(\u1/u5/X [5]),
        .I1(\u1/u5/X [4]),
        .I2(\u1/u5/X [3]),
        .I3(\u1/u5/X [2]),
        .I4(\u1/u5/X [6]),
        .I5(\u1/u5/X [1]),
        .O(\u1/out5 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__175
       (.I0(\u1/u6/X [41]),
        .I1(\u1/u6/X [40]),
        .I2(\u1/u6/X [39]),
        .I3(\u1/u6/X [38]),
        .I4(\u1/u6/X [42]),
        .I5(\u1/u6/X [37]),
        .O(\u1/out6 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__176
       (.I0(\u1/u6/X [17]),
        .I1(\u1/u6/X [16]),
        .I2(\u1/u6/X [15]),
        .I3(\u1/u6/X [14]),
        .I4(\u1/u6/X [18]),
        .I5(\u1/u6/X [13]),
        .O(\u1/out6 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__177
       (.I0(\u1/u6/X [35]),
        .I1(\u1/u6/X [34]),
        .I2(\u1/u6/X [33]),
        .I3(\u1/u6/X [32]),
        .I4(\u1/u6/X [36]),
        .I5(\u1/u6/X [31]),
        .O(\u1/out6 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__178
       (.I0(\u1/u6/X [11]),
        .I1(\u1/u6/X [10]),
        .I2(\u1/u6/X [9]),
        .I3(\u1/u6/X [8]),
        .I4(\u1/u6/X [12]),
        .I5(\u1/u6/X [7]),
        .O(\u1/out6 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__179
       (.I0(\u1/u6/X [47]),
        .I1(\u1/u6/X [46]),
        .I2(\u1/u6/X [45]),
        .I3(\u1/u6/X [44]),
        .I4(\u1/u6/X [48]),
        .I5(\u1/u6/X [43]),
        .O(\u1/out6 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__18
       (.I0(\u0/u2/X [11]),
        .I1(\u0/u2/X [10]),
        .I2(\u0/u2/X [9]),
        .I3(\u0/u2/X [8]),
        .I4(\u0/u2/X [12]),
        .I5(\u0/u2/X [7]),
        .O(\u0/out2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__180
       (.I0(\u1/u6/X [23]),
        .I1(\u1/u6/X [22]),
        .I2(\u1/u6/X [21]),
        .I3(\u1/u6/X [20]),
        .I4(\u1/u6/X [24]),
        .I5(\u1/u6/X [19]),
        .O(\u1/out6 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__181
       (.I0(\u1/u6/X [29]),
        .I1(\u1/u6/X [28]),
        .I2(\u1/u6/X [27]),
        .I3(\u1/u6/X [26]),
        .I4(\u1/u6/X [30]),
        .I5(\u1/u6/X [25]),
        .O(\u1/out6 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__182
       (.I0(\u1/u6/X [5]),
        .I1(\u1/u6/X [4]),
        .I2(\u1/u6/X [3]),
        .I3(\u1/u6/X [2]),
        .I4(\u1/u6/X [6]),
        .I5(\u1/u6/X [1]),
        .O(\u1/out6 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__183
       (.I0(\u1/u7/X [41]),
        .I1(\u1/u7/X [40]),
        .I2(\u1/u7/X [39]),
        .I3(\u1/u7/X [38]),
        .I4(\u1/u7/X [42]),
        .I5(\u1/u7/X [37]),
        .O(\u1/out7 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__184
       (.I0(\u1/u7/X [17]),
        .I1(\u1/u7/X [16]),
        .I2(\u1/u7/X [15]),
        .I3(\u1/u7/X [14]),
        .I4(\u1/u7/X [18]),
        .I5(\u1/u7/X [13]),
        .O(\u1/out7 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__185
       (.I0(\u1/u7/X [35]),
        .I1(\u1/u7/X [34]),
        .I2(\u1/u7/X [33]),
        .I3(\u1/u7/X [32]),
        .I4(\u1/u7/X [36]),
        .I5(\u1/u7/X [31]),
        .O(\u1/out7 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__186
       (.I0(\u1/u7/X [11]),
        .I1(\u1/u7/X [10]),
        .I2(\u1/u7/X [9]),
        .I3(\u1/u7/X [8]),
        .I4(\u1/u7/X [12]),
        .I5(\u1/u7/X [7]),
        .O(\u1/out7 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__187
       (.I0(\u1/u7/X [47]),
        .I1(\u1/u7/X [46]),
        .I2(\u1/u7/X [45]),
        .I3(\u1/u7/X [44]),
        .I4(\u1/u7/X [48]),
        .I5(\u1/u7/X [43]),
        .O(\u1/out7 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__188
       (.I0(\u1/u7/X [23]),
        .I1(\u1/u7/X [22]),
        .I2(\u1/u7/X [21]),
        .I3(\u1/u7/X [20]),
        .I4(\u1/u7/X [24]),
        .I5(\u1/u7/X [19]),
        .O(\u1/out7 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__189
       (.I0(\u1/u7/X [29]),
        .I1(\u1/u7/X [28]),
        .I2(\u1/u7/X [27]),
        .I3(\u1/u7/X [26]),
        .I4(\u1/u7/X [30]),
        .I5(\u1/u7/X [25]),
        .O(\u1/out7 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__19
       (.I0(\u0/u2/X [47]),
        .I1(\u0/u2/X [46]),
        .I2(\u0/u2/X [45]),
        .I3(\u0/u2/X [44]),
        .I4(\u0/u2/X [48]),
        .I5(\u0/u2/X [43]),
        .O(\u0/out2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__190
       (.I0(\u1/u7/X [5]),
        .I1(\u1/u7/X [4]),
        .I2(\u1/u7/X [3]),
        .I3(\u1/u7/X [2]),
        .I4(\u1/u7/X [6]),
        .I5(\u1/u7/X [1]),
        .O(\u1/out7 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__191
       (.I0(\u1/u8/X [41]),
        .I1(\u1/u8/X [40]),
        .I2(\u1/u8/X [39]),
        .I3(\u1/u8/X [38]),
        .I4(\u1/u8/X [42]),
        .I5(\u1/u8/X [37]),
        .O(\u1/out8 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__192
       (.I0(\u1/u8/X [17]),
        .I1(\u1/u8/X [16]),
        .I2(\u1/u8/X [15]),
        .I3(\u1/u8/X [14]),
        .I4(\u1/u8/X [18]),
        .I5(\u1/u8/X [13]),
        .O(\u1/out8 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__193
       (.I0(\u1/u8/X [35]),
        .I1(\u1/u8/X [34]),
        .I2(\u1/u8/X [33]),
        .I3(\u1/u8/X [32]),
        .I4(\u1/u8/X [36]),
        .I5(\u1/u8/X [31]),
        .O(\u1/out8 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__194
       (.I0(\u1/u8/X [11]),
        .I1(\u1/u8/X [10]),
        .I2(\u1/u8/X [9]),
        .I3(\u1/u8/X [8]),
        .I4(\u1/u8/X [12]),
        .I5(\u1/u8/X [7]),
        .O(\u1/out8 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__195
       (.I0(\u1/u8/X [47]),
        .I1(\u1/u8/X [46]),
        .I2(\u1/u8/X [45]),
        .I3(\u1/u8/X [44]),
        .I4(\u1/u8/X [48]),
        .I5(\u1/u8/X [43]),
        .O(\u1/out8 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__196
       (.I0(\u1/u8/X [23]),
        .I1(\u1/u8/X [22]),
        .I2(\u1/u8/X [21]),
        .I3(\u1/u8/X [20]),
        .I4(\u1/u8/X [24]),
        .I5(\u1/u8/X [19]),
        .O(\u1/out8 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__197
       (.I0(\u1/u8/X [29]),
        .I1(\u1/u8/X [28]),
        .I2(\u1/u8/X [27]),
        .I3(\u1/u8/X [26]),
        .I4(\u1/u8/X [30]),
        .I5(\u1/u8/X [25]),
        .O(\u1/out8 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__198
       (.I0(\u1/u8/X [5]),
        .I1(\u1/u8/X [4]),
        .I2(\u1/u8/X [3]),
        .I3(\u1/u8/X [2]),
        .I4(\u1/u8/X [6]),
        .I5(\u1/u8/X [1]),
        .O(\u1/out8 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__199
       (.I0(\u1/u9/X [41]),
        .I1(\u1/u9/X [40]),
        .I2(\u1/u9/X [39]),
        .I3(\u1/u9/X [38]),
        .I4(\u1/u9/X [42]),
        .I5(\u1/u9/X [37]),
        .O(\u1/out9 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__2
       (.I0(\u0/u0/X [11]),
        .I1(\u0/u0/X [10]),
        .I2(\u0/u0/X [9]),
        .I3(\u0/u0/X [8]),
        .I4(\u0/u0/X [12]),
        .I5(\u0/u0/X [7]),
        .O(\u0/out0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__20
       (.I0(\u0/u2/X [23]),
        .I1(\u0/u2/X [22]),
        .I2(\u0/u2/X [21]),
        .I3(\u0/u2/X [20]),
        .I4(\u0/u2/X [24]),
        .I5(\u0/u2/X [19]),
        .O(\u0/out2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__200
       (.I0(\u1/u9/X [17]),
        .I1(\u1/u9/X [16]),
        .I2(\u1/u9/X [15]),
        .I3(\u1/u9/X [14]),
        .I4(\u1/u9/X [18]),
        .I5(\u1/u9/X [13]),
        .O(\u1/out9 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__201
       (.I0(\u1/u9/X [35]),
        .I1(\u1/u9/X [34]),
        .I2(\u1/u9/X [33]),
        .I3(\u1/u9/X [32]),
        .I4(\u1/u9/X [36]),
        .I5(\u1/u9/X [31]),
        .O(\u1/out9 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__202
       (.I0(\u1/u9/X [11]),
        .I1(\u1/u9/X [10]),
        .I2(\u1/u9/X [9]),
        .I3(\u1/u9/X [8]),
        .I4(\u1/u9/X [12]),
        .I5(\u1/u9/X [7]),
        .O(\u1/out9 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__203
       (.I0(\u1/u9/X [47]),
        .I1(\u1/u9/X [46]),
        .I2(\u1/u9/X [45]),
        .I3(\u1/u9/X [44]),
        .I4(\u1/u9/X [48]),
        .I5(\u1/u9/X [43]),
        .O(\u1/out9 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__204
       (.I0(\u1/u9/X [23]),
        .I1(\u1/u9/X [22]),
        .I2(\u1/u9/X [21]),
        .I3(\u1/u9/X [20]),
        .I4(\u1/u9/X [24]),
        .I5(\u1/u9/X [19]),
        .O(\u1/out9 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__205
       (.I0(\u1/u9/X [29]),
        .I1(\u1/u9/X [28]),
        .I2(\u1/u9/X [27]),
        .I3(\u1/u9/X [26]),
        .I4(\u1/u9/X [30]),
        .I5(\u1/u9/X [25]),
        .O(\u1/out9 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__206
       (.I0(\u1/u9/X [5]),
        .I1(\u1/u9/X [4]),
        .I2(\u1/u9/X [3]),
        .I3(\u1/u9/X [2]),
        .I4(\u1/u9/X [6]),
        .I5(\u1/u9/X [1]),
        .O(\u1/out9 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__207
       (.I0(\u1/u10/X [41]),
        .I1(\u1/u10/X [40]),
        .I2(\u1/u10/X [39]),
        .I3(\u1/u10/X [38]),
        .I4(\u1/u10/X [42]),
        .I5(\u1/u10/X [37]),
        .O(\u1/out10 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__208
       (.I0(\u1/u10/X [17]),
        .I1(\u1/u10/X [16]),
        .I2(\u1/u10/X [15]),
        .I3(\u1/u10/X [14]),
        .I4(\u1/u10/X [18]),
        .I5(\u1/u10/X [13]),
        .O(\u1/out10 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__209
       (.I0(\u1/u10/X [35]),
        .I1(\u1/u10/X [34]),
        .I2(\u1/u10/X [33]),
        .I3(\u1/u10/X [32]),
        .I4(\u1/u10/X [36]),
        .I5(\u1/u10/X [31]),
        .O(\u1/out10 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__21
       (.I0(\u0/u2/X [29]),
        .I1(\u0/u2/X [28]),
        .I2(\u0/u2/X [27]),
        .I3(\u0/u2/X [26]),
        .I4(\u0/u2/X [30]),
        .I5(\u0/u2/X [25]),
        .O(\u0/out2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__210
       (.I0(\u1/u10/X [11]),
        .I1(\u1/u10/X [10]),
        .I2(\u1/u10/X [9]),
        .I3(\u1/u10/X [8]),
        .I4(\u1/u10/X [12]),
        .I5(\u1/u10/X [7]),
        .O(\u1/out10 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__211
       (.I0(\u1/u10/X [47]),
        .I1(\u1/u10/X [46]),
        .I2(\u1/u10/X [45]),
        .I3(\u1/u10/X [44]),
        .I4(\u1/u10/X [48]),
        .I5(\u1/u10/X [43]),
        .O(\u1/out10 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__212
       (.I0(\u1/u10/X [23]),
        .I1(\u1/u10/X [22]),
        .I2(\u1/u10/X [21]),
        .I3(\u1/u10/X [20]),
        .I4(\u1/u10/X [24]),
        .I5(\u1/u10/X [19]),
        .O(\u1/out10 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__213
       (.I0(\u1/u10/X [29]),
        .I1(\u1/u10/X [28]),
        .I2(\u1/u10/X [27]),
        .I3(\u1/u10/X [26]),
        .I4(\u1/u10/X [30]),
        .I5(\u1/u10/X [25]),
        .O(\u1/out10 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__214
       (.I0(\u1/u10/X [5]),
        .I1(\u1/u10/X [4]),
        .I2(\u1/u10/X [3]),
        .I3(\u1/u10/X [2]),
        .I4(\u1/u10/X [6]),
        .I5(\u1/u10/X [1]),
        .O(\u1/out10 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__215
       (.I0(\u1/u11/X [41]),
        .I1(\u1/u11/X [40]),
        .I2(\u1/u11/X [39]),
        .I3(\u1/u11/X [38]),
        .I4(\u1/u11/X [42]),
        .I5(\u1/u11/X [37]),
        .O(\u1/out11 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__216
       (.I0(\u1/u11/X [17]),
        .I1(\u1/u11/X [16]),
        .I2(\u1/u11/X [15]),
        .I3(\u1/u11/X [14]),
        .I4(\u1/u11/X [18]),
        .I5(\u1/u11/X [13]),
        .O(\u1/out11 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__217
       (.I0(\u1/u11/X [35]),
        .I1(\u1/u11/X [34]),
        .I2(\u1/u11/X [33]),
        .I3(\u1/u11/X [32]),
        .I4(\u1/u11/X [36]),
        .I5(\u1/u11/X [31]),
        .O(\u1/out11 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__218
       (.I0(\u1/u11/X [11]),
        .I1(\u1/u11/X [10]),
        .I2(\u1/u11/X [9]),
        .I3(\u1/u11/X [8]),
        .I4(\u1/u11/X [12]),
        .I5(\u1/u11/X [7]),
        .O(\u1/out11 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__219
       (.I0(\u1/u11/X [47]),
        .I1(\u1/u11/X [46]),
        .I2(\u1/u11/X [45]),
        .I3(\u1/u11/X [44]),
        .I4(\u1/u11/X [48]),
        .I5(\u1/u11/X [43]),
        .O(\u1/out11 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__22
       (.I0(\u0/u2/X [5]),
        .I1(\u0/u2/X [4]),
        .I2(\u0/u2/X [3]),
        .I3(\u0/u2/X [2]),
        .I4(\u0/u2/X [6]),
        .I5(\u0/u2/X [1]),
        .O(\u0/out2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__220
       (.I0(\u1/u11/X [23]),
        .I1(\u1/u11/X [22]),
        .I2(\u1/u11/X [21]),
        .I3(\u1/u11/X [20]),
        .I4(\u1/u11/X [24]),
        .I5(\u1/u11/X [19]),
        .O(\u1/out11 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__221
       (.I0(\u1/u11/X [29]),
        .I1(\u1/u11/X [28]),
        .I2(\u1/u11/X [27]),
        .I3(\u1/u11/X [26]),
        .I4(\u1/u11/X [30]),
        .I5(\u1/u11/X [25]),
        .O(\u1/out11 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__222
       (.I0(\u1/u11/X [5]),
        .I1(\u1/u11/X [4]),
        .I2(\u1/u11/X [3]),
        .I3(\u1/u11/X [2]),
        .I4(\u1/u11/X [6]),
        .I5(\u1/u11/X [1]),
        .O(\u1/out11 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__223
       (.I0(\u1/u12/X [41]),
        .I1(\u1/u12/X [40]),
        .I2(\u1/u12/X [39]),
        .I3(\u1/u12/X [38]),
        .I4(\u1/u12/X [42]),
        .I5(\u1/u12/X [37]),
        .O(\u1/out12 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__224
       (.I0(\u1/u12/X [17]),
        .I1(\u1/u12/X [16]),
        .I2(\u1/u12/X [15]),
        .I3(\u1/u12/X [14]),
        .I4(\u1/u12/X [18]),
        .I5(\u1/u12/X [13]),
        .O(\u1/out12 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__225
       (.I0(\u1/u12/X [35]),
        .I1(\u1/u12/X [34]),
        .I2(\u1/u12/X [33]),
        .I3(\u1/u12/X [32]),
        .I4(\u1/u12/X [36]),
        .I5(\u1/u12/X [31]),
        .O(\u1/out12 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__226
       (.I0(\u1/u12/X [11]),
        .I1(\u1/u12/X [10]),
        .I2(\u1/u12/X [9]),
        .I3(\u1/u12/X [8]),
        .I4(\u1/u12/X [12]),
        .I5(\u1/u12/X [7]),
        .O(\u1/out12 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__227
       (.I0(\u1/u12/X [47]),
        .I1(\u1/u12/X [46]),
        .I2(\u1/u12/X [45]),
        .I3(\u1/u12/X [44]),
        .I4(\u1/u12/X [48]),
        .I5(\u1/u12/X [43]),
        .O(\u1/out12 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__228
       (.I0(\u1/u12/X [23]),
        .I1(\u1/u12/X [22]),
        .I2(\u1/u12/X [21]),
        .I3(\u1/u12/X [20]),
        .I4(\u1/u12/X [24]),
        .I5(\u1/u12/X [19]),
        .O(\u1/out12 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__229
       (.I0(\u1/u12/X [29]),
        .I1(\u1/u12/X [28]),
        .I2(\u1/u12/X [27]),
        .I3(\u1/u12/X [26]),
        .I4(\u1/u12/X [30]),
        .I5(\u1/u12/X [25]),
        .O(\u1/out12 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__23
       (.I0(\u0/u3/X [41]),
        .I1(\u0/u3/X [40]),
        .I2(\u0/u3/X [39]),
        .I3(\u0/u3/X [38]),
        .I4(\u0/u3/X [42]),
        .I5(\u0/u3/X [37]),
        .O(\u0/out3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__230
       (.I0(\u1/u12/X [5]),
        .I1(\u1/u12/X [4]),
        .I2(\u1/u12/X [3]),
        .I3(\u1/u12/X [2]),
        .I4(\u1/u12/X [6]),
        .I5(\u1/u12/X [1]),
        .O(\u1/out12 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__231
       (.I0(\u1/u13/X [41]),
        .I1(\u1/u13/X [40]),
        .I2(\u1/u13/X [39]),
        .I3(\u1/u13/X [38]),
        .I4(\u1/u13/X [42]),
        .I5(\u1/u13/X [37]),
        .O(\u1/out13 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__232
       (.I0(\u1/u13/X [17]),
        .I1(\u1/u13/X [16]),
        .I2(\u1/u13/X [15]),
        .I3(\u1/u13/X [14]),
        .I4(\u1/u13/X [18]),
        .I5(\u1/u13/X [13]),
        .O(\u1/out13 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__233
       (.I0(\u1/u13/X [35]),
        .I1(\u1/u13/X [34]),
        .I2(\u1/u13/X [33]),
        .I3(\u1/u13/X [32]),
        .I4(\u1/u13/X [36]),
        .I5(\u1/u13/X [31]),
        .O(\u1/out13 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__234
       (.I0(\u1/u13/X [11]),
        .I1(\u1/u13/X [10]),
        .I2(\u1/u13/X [9]),
        .I3(\u1/u13/X [8]),
        .I4(\u1/u13/X [12]),
        .I5(\u1/u13/X [7]),
        .O(\u1/out13 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__235
       (.I0(\u1/u13/X [47]),
        .I1(\u1/u13/X [46]),
        .I2(\u1/u13/X [45]),
        .I3(\u1/u13/X [44]),
        .I4(\u1/u13/X [48]),
        .I5(\u1/u13/X [43]),
        .O(\u1/out13 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__236
       (.I0(\u1/u13/X [23]),
        .I1(\u1/u13/X [22]),
        .I2(\u1/u13/X [21]),
        .I3(\u1/u13/X [20]),
        .I4(\u1/u13/X [24]),
        .I5(\u1/u13/X [19]),
        .O(\u1/out13 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__237
       (.I0(\u1/u13/X [29]),
        .I1(\u1/u13/X [28]),
        .I2(\u1/u13/X [27]),
        .I3(\u1/u13/X [26]),
        .I4(\u1/u13/X [30]),
        .I5(\u1/u13/X [25]),
        .O(\u1/out13 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__238
       (.I0(\u1/u13/X [5]),
        .I1(\u1/u13/X [4]),
        .I2(\u1/u13/X [3]),
        .I3(\u1/u13/X [2]),
        .I4(\u1/u13/X [6]),
        .I5(\u1/u13/X [1]),
        .O(\u1/out13 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__239
       (.I0(\u1/u14/X [41]),
        .I1(\u1/u14/X [40]),
        .I2(\u1/u14/X [39]),
        .I3(\u1/u14/X [38]),
        .I4(\u1/u14/X [42]),
        .I5(\u1/u14/X [37]),
        .O(\u1/out14 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__24
       (.I0(\u0/u3/X [17]),
        .I1(\u0/u3/X [16]),
        .I2(\u0/u3/X [15]),
        .I3(\u0/u3/X [14]),
        .I4(\u0/u3/X [18]),
        .I5(\u0/u3/X [13]),
        .O(\u0/out3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__240
       (.I0(\u1/u14/X [17]),
        .I1(\u1/u14/X [16]),
        .I2(\u1/u14/X [15]),
        .I3(\u1/u14/X [14]),
        .I4(\u1/u14/X [18]),
        .I5(\u1/u14/X [13]),
        .O(\u1/out14 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__241
       (.I0(\u1/u14/X [35]),
        .I1(\u1/u14/X [34]),
        .I2(\u1/u14/X [33]),
        .I3(\u1/u14/X [32]),
        .I4(\u1/u14/X [36]),
        .I5(\u1/u14/X [31]),
        .O(\u1/out14 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__242
       (.I0(\u1/u14/X [11]),
        .I1(\u1/u14/X [10]),
        .I2(\u1/u14/X [9]),
        .I3(\u1/u14/X [8]),
        .I4(\u1/u14/X [12]),
        .I5(\u1/u14/X [7]),
        .O(\u1/out14 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__243
       (.I0(\u1/u14/X [47]),
        .I1(\u1/u14/X [46]),
        .I2(\u1/u14/X [45]),
        .I3(\u1/u14/X [44]),
        .I4(\u1/u14/X [48]),
        .I5(\u1/u14/X [43]),
        .O(\u1/out14 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__244
       (.I0(\u1/u14/X [23]),
        .I1(\u1/u14/X [22]),
        .I2(\u1/u14/X [21]),
        .I3(\u1/u14/X [20]),
        .I4(\u1/u14/X [24]),
        .I5(\u1/u14/X [19]),
        .O(\u1/out14 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__245
       (.I0(\u1/u14/X [29]),
        .I1(\u1/u14/X [28]),
        .I2(\u1/u14/X [27]),
        .I3(\u1/u14/X [26]),
        .I4(\u1/u14/X [30]),
        .I5(\u1/u14/X [25]),
        .O(\u1/out14 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__246
       (.I0(\u1/u14/X [5]),
        .I1(\u1/u14/X [4]),
        .I2(\u1/u14/X [3]),
        .I3(\u1/u14/X [2]),
        .I4(\u1/u14/X [6]),
        .I5(\u1/u14/X [1]),
        .O(\u1/out14 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__247
       (.I0(\u1/u15/X [41]),
        .I1(\u1/u15/X [40]),
        .I2(\u1/u15/X [39]),
        .I3(\u1/u15/X [38]),
        .I4(\u1/u15/X [42]),
        .I5(\u1/u15/X [37]),
        .O(\u1/out15 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__248
       (.I0(\u1/u15/X [17]),
        .I1(\u1/u15/X [16]),
        .I2(\u1/u15/X [15]),
        .I3(\u1/u15/X [14]),
        .I4(\u1/u15/X [18]),
        .I5(\u1/u15/X [13]),
        .O(\u1/out15 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__249
       (.I0(\u1/u15/X [35]),
        .I1(\u1/u15/X [34]),
        .I2(\u1/u15/X [33]),
        .I3(\u1/u15/X [32]),
        .I4(\u1/u15/X [36]),
        .I5(\u1/u15/X [31]),
        .O(\u1/out15 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__25
       (.I0(\u0/u3/X [35]),
        .I1(\u0/u3/X [34]),
        .I2(\u0/u3/X [33]),
        .I3(\u0/u3/X [32]),
        .I4(\u0/u3/X [36]),
        .I5(\u0/u3/X [31]),
        .O(\u0/out3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__250
       (.I0(\u1/u15/X [11]),
        .I1(\u1/u15/X [10]),
        .I2(\u1/u15/X [9]),
        .I3(\u1/u15/X [8]),
        .I4(\u1/u15/X [12]),
        .I5(\u1/u15/X [7]),
        .O(\u1/out15 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__251
       (.I0(\u1/u15/X [47]),
        .I1(\u1/u15/X [46]),
        .I2(\u1/u15/X [45]),
        .I3(\u1/u15/X [44]),
        .I4(\u1/u15/X [48]),
        .I5(\u1/u15/X [43]),
        .O(\u1/out15 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__252
       (.I0(\u1/u15/X [23]),
        .I1(\u1/u15/X [22]),
        .I2(\u1/u15/X [21]),
        .I3(\u1/u15/X [20]),
        .I4(\u1/u15/X [24]),
        .I5(\u1/u15/X [19]),
        .O(\u1/out15 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__253
       (.I0(\u1/u15/X [29]),
        .I1(\u1/u15/X [28]),
        .I2(\u1/u15/X [27]),
        .I3(\u1/u15/X [26]),
        .I4(\u1/u15/X [30]),
        .I5(\u1/u15/X [25]),
        .O(\u1/out15 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__254
       (.I0(\u1/u15/X [5]),
        .I1(\u1/u15/X [4]),
        .I2(\u1/u15/X [3]),
        .I3(\u1/u15/X [2]),
        .I4(\u1/u15/X [6]),
        .I5(\u1/u15/X [1]),
        .O(\u1/out15 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__255
       (.I0(\u2/u0/X [41]),
        .I1(\u2/u0/X [40]),
        .I2(\u2/u0/X [39]),
        .I3(\u2/u0/X [38]),
        .I4(\u2/u0/X [42]),
        .I5(\u2/u0/X [37]),
        .O(\u2/out0 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__256
       (.I0(\u2/u0/X [17]),
        .I1(\u2/u0/X [16]),
        .I2(\u2/u0/X [15]),
        .I3(\u2/u0/X [14]),
        .I4(\u2/u0/X [18]),
        .I5(\u2/u0/X [13]),
        .O(\u2/out0 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__257
       (.I0(\u2/u0/X [35]),
        .I1(\u2/u0/X [34]),
        .I2(\u2/u0/X [33]),
        .I3(\u2/u0/X [32]),
        .I4(\u2/u0/X [36]),
        .I5(\u2/u0/X [31]),
        .O(\u2/out0 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__258
       (.I0(\u2/u0/X [11]),
        .I1(\u2/u0/X [10]),
        .I2(\u2/u0/X [9]),
        .I3(\u2/u0/X [8]),
        .I4(\u2/u0/X [12]),
        .I5(\u2/u0/X [7]),
        .O(\u2/out0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__259
       (.I0(\u2/u0/X [47]),
        .I1(\u2/u0/X [46]),
        .I2(\u2/u0/X [45]),
        .I3(\u2/u0/X [44]),
        .I4(\u2/u0/X [48]),
        .I5(\u2/u0/X [43]),
        .O(\u2/out0 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__26
       (.I0(\u0/u3/X [11]),
        .I1(\u0/u3/X [10]),
        .I2(\u0/u3/X [9]),
        .I3(\u0/u3/X [8]),
        .I4(\u0/u3/X [12]),
        .I5(\u0/u3/X [7]),
        .O(\u0/out3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__260
       (.I0(\u2/u0/X [23]),
        .I1(\u2/u0/X [22]),
        .I2(\u2/u0/X [21]),
        .I3(\u2/u0/X [20]),
        .I4(\u2/u0/X [24]),
        .I5(\u2/u0/X [19]),
        .O(\u2/out0 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__261
       (.I0(\u2/u0/X [29]),
        .I1(\u2/u0/X [28]),
        .I2(\u2/u0/X [27]),
        .I3(\u2/u0/X [26]),
        .I4(\u2/u0/X [30]),
        .I5(\u2/u0/X [25]),
        .O(\u2/out0 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__262
       (.I0(\u2/u0/X [5]),
        .I1(\u2/u0/X [4]),
        .I2(\u2/u0/X [3]),
        .I3(\u2/u0/X [2]),
        .I4(\u2/u0/X [6]),
        .I5(\u2/u0/X [1]),
        .O(\u2/out0 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__263
       (.I0(\u2/u1/X [41]),
        .I1(\u2/u1/X [40]),
        .I2(\u2/u1/X [39]),
        .I3(\u2/u1/X [38]),
        .I4(\u2/u1/X [42]),
        .I5(\u2/u1/X [37]),
        .O(\u2/out1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__264
       (.I0(\u2/u1/X [17]),
        .I1(\u2/u1/X [16]),
        .I2(\u2/u1/X [15]),
        .I3(\u2/u1/X [14]),
        .I4(\u2/u1/X [18]),
        .I5(\u2/u1/X [13]),
        .O(\u2/out1 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__265
       (.I0(\u2/u1/X [35]),
        .I1(\u2/u1/X [34]),
        .I2(\u2/u1/X [33]),
        .I3(\u2/u1/X [32]),
        .I4(\u2/u1/X [36]),
        .I5(\u2/u1/X [31]),
        .O(\u2/out1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__266
       (.I0(\u2/u1/X [11]),
        .I1(\u2/u1/X [10]),
        .I2(\u2/u1/X [9]),
        .I3(\u2/u1/X [8]),
        .I4(\u2/u1/X [12]),
        .I5(\u2/u1/X [7]),
        .O(\u2/out1 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__267
       (.I0(\u2/u1/X [47]),
        .I1(\u2/u1/X [46]),
        .I2(\u2/u1/X [45]),
        .I3(\u2/u1/X [44]),
        .I4(\u2/u1/X [48]),
        .I5(\u2/u1/X [43]),
        .O(\u2/out1 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__268
       (.I0(\u2/u1/X [23]),
        .I1(\u2/u1/X [22]),
        .I2(\u2/u1/X [21]),
        .I3(\u2/u1/X [20]),
        .I4(\u2/u1/X [24]),
        .I5(\u2/u1/X [19]),
        .O(\u2/out1 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__269
       (.I0(\u2/u1/X [29]),
        .I1(\u2/u1/X [28]),
        .I2(\u2/u1/X [27]),
        .I3(\u2/u1/X [26]),
        .I4(\u2/u1/X [30]),
        .I5(\u2/u1/X [25]),
        .O(\u2/out1 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__27
       (.I0(\u0/u3/X [47]),
        .I1(\u0/u3/X [46]),
        .I2(\u0/u3/X [45]),
        .I3(\u0/u3/X [44]),
        .I4(\u0/u3/X [48]),
        .I5(\u0/u3/X [43]),
        .O(\u0/out3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__270
       (.I0(\u2/u1/X [5]),
        .I1(\u2/u1/X [4]),
        .I2(\u2/u1/X [3]),
        .I3(\u2/u1/X [2]),
        .I4(\u2/u1/X [6]),
        .I5(\u2/u1/X [1]),
        .O(\u2/out1 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__271
       (.I0(\u2/u2/X [41]),
        .I1(\u2/u2/X [40]),
        .I2(\u2/u2/X [39]),
        .I3(\u2/u2/X [38]),
        .I4(\u2/u2/X [42]),
        .I5(\u2/u2/X [37]),
        .O(\u2/out2 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__272
       (.I0(\u2/u2/X [17]),
        .I1(\u2/u2/X [16]),
        .I2(\u2/u2/X [15]),
        .I3(\u2/u2/X [14]),
        .I4(\u2/u2/X [18]),
        .I5(\u2/u2/X [13]),
        .O(\u2/out2 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__273
       (.I0(\u2/u2/X [35]),
        .I1(\u2/u2/X [34]),
        .I2(\u2/u2/X [33]),
        .I3(\u2/u2/X [32]),
        .I4(\u2/u2/X [36]),
        .I5(\u2/u2/X [31]),
        .O(\u2/out2 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__274
       (.I0(\u2/u2/X [11]),
        .I1(\u2/u2/X [10]),
        .I2(\u2/u2/X [9]),
        .I3(\u2/u2/X [8]),
        .I4(\u2/u2/X [12]),
        .I5(\u2/u2/X [7]),
        .O(\u2/out2 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__275
       (.I0(\u2/u2/X [47]),
        .I1(\u2/u2/X [46]),
        .I2(\u2/u2/X [45]),
        .I3(\u2/u2/X [44]),
        .I4(\u2/u2/X [48]),
        .I5(\u2/u2/X [43]),
        .O(\u2/out2 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__276
       (.I0(\u2/u2/X [23]),
        .I1(\u2/u2/X [22]),
        .I2(\u2/u2/X [21]),
        .I3(\u2/u2/X [20]),
        .I4(\u2/u2/X [24]),
        .I5(\u2/u2/X [19]),
        .O(\u2/out2 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__277
       (.I0(\u2/u2/X [29]),
        .I1(\u2/u2/X [28]),
        .I2(\u2/u2/X [27]),
        .I3(\u2/u2/X [26]),
        .I4(\u2/u2/X [30]),
        .I5(\u2/u2/X [25]),
        .O(\u2/out2 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__278
       (.I0(\u2/u2/X [5]),
        .I1(\u2/u2/X [4]),
        .I2(\u2/u2/X [3]),
        .I3(\u2/u2/X [2]),
        .I4(\u2/u2/X [6]),
        .I5(\u2/u2/X [1]),
        .O(\u2/out2 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__279
       (.I0(\u2/u3/X [41]),
        .I1(\u2/u3/X [40]),
        .I2(\u2/u3/X [39]),
        .I3(\u2/u3/X [38]),
        .I4(\u2/u3/X [42]),
        .I5(\u2/u3/X [37]),
        .O(\u2/out3 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__28
       (.I0(\u0/u3/X [23]),
        .I1(\u0/u3/X [22]),
        .I2(\u0/u3/X [21]),
        .I3(\u0/u3/X [20]),
        .I4(\u0/u3/X [24]),
        .I5(\u0/u3/X [19]),
        .O(\u0/out3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__280
       (.I0(\u2/u3/X [17]),
        .I1(\u2/u3/X [16]),
        .I2(\u2/u3/X [15]),
        .I3(\u2/u3/X [14]),
        .I4(\u2/u3/X [18]),
        .I5(\u2/u3/X [13]),
        .O(\u2/out3 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__281
       (.I0(\u2/u3/X [35]),
        .I1(\u2/u3/X [34]),
        .I2(\u2/u3/X [33]),
        .I3(\u2/u3/X [32]),
        .I4(\u2/u3/X [36]),
        .I5(\u2/u3/X [31]),
        .O(\u2/out3 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__282
       (.I0(\u2/u3/X [11]),
        .I1(\u2/u3/X [10]),
        .I2(\u2/u3/X [9]),
        .I3(\u2/u3/X [8]),
        .I4(\u2/u3/X [12]),
        .I5(\u2/u3/X [7]),
        .O(\u2/out3 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__283
       (.I0(\u2/u3/X [47]),
        .I1(\u2/u3/X [46]),
        .I2(\u2/u3/X [45]),
        .I3(\u2/u3/X [44]),
        .I4(\u2/u3/X [48]),
        .I5(\u2/u3/X [43]),
        .O(\u2/out3 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__284
       (.I0(\u2/u3/X [23]),
        .I1(\u2/u3/X [22]),
        .I2(\u2/u3/X [21]),
        .I3(\u2/u3/X [20]),
        .I4(\u2/u3/X [24]),
        .I5(\u2/u3/X [19]),
        .O(\u2/out3 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__285
       (.I0(\u2/u3/X [29]),
        .I1(\u2/u3/X [28]),
        .I2(\u2/u3/X [27]),
        .I3(\u2/u3/X [26]),
        .I4(\u2/u3/X [30]),
        .I5(\u2/u3/X [25]),
        .O(\u2/out3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__286
       (.I0(\u2/u3/X [5]),
        .I1(\u2/u3/X [4]),
        .I2(\u2/u3/X [3]),
        .I3(\u2/u3/X [2]),
        .I4(\u2/u3/X [6]),
        .I5(\u2/u3/X [1]),
        .O(\u2/out3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__287
       (.I0(\u2/u4/X [41]),
        .I1(\u2/u4/X [40]),
        .I2(\u2/u4/X [39]),
        .I3(\u2/u4/X [38]),
        .I4(\u2/u4/X [42]),
        .I5(\u2/u4/X [37]),
        .O(\u2/out4 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__288
       (.I0(\u2/u4/X [17]),
        .I1(\u2/u4/X [16]),
        .I2(\u2/u4/X [15]),
        .I3(\u2/u4/X [14]),
        .I4(\u2/u4/X [18]),
        .I5(\u2/u4/X [13]),
        .O(\u2/out4 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__289
       (.I0(\u2/u4/X [35]),
        .I1(\u2/u4/X [34]),
        .I2(\u2/u4/X [33]),
        .I3(\u2/u4/X [32]),
        .I4(\u2/u4/X [36]),
        .I5(\u2/u4/X [31]),
        .O(\u2/out4 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__29
       (.I0(\u0/u3/X [29]),
        .I1(\u0/u3/X [28]),
        .I2(\u0/u3/X [27]),
        .I3(\u0/u3/X [26]),
        .I4(\u0/u3/X [30]),
        .I5(\u0/u3/X [25]),
        .O(\u0/out3 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__290
       (.I0(\u2/u4/X [11]),
        .I1(\u2/u4/X [10]),
        .I2(\u2/u4/X [9]),
        .I3(\u2/u4/X [8]),
        .I4(\u2/u4/X [12]),
        .I5(\u2/u4/X [7]),
        .O(\u2/out4 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__291
       (.I0(\u2/u4/X [47]),
        .I1(\u2/u4/X [46]),
        .I2(\u2/u4/X [45]),
        .I3(\u2/u4/X [44]),
        .I4(\u2/u4/X [48]),
        .I5(\u2/u4/X [43]),
        .O(\u2/out4 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__292
       (.I0(\u2/u4/X [23]),
        .I1(\u2/u4/X [22]),
        .I2(\u2/u4/X [21]),
        .I3(\u2/u4/X [20]),
        .I4(\u2/u4/X [24]),
        .I5(\u2/u4/X [19]),
        .O(\u2/out4 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__293
       (.I0(\u2/u4/X [29]),
        .I1(\u2/u4/X [28]),
        .I2(\u2/u4/X [27]),
        .I3(\u2/u4/X [26]),
        .I4(\u2/u4/X [30]),
        .I5(\u2/u4/X [25]),
        .O(\u2/out4 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__294
       (.I0(\u2/u4/X [5]),
        .I1(\u2/u4/X [4]),
        .I2(\u2/u4/X [3]),
        .I3(\u2/u4/X [2]),
        .I4(\u2/u4/X [6]),
        .I5(\u2/u4/X [1]),
        .O(\u2/out4 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__295
       (.I0(\u2/u5/X [41]),
        .I1(\u2/u5/X [40]),
        .I2(\u2/u5/X [39]),
        .I3(\u2/u5/X [38]),
        .I4(\u2/u5/X [42]),
        .I5(\u2/u5/X [37]),
        .O(\u2/out5 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__296
       (.I0(\u2/u5/X [17]),
        .I1(\u2/u5/X [16]),
        .I2(\u2/u5/X [15]),
        .I3(\u2/u5/X [14]),
        .I4(\u2/u5/X [18]),
        .I5(\u2/u5/X [13]),
        .O(\u2/out5 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__297
       (.I0(\u2/u5/X [35]),
        .I1(\u2/u5/X [34]),
        .I2(\u2/u5/X [33]),
        .I3(\u2/u5/X [32]),
        .I4(\u2/u5/X [36]),
        .I5(\u2/u5/X [31]),
        .O(\u2/out5 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__298
       (.I0(\u2/u5/X [11]),
        .I1(\u2/u5/X [10]),
        .I2(\u2/u5/X [9]),
        .I3(\u2/u5/X [8]),
        .I4(\u2/u5/X [12]),
        .I5(\u2/u5/X [7]),
        .O(\u2/out5 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__299
       (.I0(\u2/u5/X [47]),
        .I1(\u2/u5/X [46]),
        .I2(\u2/u5/X [45]),
        .I3(\u2/u5/X [44]),
        .I4(\u2/u5/X [48]),
        .I5(\u2/u5/X [43]),
        .O(\u2/out5 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__3
       (.I0(\u0/u0/X [47]),
        .I1(\u0/u0/X [46]),
        .I2(\u0/u0/X [45]),
        .I3(\u0/u0/X [44]),
        .I4(\u0/u0/X [48]),
        .I5(\u0/u0/X [43]),
        .O(\u0/out0 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__30
       (.I0(\u0/u3/X [5]),
        .I1(\u0/u3/X [4]),
        .I2(\u0/u3/X [3]),
        .I3(\u0/u3/X [2]),
        .I4(\u0/u3/X [6]),
        .I5(\u0/u3/X [1]),
        .O(\u0/out3 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__300
       (.I0(\u2/u5/X [23]),
        .I1(\u2/u5/X [22]),
        .I2(\u2/u5/X [21]),
        .I3(\u2/u5/X [20]),
        .I4(\u2/u5/X [24]),
        .I5(\u2/u5/X [19]),
        .O(\u2/out5 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__301
       (.I0(\u2/u5/X [29]),
        .I1(\u2/u5/X [28]),
        .I2(\u2/u5/X [27]),
        .I3(\u2/u5/X [26]),
        .I4(\u2/u5/X [30]),
        .I5(\u2/u5/X [25]),
        .O(\u2/out5 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__302
       (.I0(\u2/u5/X [5]),
        .I1(\u2/u5/X [4]),
        .I2(\u2/u5/X [3]),
        .I3(\u2/u5/X [2]),
        .I4(\u2/u5/X [6]),
        .I5(\u2/u5/X [1]),
        .O(\u2/out5 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__303
       (.I0(\u2/u6/X [41]),
        .I1(\u2/u6/X [40]),
        .I2(\u2/u6/X [39]),
        .I3(\u2/u6/X [38]),
        .I4(\u2/u6/X [42]),
        .I5(\u2/u6/X [37]),
        .O(\u2/out6 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__304
       (.I0(\u2/u6/X [17]),
        .I1(\u2/u6/X [16]),
        .I2(\u2/u6/X [15]),
        .I3(\u2/u6/X [14]),
        .I4(\u2/u6/X [18]),
        .I5(\u2/u6/X [13]),
        .O(\u2/out6 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__305
       (.I0(\u2/u6/X [35]),
        .I1(\u2/u6/X [34]),
        .I2(\u2/u6/X [33]),
        .I3(\u2/u6/X [32]),
        .I4(\u2/u6/X [36]),
        .I5(\u2/u6/X [31]),
        .O(\u2/out6 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__306
       (.I0(\u2/u6/X [11]),
        .I1(\u2/u6/X [10]),
        .I2(\u2/u6/X [9]),
        .I3(\u2/u6/X [8]),
        .I4(\u2/u6/X [12]),
        .I5(\u2/u6/X [7]),
        .O(\u2/out6 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__307
       (.I0(\u2/u6/X [47]),
        .I1(\u2/u6/X [46]),
        .I2(\u2/u6/X [45]),
        .I3(\u2/u6/X [44]),
        .I4(\u2/u6/X [48]),
        .I5(\u2/u6/X [43]),
        .O(\u2/out6 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__308
       (.I0(\u2/u6/X [23]),
        .I1(\u2/u6/X [22]),
        .I2(\u2/u6/X [21]),
        .I3(\u2/u6/X [20]),
        .I4(\u2/u6/X [24]),
        .I5(\u2/u6/X [19]),
        .O(\u2/out6 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__309
       (.I0(\u2/u6/X [29]),
        .I1(\u2/u6/X [28]),
        .I2(\u2/u6/X [27]),
        .I3(\u2/u6/X [26]),
        .I4(\u2/u6/X [30]),
        .I5(\u2/u6/X [25]),
        .O(\u2/out6 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__31
       (.I0(\u0/u4/X [41]),
        .I1(\u0/u4/X [40]),
        .I2(\u0/u4/X [39]),
        .I3(\u0/u4/X [38]),
        .I4(\u0/u4/X [42]),
        .I5(\u0/u4/X [37]),
        .O(\u0/out4 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__310
       (.I0(\u2/u6/X [5]),
        .I1(\u2/u6/X [4]),
        .I2(\u2/u6/X [3]),
        .I3(\u2/u6/X [2]),
        .I4(\u2/u6/X [6]),
        .I5(\u2/u6/X [1]),
        .O(\u2/out6 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__311
       (.I0(\u2/u7/X [41]),
        .I1(\u2/u7/X [40]),
        .I2(\u2/u7/X [39]),
        .I3(\u2/u7/X [38]),
        .I4(\u2/u7/X [42]),
        .I5(\u2/u7/X [37]),
        .O(\u2/out7 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__312
       (.I0(\u2/u7/X [17]),
        .I1(\u2/u7/X [16]),
        .I2(\u2/u7/X [15]),
        .I3(\u2/u7/X [14]),
        .I4(\u2/u7/X [18]),
        .I5(\u2/u7/X [13]),
        .O(\u2/out7 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__313
       (.I0(\u2/u7/X [35]),
        .I1(\u2/u7/X [34]),
        .I2(\u2/u7/X [33]),
        .I3(\u2/u7/X [32]),
        .I4(\u2/u7/X [36]),
        .I5(\u2/u7/X [31]),
        .O(\u2/out7 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__314
       (.I0(\u2/u7/X [11]),
        .I1(\u2/u7/X [10]),
        .I2(\u2/u7/X [9]),
        .I3(\u2/u7/X [8]),
        .I4(\u2/u7/X [12]),
        .I5(\u2/u7/X [7]),
        .O(\u2/out7 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__315
       (.I0(\u2/u7/X [47]),
        .I1(\u2/u7/X [46]),
        .I2(\u2/u7/X [45]),
        .I3(\u2/u7/X [44]),
        .I4(\u2/u7/X [48]),
        .I5(\u2/u7/X [43]),
        .O(\u2/out7 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__316
       (.I0(\u2/u7/X [23]),
        .I1(\u2/u7/X [22]),
        .I2(\u2/u7/X [21]),
        .I3(\u2/u7/X [20]),
        .I4(\u2/u7/X [24]),
        .I5(\u2/u7/X [19]),
        .O(\u2/out7 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__317
       (.I0(\u2/u7/X [29]),
        .I1(\u2/u7/X [28]),
        .I2(\u2/u7/X [27]),
        .I3(\u2/u7/X [26]),
        .I4(\u2/u7/X [30]),
        .I5(\u2/u7/X [25]),
        .O(\u2/out7 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__318
       (.I0(\u2/u7/X [5]),
        .I1(\u2/u7/X [4]),
        .I2(\u2/u7/X [3]),
        .I3(\u2/u7/X [2]),
        .I4(\u2/u7/X [6]),
        .I5(\u2/u7/X [1]),
        .O(\u2/out7 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__319
       (.I0(\u2/u8/X [41]),
        .I1(\u2/u8/X [40]),
        .I2(\u2/u8/X [39]),
        .I3(\u2/u8/X [38]),
        .I4(\u2/u8/X [42]),
        .I5(\u2/u8/X [37]),
        .O(\u2/out8 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__32
       (.I0(\u0/u4/X [17]),
        .I1(\u0/u4/X [16]),
        .I2(\u0/u4/X [15]),
        .I3(\u0/u4/X [14]),
        .I4(\u0/u4/X [18]),
        .I5(\u0/u4/X [13]),
        .O(\u0/out4 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__320
       (.I0(\u2/u8/X [17]),
        .I1(\u2/u8/X [16]),
        .I2(\u2/u8/X [15]),
        .I3(\u2/u8/X [14]),
        .I4(\u2/u8/X [18]),
        .I5(\u2/u8/X [13]),
        .O(\u2/out8 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__321
       (.I0(\u2/u8/X [35]),
        .I1(\u2/u8/X [34]),
        .I2(\u2/u8/X [33]),
        .I3(\u2/u8/X [32]),
        .I4(\u2/u8/X [36]),
        .I5(\u2/u8/X [31]),
        .O(\u2/out8 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__322
       (.I0(\u2/u8/X [11]),
        .I1(\u2/u8/X [10]),
        .I2(\u2/u8/X [9]),
        .I3(\u2/u8/X [8]),
        .I4(\u2/u8/X [12]),
        .I5(\u2/u8/X [7]),
        .O(\u2/out8 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__323
       (.I0(\u2/u8/X [47]),
        .I1(\u2/u8/X [46]),
        .I2(\u2/u8/X [45]),
        .I3(\u2/u8/X [44]),
        .I4(\u2/u8/X [48]),
        .I5(\u2/u8/X [43]),
        .O(\u2/out8 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__324
       (.I0(\u2/u8/X [23]),
        .I1(\u2/u8/X [22]),
        .I2(\u2/u8/X [21]),
        .I3(\u2/u8/X [20]),
        .I4(\u2/u8/X [24]),
        .I5(\u2/u8/X [19]),
        .O(\u2/out8 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__325
       (.I0(\u2/u8/X [29]),
        .I1(\u2/u8/X [28]),
        .I2(\u2/u8/X [27]),
        .I3(\u2/u8/X [26]),
        .I4(\u2/u8/X [30]),
        .I5(\u2/u8/X [25]),
        .O(\u2/out8 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__326
       (.I0(\u2/u8/X [5]),
        .I1(\u2/u8/X [4]),
        .I2(\u2/u8/X [3]),
        .I3(\u2/u8/X [2]),
        .I4(\u2/u8/X [6]),
        .I5(\u2/u8/X [1]),
        .O(\u2/out8 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__327
       (.I0(\u2/u9/X [41]),
        .I1(\u2/u9/X [40]),
        .I2(\u2/u9/X [39]),
        .I3(\u2/u9/X [38]),
        .I4(\u2/u9/X [42]),
        .I5(\u2/u9/X [37]),
        .O(\u2/out9 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__328
       (.I0(\u2/u9/X [17]),
        .I1(\u2/u9/X [16]),
        .I2(\u2/u9/X [15]),
        .I3(\u2/u9/X [14]),
        .I4(\u2/u9/X [18]),
        .I5(\u2/u9/X [13]),
        .O(\u2/out9 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__329
       (.I0(\u2/u9/X [35]),
        .I1(\u2/u9/X [34]),
        .I2(\u2/u9/X [33]),
        .I3(\u2/u9/X [32]),
        .I4(\u2/u9/X [36]),
        .I5(\u2/u9/X [31]),
        .O(\u2/out9 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__33
       (.I0(\u0/u4/X [35]),
        .I1(\u0/u4/X [34]),
        .I2(\u0/u4/X [33]),
        .I3(\u0/u4/X [32]),
        .I4(\u0/u4/X [36]),
        .I5(\u0/u4/X [31]),
        .O(\u0/out4 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__330
       (.I0(\u2/u9/X [11]),
        .I1(\u2/u9/X [10]),
        .I2(\u2/u9/X [9]),
        .I3(\u2/u9/X [8]),
        .I4(\u2/u9/X [12]),
        .I5(\u2/u9/X [7]),
        .O(\u2/out9 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__331
       (.I0(\u2/u9/X [47]),
        .I1(\u2/u9/X [46]),
        .I2(\u2/u9/X [45]),
        .I3(\u2/u9/X [44]),
        .I4(\u2/u9/X [48]),
        .I5(\u2/u9/X [43]),
        .O(\u2/out9 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__332
       (.I0(\u2/u9/X [23]),
        .I1(\u2/u9/X [22]),
        .I2(\u2/u9/X [21]),
        .I3(\u2/u9/X [20]),
        .I4(\u2/u9/X [24]),
        .I5(\u2/u9/X [19]),
        .O(\u2/out9 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__333
       (.I0(\u2/u9/X [29]),
        .I1(\u2/u9/X [28]),
        .I2(\u2/u9/X [27]),
        .I3(\u2/u9/X [26]),
        .I4(\u2/u9/X [30]),
        .I5(\u2/u9/X [25]),
        .O(\u2/out9 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__334
       (.I0(\u2/u9/X [5]),
        .I1(\u2/u9/X [4]),
        .I2(\u2/u9/X [3]),
        .I3(\u2/u9/X [2]),
        .I4(\u2/u9/X [6]),
        .I5(\u2/u9/X [1]),
        .O(\u2/out9 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__335
       (.I0(\u2/u10/X [41]),
        .I1(\u2/u10/X [40]),
        .I2(\u2/u10/X [39]),
        .I3(\u2/u10/X [38]),
        .I4(\u2/u10/X [42]),
        .I5(\u2/u10/X [37]),
        .O(\u2/out10 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__336
       (.I0(\u2/u10/X [17]),
        .I1(\u2/u10/X [16]),
        .I2(\u2/u10/X [15]),
        .I3(\u2/u10/X [14]),
        .I4(\u2/u10/X [18]),
        .I5(\u2/u10/X [13]),
        .O(\u2/out10 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__337
       (.I0(\u2/u10/X [35]),
        .I1(\u2/u10/X [34]),
        .I2(\u2/u10/X [33]),
        .I3(\u2/u10/X [32]),
        .I4(\u2/u10/X [36]),
        .I5(\u2/u10/X [31]),
        .O(\u2/out10 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__338
       (.I0(\u2/u10/X [11]),
        .I1(\u2/u10/X [10]),
        .I2(\u2/u10/X [9]),
        .I3(\u2/u10/X [8]),
        .I4(\u2/u10/X [12]),
        .I5(\u2/u10/X [7]),
        .O(\u2/out10 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__339
       (.I0(\u2/u10/X [47]),
        .I1(\u2/u10/X [46]),
        .I2(\u2/u10/X [45]),
        .I3(\u2/u10/X [44]),
        .I4(\u2/u10/X [48]),
        .I5(\u2/u10/X [43]),
        .O(\u2/out10 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__34
       (.I0(\u0/u4/X [11]),
        .I1(\u0/u4/X [10]),
        .I2(\u0/u4/X [9]),
        .I3(\u0/u4/X [8]),
        .I4(\u0/u4/X [12]),
        .I5(\u0/u4/X [7]),
        .O(\u0/out4 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__340
       (.I0(\u2/u10/X [23]),
        .I1(\u2/u10/X [22]),
        .I2(\u2/u10/X [21]),
        .I3(\u2/u10/X [20]),
        .I4(\u2/u10/X [24]),
        .I5(\u2/u10/X [19]),
        .O(\u2/out10 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__341
       (.I0(\u2/u10/X [29]),
        .I1(\u2/u10/X [28]),
        .I2(\u2/u10/X [27]),
        .I3(\u2/u10/X [26]),
        .I4(\u2/u10/X [30]),
        .I5(\u2/u10/X [25]),
        .O(\u2/out10 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__342
       (.I0(\u2/u10/X [5]),
        .I1(\u2/u10/X [4]),
        .I2(\u2/u10/X [3]),
        .I3(\u2/u10/X [2]),
        .I4(\u2/u10/X [6]),
        .I5(\u2/u10/X [1]),
        .O(\u2/out10 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__343
       (.I0(\u2/u11/X [41]),
        .I1(\u2/u11/X [40]),
        .I2(\u2/u11/X [39]),
        .I3(\u2/u11/X [38]),
        .I4(\u2/u11/X [42]),
        .I5(\u2/u11/X [37]),
        .O(\u2/out11 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__344
       (.I0(\u2/u11/X [17]),
        .I1(\u2/u11/X [16]),
        .I2(\u2/u11/X [15]),
        .I3(\u2/u11/X [14]),
        .I4(\u2/u11/X [18]),
        .I5(\u2/u11/X [13]),
        .O(\u2/out11 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__345
       (.I0(\u2/u11/X [35]),
        .I1(\u2/u11/X [34]),
        .I2(\u2/u11/X [33]),
        .I3(\u2/u11/X [32]),
        .I4(\u2/u11/X [36]),
        .I5(\u2/u11/X [31]),
        .O(\u2/out11 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__346
       (.I0(\u2/u11/X [11]),
        .I1(\u2/u11/X [10]),
        .I2(\u2/u11/X [9]),
        .I3(\u2/u11/X [8]),
        .I4(\u2/u11/X [12]),
        .I5(\u2/u11/X [7]),
        .O(\u2/out11 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__347
       (.I0(\u2/u11/X [47]),
        .I1(\u2/u11/X [46]),
        .I2(\u2/u11/X [45]),
        .I3(\u2/u11/X [44]),
        .I4(\u2/u11/X [48]),
        .I5(\u2/u11/X [43]),
        .O(\u2/out11 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__348
       (.I0(\u2/u11/X [23]),
        .I1(\u2/u11/X [22]),
        .I2(\u2/u11/X [21]),
        .I3(\u2/u11/X [20]),
        .I4(\u2/u11/X [24]),
        .I5(\u2/u11/X [19]),
        .O(\u2/out11 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__349
       (.I0(\u2/u11/X [29]),
        .I1(\u2/u11/X [28]),
        .I2(\u2/u11/X [27]),
        .I3(\u2/u11/X [26]),
        .I4(\u2/u11/X [30]),
        .I5(\u2/u11/X [25]),
        .O(\u2/out11 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__35
       (.I0(\u0/u4/X [47]),
        .I1(\u0/u4/X [46]),
        .I2(\u0/u4/X [45]),
        .I3(\u0/u4/X [44]),
        .I4(\u0/u4/X [48]),
        .I5(\u0/u4/X [43]),
        .O(\u0/out4 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__350
       (.I0(\u2/u11/X [5]),
        .I1(\u2/u11/X [4]),
        .I2(\u2/u11/X [3]),
        .I3(\u2/u11/X [2]),
        .I4(\u2/u11/X [6]),
        .I5(\u2/u11/X [1]),
        .O(\u2/out11 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__351
       (.I0(\u2/u12/X [41]),
        .I1(\u2/u12/X [40]),
        .I2(\u2/u12/X [39]),
        .I3(\u2/u12/X [38]),
        .I4(\u2/u12/X [42]),
        .I5(\u2/u12/X [37]),
        .O(\u2/out12 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__352
       (.I0(\u2/u12/X [17]),
        .I1(\u2/u12/X [16]),
        .I2(\u2/u12/X [15]),
        .I3(\u2/u12/X [14]),
        .I4(\u2/u12/X [18]),
        .I5(\u2/u12/X [13]),
        .O(\u2/out12 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__353
       (.I0(\u2/u12/X [35]),
        .I1(\u2/u12/X [34]),
        .I2(\u2/u12/X [33]),
        .I3(\u2/u12/X [32]),
        .I4(\u2/u12/X [36]),
        .I5(\u2/u12/X [31]),
        .O(\u2/out12 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__354
       (.I0(\u2/u12/X [11]),
        .I1(\u2/u12/X [10]),
        .I2(\u2/u12/X [9]),
        .I3(\u2/u12/X [8]),
        .I4(\u2/u12/X [12]),
        .I5(\u2/u12/X [7]),
        .O(\u2/out12 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__355
       (.I0(\u2/u12/X [47]),
        .I1(\u2/u12/X [46]),
        .I2(\u2/u12/X [45]),
        .I3(\u2/u12/X [44]),
        .I4(\u2/u12/X [48]),
        .I5(\u2/u12/X [43]),
        .O(\u2/out12 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__356
       (.I0(\u2/u12/X [23]),
        .I1(\u2/u12/X [22]),
        .I2(\u2/u12/X [21]),
        .I3(\u2/u12/X [20]),
        .I4(\u2/u12/X [24]),
        .I5(\u2/u12/X [19]),
        .O(\u2/out12 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__357
       (.I0(\u2/u12/X [29]),
        .I1(\u2/u12/X [28]),
        .I2(\u2/u12/X [27]),
        .I3(\u2/u12/X [26]),
        .I4(\u2/u12/X [30]),
        .I5(\u2/u12/X [25]),
        .O(\u2/out12 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__358
       (.I0(\u2/u12/X [5]),
        .I1(\u2/u12/X [4]),
        .I2(\u2/u12/X [3]),
        .I3(\u2/u12/X [2]),
        .I4(\u2/u12/X [6]),
        .I5(\u2/u12/X [1]),
        .O(\u2/out12 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__359
       (.I0(\u2/u13/X [41]),
        .I1(\u2/u13/X [40]),
        .I2(\u2/u13/X [39]),
        .I3(\u2/u13/X [38]),
        .I4(\u2/u13/X [42]),
        .I5(\u2/u13/X [37]),
        .O(\u2/out13 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__36
       (.I0(\u0/u4/X [23]),
        .I1(\u0/u4/X [22]),
        .I2(\u0/u4/X [21]),
        .I3(\u0/u4/X [20]),
        .I4(\u0/u4/X [24]),
        .I5(\u0/u4/X [19]),
        .O(\u0/out4 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__360
       (.I0(\u2/u13/X [17]),
        .I1(\u2/u13/X [16]),
        .I2(\u2/u13/X [15]),
        .I3(\u2/u13/X [14]),
        .I4(\u2/u13/X [18]),
        .I5(\u2/u13/X [13]),
        .O(\u2/out13 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__361
       (.I0(\u2/u13/X [35]),
        .I1(\u2/u13/X [34]),
        .I2(\u2/u13/X [33]),
        .I3(\u2/u13/X [32]),
        .I4(\u2/u13/X [36]),
        .I5(\u2/u13/X [31]),
        .O(\u2/out13 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__362
       (.I0(\u2/u13/X [11]),
        .I1(\u2/u13/X [10]),
        .I2(\u2/u13/X [9]),
        .I3(\u2/u13/X [8]),
        .I4(\u2/u13/X [12]),
        .I5(\u2/u13/X [7]),
        .O(\u2/out13 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__363
       (.I0(\u2/u13/X [47]),
        .I1(\u2/u13/X [46]),
        .I2(\u2/u13/X [45]),
        .I3(\u2/u13/X [44]),
        .I4(\u2/u13/X [48]),
        .I5(\u2/u13/X [43]),
        .O(\u2/out13 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__364
       (.I0(\u2/u13/X [23]),
        .I1(\u2/u13/X [22]),
        .I2(\u2/u13/X [21]),
        .I3(\u2/u13/X [20]),
        .I4(\u2/u13/X [24]),
        .I5(\u2/u13/X [19]),
        .O(\u2/out13 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__365
       (.I0(\u2/u13/X [29]),
        .I1(\u2/u13/X [28]),
        .I2(\u2/u13/X [27]),
        .I3(\u2/u13/X [26]),
        .I4(\u2/u13/X [30]),
        .I5(\u2/u13/X [25]),
        .O(\u2/out13 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__366
       (.I0(\u2/u13/X [5]),
        .I1(\u2/u13/X [4]),
        .I2(\u2/u13/X [3]),
        .I3(\u2/u13/X [2]),
        .I4(\u2/u13/X [6]),
        .I5(\u2/u13/X [1]),
        .O(\u2/out13 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__367
       (.I0(\u2/u14/X [41]),
        .I1(\u2/u14/X [40]),
        .I2(\u2/u14/X [39]),
        .I3(\u2/u14/X [38]),
        .I4(\u2/u14/X [42]),
        .I5(\u2/u14/X [37]),
        .O(\u2/out14 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__368
       (.I0(\u2/u14/X [17]),
        .I1(\u2/u14/X [16]),
        .I2(\u2/u14/X [15]),
        .I3(\u2/u14/X [14]),
        .I4(\u2/u14/X [18]),
        .I5(\u2/u14/X [13]),
        .O(\u2/out14 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__369
       (.I0(\u2/u14/X [35]),
        .I1(\u2/u14/X [34]),
        .I2(\u2/u14/X [33]),
        .I3(\u2/u14/X [32]),
        .I4(\u2/u14/X [36]),
        .I5(\u2/u14/X [31]),
        .O(\u2/out14 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__37
       (.I0(\u0/u4/X [29]),
        .I1(\u0/u4/X [28]),
        .I2(\u0/u4/X [27]),
        .I3(\u0/u4/X [26]),
        .I4(\u0/u4/X [30]),
        .I5(\u0/u4/X [25]),
        .O(\u0/out4 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__370
       (.I0(\u2/u14/X [11]),
        .I1(\u2/u14/X [10]),
        .I2(\u2/u14/X [9]),
        .I3(\u2/u14/X [8]),
        .I4(\u2/u14/X [12]),
        .I5(\u2/u14/X [7]),
        .O(\u2/out14 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__371
       (.I0(\u2/u14/X [47]),
        .I1(\u2/u14/X [46]),
        .I2(\u2/u14/X [45]),
        .I3(\u2/u14/X [44]),
        .I4(\u2/u14/X [48]),
        .I5(\u2/u14/X [43]),
        .O(\u2/out14 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__372
       (.I0(\u2/u14/X [23]),
        .I1(\u2/u14/X [22]),
        .I2(\u2/u14/X [21]),
        .I3(\u2/u14/X [20]),
        .I4(\u2/u14/X [24]),
        .I5(\u2/u14/X [19]),
        .O(\u2/out14 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__373
       (.I0(\u2/u14/X [29]),
        .I1(\u2/u14/X [28]),
        .I2(\u2/u14/X [27]),
        .I3(\u2/u14/X [26]),
        .I4(\u2/u14/X [30]),
        .I5(\u2/u14/X [25]),
        .O(\u2/out14 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__374
       (.I0(\u2/u14/X [5]),
        .I1(\u2/u14/X [4]),
        .I2(\u2/u14/X [3]),
        .I3(\u2/u14/X [2]),
        .I4(\u2/u14/X [6]),
        .I5(\u2/u14/X [1]),
        .O(\u2/out14 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__375
       (.I0(\u2/u15/X [41]),
        .I1(\u2/u15/X [40]),
        .I2(\u2/u15/X [39]),
        .I3(\u2/u15/X [38]),
        .I4(\u2/u15/X [42]),
        .I5(\u2/u15/X [37]),
        .O(\u2/out15 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__376
       (.I0(\u2/u15/X [17]),
        .I1(\u2/u15/X [16]),
        .I2(\u2/u15/X [15]),
        .I3(\u2/u15/X [14]),
        .I4(\u2/u15/X [18]),
        .I5(\u2/u15/X [13]),
        .O(\u2/out15 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__377
       (.I0(\u2/u15/X [35]),
        .I1(\u2/u15/X [34]),
        .I2(\u2/u15/X [33]),
        .I3(\u2/u15/X [32]),
        .I4(\u2/u15/X [36]),
        .I5(\u2/u15/X [31]),
        .O(\u2/out15 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__378
       (.I0(\u2/u15/X [11]),
        .I1(\u2/u15/X [10]),
        .I2(\u2/u15/X [9]),
        .I3(\u2/u15/X [8]),
        .I4(\u2/u15/X [12]),
        .I5(\u2/u15/X [7]),
        .O(\u2/out15 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__379
       (.I0(\u2/u15/X [47]),
        .I1(\u2/u15/X [46]),
        .I2(\u2/u15/X [45]),
        .I3(\u2/u15/X [44]),
        .I4(\u2/u15/X [48]),
        .I5(\u2/u15/X [43]),
        .O(\u2/out15 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__38
       (.I0(\u0/u4/X [5]),
        .I1(\u0/u4/X [4]),
        .I2(\u0/u4/X [3]),
        .I3(\u0/u4/X [2]),
        .I4(\u0/u4/X [6]),
        .I5(\u0/u4/X [1]),
        .O(\u0/out4 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__380
       (.I0(\u2/u15/X [23]),
        .I1(\u2/u15/X [22]),
        .I2(\u2/u15/X [21]),
        .I3(\u2/u15/X [20]),
        .I4(\u2/u15/X [24]),
        .I5(\u2/u15/X [19]),
        .O(\u2/out15 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__381
       (.I0(\u2/u15/X [29]),
        .I1(\u2/u15/X [28]),
        .I2(\u2/u15/X [27]),
        .I3(\u2/u15/X [26]),
        .I4(\u2/u15/X [30]),
        .I5(\u2/u15/X [25]),
        .O(\u2/out15 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__382
       (.I0(\u2/u15/X [5]),
        .I1(\u2/u15/X [4]),
        .I2(\u2/u15/X [3]),
        .I3(\u2/u15/X [2]),
        .I4(\u2/u15/X [6]),
        .I5(\u2/u15/X [1]),
        .O(\u2/out15 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__39
       (.I0(\u0/u5/X [41]),
        .I1(\u0/u5/X [40]),
        .I2(\u0/u5/X [39]),
        .I3(\u0/u5/X [38]),
        .I4(\u0/u5/X [42]),
        .I5(\u0/u5/X [37]),
        .O(\u0/out5 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__4
       (.I0(\u0/u0/X [23]),
        .I1(\u0/u0/X [22]),
        .I2(\u0/u0/X [21]),
        .I3(\u0/u0/X [20]),
        .I4(\u0/u0/X [24]),
        .I5(\u0/u0/X [19]),
        .O(\u0/out0 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__40
       (.I0(\u0/u5/X [17]),
        .I1(\u0/u5/X [16]),
        .I2(\u0/u5/X [15]),
        .I3(\u0/u5/X [14]),
        .I4(\u0/u5/X [18]),
        .I5(\u0/u5/X [13]),
        .O(\u0/out5 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__41
       (.I0(\u0/u5/X [35]),
        .I1(\u0/u5/X [34]),
        .I2(\u0/u5/X [33]),
        .I3(\u0/u5/X [32]),
        .I4(\u0/u5/X [36]),
        .I5(\u0/u5/X [31]),
        .O(\u0/out5 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__42
       (.I0(\u0/u5/X [11]),
        .I1(\u0/u5/X [10]),
        .I2(\u0/u5/X [9]),
        .I3(\u0/u5/X [8]),
        .I4(\u0/u5/X [12]),
        .I5(\u0/u5/X [7]),
        .O(\u0/out5 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__43
       (.I0(\u0/u5/X [47]),
        .I1(\u0/u5/X [46]),
        .I2(\u0/u5/X [45]),
        .I3(\u0/u5/X [44]),
        .I4(\u0/u5/X [48]),
        .I5(\u0/u5/X [43]),
        .O(\u0/out5 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__44
       (.I0(\u0/u5/X [23]),
        .I1(\u0/u5/X [22]),
        .I2(\u0/u5/X [21]),
        .I3(\u0/u5/X [20]),
        .I4(\u0/u5/X [24]),
        .I5(\u0/u5/X [19]),
        .O(\u0/out5 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__45
       (.I0(\u0/u5/X [29]),
        .I1(\u0/u5/X [28]),
        .I2(\u0/u5/X [27]),
        .I3(\u0/u5/X [26]),
        .I4(\u0/u5/X [30]),
        .I5(\u0/u5/X [25]),
        .O(\u0/out5 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__46
       (.I0(\u0/u5/X [5]),
        .I1(\u0/u5/X [4]),
        .I2(\u0/u5/X [3]),
        .I3(\u0/u5/X [2]),
        .I4(\u0/u5/X [6]),
        .I5(\u0/u5/X [1]),
        .O(\u0/out5 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__47
       (.I0(\u0/u6/X [41]),
        .I1(\u0/u6/X [40]),
        .I2(\u0/u6/X [39]),
        .I3(\u0/u6/X [38]),
        .I4(\u0/u6/X [42]),
        .I5(\u0/u6/X [37]),
        .O(\u0/out6 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__48
       (.I0(\u0/u6/X [17]),
        .I1(\u0/u6/X [16]),
        .I2(\u0/u6/X [15]),
        .I3(\u0/u6/X [14]),
        .I4(\u0/u6/X [18]),
        .I5(\u0/u6/X [13]),
        .O(\u0/out6 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__49
       (.I0(\u0/u6/X [35]),
        .I1(\u0/u6/X [34]),
        .I2(\u0/u6/X [33]),
        .I3(\u0/u6/X [32]),
        .I4(\u0/u6/X [36]),
        .I5(\u0/u6/X [31]),
        .O(\u0/out6 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__5
       (.I0(\u0/u0/X [29]),
        .I1(\u0/u0/X [28]),
        .I2(\u0/u0/X [27]),
        .I3(\u0/u0/X [26]),
        .I4(\u0/u0/X [30]),
        .I5(\u0/u0/X [25]),
        .O(\u0/out0 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__50
       (.I0(\u0/u6/X [11]),
        .I1(\u0/u6/X [10]),
        .I2(\u0/u6/X [9]),
        .I3(\u0/u6/X [8]),
        .I4(\u0/u6/X [12]),
        .I5(\u0/u6/X [7]),
        .O(\u0/out6 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__51
       (.I0(\u0/u6/X [47]),
        .I1(\u0/u6/X [46]),
        .I2(\u0/u6/X [45]),
        .I3(\u0/u6/X [44]),
        .I4(\u0/u6/X [48]),
        .I5(\u0/u6/X [43]),
        .O(\u0/out6 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__52
       (.I0(\u0/u6/X [23]),
        .I1(\u0/u6/X [22]),
        .I2(\u0/u6/X [21]),
        .I3(\u0/u6/X [20]),
        .I4(\u0/u6/X [24]),
        .I5(\u0/u6/X [19]),
        .O(\u0/out6 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__53
       (.I0(\u0/u6/X [29]),
        .I1(\u0/u6/X [28]),
        .I2(\u0/u6/X [27]),
        .I3(\u0/u6/X [26]),
        .I4(\u0/u6/X [30]),
        .I5(\u0/u6/X [25]),
        .O(\u0/out6 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__54
       (.I0(\u0/u6/X [5]),
        .I1(\u0/u6/X [4]),
        .I2(\u0/u6/X [3]),
        .I3(\u0/u6/X [2]),
        .I4(\u0/u6/X [6]),
        .I5(\u0/u6/X [1]),
        .O(\u0/out6 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__55
       (.I0(\u0/u7/X [41]),
        .I1(\u0/u7/X [40]),
        .I2(\u0/u7/X [39]),
        .I3(\u0/u7/X [38]),
        .I4(\u0/u7/X [42]),
        .I5(\u0/u7/X [37]),
        .O(\u0/out7 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__56
       (.I0(\u0/u7/X [17]),
        .I1(\u0/u7/X [16]),
        .I2(\u0/u7/X [15]),
        .I3(\u0/u7/X [14]),
        .I4(\u0/u7/X [18]),
        .I5(\u0/u7/X [13]),
        .O(\u0/out7 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__57
       (.I0(\u0/u7/X [35]),
        .I1(\u0/u7/X [34]),
        .I2(\u0/u7/X [33]),
        .I3(\u0/u7/X [32]),
        .I4(\u0/u7/X [36]),
        .I5(\u0/u7/X [31]),
        .O(\u0/out7 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__58
       (.I0(\u0/u7/X [11]),
        .I1(\u0/u7/X [10]),
        .I2(\u0/u7/X [9]),
        .I3(\u0/u7/X [8]),
        .I4(\u0/u7/X [12]),
        .I5(\u0/u7/X [7]),
        .O(\u0/out7 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__59
       (.I0(\u0/u7/X [47]),
        .I1(\u0/u7/X [46]),
        .I2(\u0/u7/X [45]),
        .I3(\u0/u7/X [44]),
        .I4(\u0/u7/X [48]),
        .I5(\u0/u7/X [43]),
        .O(\u0/out7 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__6
       (.I0(\u0/u0/X [5]),
        .I1(\u0/u0/X [4]),
        .I2(\u0/u0/X [3]),
        .I3(\u0/u0/X [2]),
        .I4(\u0/u0/X [6]),
        .I5(\u0/u0/X [1]),
        .O(\u0/out0 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__60
       (.I0(\u0/u7/X [23]),
        .I1(\u0/u7/X [22]),
        .I2(\u0/u7/X [21]),
        .I3(\u0/u7/X [20]),
        .I4(\u0/u7/X [24]),
        .I5(\u0/u7/X [19]),
        .O(\u0/out7 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__61
       (.I0(\u0/u7/X [29]),
        .I1(\u0/u7/X [28]),
        .I2(\u0/u7/X [27]),
        .I3(\u0/u7/X [26]),
        .I4(\u0/u7/X [30]),
        .I5(\u0/u7/X [25]),
        .O(\u0/out7 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__62
       (.I0(\u0/u7/X [5]),
        .I1(\u0/u7/X [4]),
        .I2(\u0/u7/X [3]),
        .I3(\u0/u7/X [2]),
        .I4(\u0/u7/X [6]),
        .I5(\u0/u7/X [1]),
        .O(\u0/out7 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__63
       (.I0(\u0/u8/X [41]),
        .I1(\u0/u8/X [40]),
        .I2(\u0/u8/X [39]),
        .I3(\u0/u8/X [38]),
        .I4(\u0/u8/X [42]),
        .I5(\u0/u8/X [37]),
        .O(\u0/out8 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__64
       (.I0(\u0/u8/X [17]),
        .I1(\u0/u8/X [16]),
        .I2(\u0/u8/X [15]),
        .I3(\u0/u8/X [14]),
        .I4(\u0/u8/X [18]),
        .I5(\u0/u8/X [13]),
        .O(\u0/out8 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__65
       (.I0(\u0/u8/X [35]),
        .I1(\u0/u8/X [34]),
        .I2(\u0/u8/X [33]),
        .I3(\u0/u8/X [32]),
        .I4(\u0/u8/X [36]),
        .I5(\u0/u8/X [31]),
        .O(\u0/out8 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__66
       (.I0(\u0/u8/X [11]),
        .I1(\u0/u8/X [10]),
        .I2(\u0/u8/X [9]),
        .I3(\u0/u8/X [8]),
        .I4(\u0/u8/X [12]),
        .I5(\u0/u8/X [7]),
        .O(\u0/out8 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__67
       (.I0(\u0/u8/X [47]),
        .I1(\u0/u8/X [46]),
        .I2(\u0/u8/X [45]),
        .I3(\u0/u8/X [44]),
        .I4(\u0/u8/X [48]),
        .I5(\u0/u8/X [43]),
        .O(\u0/out8 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__68
       (.I0(\u0/u8/X [23]),
        .I1(\u0/u8/X [22]),
        .I2(\u0/u8/X [21]),
        .I3(\u0/u8/X [20]),
        .I4(\u0/u8/X [24]),
        .I5(\u0/u8/X [19]),
        .O(\u0/out8 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__69
       (.I0(\u0/u8/X [29]),
        .I1(\u0/u8/X [28]),
        .I2(\u0/u8/X [27]),
        .I3(\u0/u8/X [26]),
        .I4(\u0/u8/X [30]),
        .I5(\u0/u8/X [25]),
        .O(\u0/out8 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__7
       (.I0(\u0/u1/X [41]),
        .I1(\u0/u1/X [40]),
        .I2(\u0/u1/X [39]),
        .I3(\u0/u1/X [38]),
        .I4(\u0/u1/X [42]),
        .I5(\u0/u1/X [37]),
        .O(\u0/out1 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__70
       (.I0(\u0/u8/X [5]),
        .I1(\u0/u8/X [4]),
        .I2(\u0/u8/X [3]),
        .I3(\u0/u8/X [2]),
        .I4(\u0/u8/X [6]),
        .I5(\u0/u8/X [1]),
        .O(\u0/out8 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__71
       (.I0(\u0/u9/X [41]),
        .I1(\u0/u9/X [40]),
        .I2(\u0/u9/X [39]),
        .I3(\u0/u9/X [38]),
        .I4(\u0/u9/X [42]),
        .I5(\u0/u9/X [37]),
        .O(\u0/out9 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__72
       (.I0(\u0/u9/X [17]),
        .I1(\u0/u9/X [16]),
        .I2(\u0/u9/X [15]),
        .I3(\u0/u9/X [14]),
        .I4(\u0/u9/X [18]),
        .I5(\u0/u9/X [13]),
        .O(\u0/out9 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__73
       (.I0(\u0/u9/X [35]),
        .I1(\u0/u9/X [34]),
        .I2(\u0/u9/X [33]),
        .I3(\u0/u9/X [32]),
        .I4(\u0/u9/X [36]),
        .I5(\u0/u9/X [31]),
        .O(\u0/out9 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__74
       (.I0(\u0/u9/X [11]),
        .I1(\u0/u9/X [10]),
        .I2(\u0/u9/X [9]),
        .I3(\u0/u9/X [8]),
        .I4(\u0/u9/X [12]),
        .I5(\u0/u9/X [7]),
        .O(\u0/out9 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__75
       (.I0(\u0/u9/X [47]),
        .I1(\u0/u9/X [46]),
        .I2(\u0/u9/X [45]),
        .I3(\u0/u9/X [44]),
        .I4(\u0/u9/X [48]),
        .I5(\u0/u9/X [43]),
        .O(\u0/out9 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__76
       (.I0(\u0/u9/X [23]),
        .I1(\u0/u9/X [22]),
        .I2(\u0/u9/X [21]),
        .I3(\u0/u9/X [20]),
        .I4(\u0/u9/X [24]),
        .I5(\u0/u9/X [19]),
        .O(\u0/out9 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__77
       (.I0(\u0/u9/X [29]),
        .I1(\u0/u9/X [28]),
        .I2(\u0/u9/X [27]),
        .I3(\u0/u9/X [26]),
        .I4(\u0/u9/X [30]),
        .I5(\u0/u9/X [25]),
        .O(\u0/out9 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__78
       (.I0(\u0/u9/X [5]),
        .I1(\u0/u9/X [4]),
        .I2(\u0/u9/X [3]),
        .I3(\u0/u9/X [2]),
        .I4(\u0/u9/X [6]),
        .I5(\u0/u9/X [1]),
        .O(\u0/out9 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__79
       (.I0(\u0/u10/X [41]),
        .I1(\u0/u10/X [40]),
        .I2(\u0/u10/X [39]),
        .I3(\u0/u10/X [38]),
        .I4(\u0/u10/X [42]),
        .I5(\u0/u10/X [37]),
        .O(\u0/out10 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__8
       (.I0(\u0/u1/X [17]),
        .I1(\u0/u1/X [16]),
        .I2(\u0/u1/X [15]),
        .I3(\u0/u1/X [14]),
        .I4(\u0/u1/X [18]),
        .I5(\u0/u1/X [13]),
        .O(\u0/out1 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__80
       (.I0(\u0/u10/X [17]),
        .I1(\u0/u10/X [16]),
        .I2(\u0/u10/X [15]),
        .I3(\u0/u10/X [14]),
        .I4(\u0/u10/X [18]),
        .I5(\u0/u10/X [13]),
        .O(\u0/out10 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__81
       (.I0(\u0/u10/X [35]),
        .I1(\u0/u10/X [34]),
        .I2(\u0/u10/X [33]),
        .I3(\u0/u10/X [32]),
        .I4(\u0/u10/X [36]),
        .I5(\u0/u10/X [31]),
        .O(\u0/out10 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__82
       (.I0(\u0/u10/X [11]),
        .I1(\u0/u10/X [10]),
        .I2(\u0/u10/X [9]),
        .I3(\u0/u10/X [8]),
        .I4(\u0/u10/X [12]),
        .I5(\u0/u10/X [7]),
        .O(\u0/out10 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__83
       (.I0(\u0/u10/X [47]),
        .I1(\u0/u10/X [46]),
        .I2(\u0/u10/X [45]),
        .I3(\u0/u10/X [44]),
        .I4(\u0/u10/X [48]),
        .I5(\u0/u10/X [43]),
        .O(\u0/out10 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__84
       (.I0(\u0/u10/X [23]),
        .I1(\u0/u10/X [22]),
        .I2(\u0/u10/X [21]),
        .I3(\u0/u10/X [20]),
        .I4(\u0/u10/X [24]),
        .I5(\u0/u10/X [19]),
        .O(\u0/out10 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__85
       (.I0(\u0/u10/X [29]),
        .I1(\u0/u10/X [28]),
        .I2(\u0/u10/X [27]),
        .I3(\u0/u10/X [26]),
        .I4(\u0/u10/X [30]),
        .I5(\u0/u10/X [25]),
        .O(\u0/out10 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__86
       (.I0(\u0/u10/X [5]),
        .I1(\u0/u10/X [4]),
        .I2(\u0/u10/X [3]),
        .I3(\u0/u10/X [2]),
        .I4(\u0/u10/X [6]),
        .I5(\u0/u10/X [1]),
        .O(\u0/out10 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__87
       (.I0(\u0/u11/X [41]),
        .I1(\u0/u11/X [40]),
        .I2(\u0/u11/X [39]),
        .I3(\u0/u11/X [38]),
        .I4(\u0/u11/X [42]),
        .I5(\u0/u11/X [37]),
        .O(\u0/out11 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__88
       (.I0(\u0/u11/X [17]),
        .I1(\u0/u11/X [16]),
        .I2(\u0/u11/X [15]),
        .I3(\u0/u11/X [14]),
        .I4(\u0/u11/X [18]),
        .I5(\u0/u11/X [13]),
        .O(\u0/out11 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__89
       (.I0(\u0/u11/X [35]),
        .I1(\u0/u11/X [34]),
        .I2(\u0/u11/X [33]),
        .I3(\u0/u11/X [32]),
        .I4(\u0/u11/X [36]),
        .I5(\u0/u11/X [31]),
        .O(\u0/out11 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__9
       (.I0(\u0/u1/X [35]),
        .I1(\u0/u1/X [34]),
        .I2(\u0/u1/X [33]),
        .I3(\u0/u1/X [32]),
        .I4(\u0/u1/X [36]),
        .I5(\u0/u1/X [31]),
        .O(\u0/out1 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__90
       (.I0(\u0/u11/X [11]),
        .I1(\u0/u11/X [10]),
        .I2(\u0/u11/X [9]),
        .I3(\u0/u11/X [8]),
        .I4(\u0/u11/X [12]),
        .I5(\u0/u11/X [7]),
        .O(\u0/out11 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__91
       (.I0(\u0/u11/X [47]),
        .I1(\u0/u11/X [46]),
        .I2(\u0/u11/X [45]),
        .I3(\u0/u11/X [44]),
        .I4(\u0/u11/X [48]),
        .I5(\u0/u11/X [43]),
        .O(\u0/out11 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE81B2D6366B492AD)) 
    g0_b1__92
       (.I0(\u0/u11/X [23]),
        .I1(\u0/u11/X [22]),
        .I2(\u0/u11/X [21]),
        .I3(\u0/u11/X [20]),
        .I4(\u0/u11/X [24]),
        .I5(\u0/u11/X [19]),
        .O(\u0/out11 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9369B15A9C274CF1)) 
    g0_b1__93
       (.I0(\u0/u11/X [29]),
        .I1(\u0/u11/X [28]),
        .I2(\u0/u11/X [27]),
        .I3(\u0/u11/X [26]),
        .I4(\u0/u11/X [30]),
        .I5(\u0/u11/X [25]),
        .O(\u0/out11 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E8939E44B368771)) 
    g0_b1__94
       (.I0(\u0/u11/X [5]),
        .I1(\u0/u11/X [4]),
        .I2(\u0/u11/X [3]),
        .I3(\u0/u11/X [2]),
        .I4(\u0/u11/X [6]),
        .I5(\u0/u11/X [1]),
        .O(\u0/out11 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h78C387E4B38C691E)) 
    g0_b1__95
       (.I0(\u0/u12/X [41]),
        .I1(\u0/u12/X [40]),
        .I2(\u0/u12/X [39]),
        .I3(\u0/u12/X [38]),
        .I4(\u0/u12/X [42]),
        .I5(\u0/u12/X [37]),
        .O(\u0/out12 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5E92E56269D25879)) 
    g0_b1__96
       (.I0(\u0/u12/X [17]),
        .I1(\u0/u12/X [16]),
        .I2(\u0/u12/X [15]),
        .I3(\u0/u12/X [14]),
        .I4(\u0/u12/X [18]),
        .I5(\u0/u12/X [13]),
        .O(\u0/out12 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1BC6C996691BB46C)) 
    g0_b1__97
       (.I0(\u0/u12/X [35]),
        .I1(\u0/u12/X [34]),
        .I2(\u0/u12/X [33]),
        .I3(\u0/u12/X [32]),
        .I4(\u0/u12/X [36]),
        .I5(\u0/u12/X [31]),
        .O(\u0/out12 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h47B4E81E58B98679)) 
    g0_b1__98
       (.I0(\u0/u12/X [11]),
        .I1(\u0/u12/X [10]),
        .I2(\u0/u12/X [9]),
        .I3(\u0/u12/X [8]),
        .I4(\u0/u12/X [12]),
        .I5(\u0/u12/X [7]),
        .O(\u0/out12 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD12D36C3AC728D72)) 
    g0_b1__99
       (.I0(\u0/u12/X [47]),
        .I1(\u0/u12/X [46]),
        .I2(\u0/u12/X [45]),
        .I3(\u0/u12/X [44]),
        .I4(\u0/u12/X [48]),
        .I5(\u0/u12/X [43]),
        .O(\u0/out12 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2
       (.I0(\u0/u0/X [41]),
        .I1(\u0/u0/X [40]),
        .I2(\u0/u0/X [39]),
        .I3(\u0/u0/X [38]),
        .I4(\u0/u0/X [42]),
        .I5(\u0/u0/X [37]),
        .O(\u0/out0 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__0
       (.I0(\u0/u0/X [17]),
        .I1(\u0/u0/X [16]),
        .I2(\u0/u0/X [15]),
        .I3(\u0/u0/X [14]),
        .I4(\u0/u0/X [18]),
        .I5(\u0/u0/X [13]),
        .O(\u0/out0 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__1
       (.I0(\u0/u0/X [35]),
        .I1(\u0/u0/X [34]),
        .I2(\u0/u0/X [33]),
        .I3(\u0/u0/X [32]),
        .I4(\u0/u0/X [36]),
        .I5(\u0/u0/X [31]),
        .O(\u0/out0 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__10
       (.I0(\u0/u1/X [11]),
        .I1(\u0/u1/X [10]),
        .I2(\u0/u1/X [9]),
        .I3(\u0/u1/X [8]),
        .I4(\u0/u1/X [12]),
        .I5(\u0/u1/X [7]),
        .O(\u0/out1 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__100
       (.I0(\u0/u12/X [23]),
        .I1(\u0/u12/X [22]),
        .I2(\u0/u12/X [21]),
        .I3(\u0/u12/X [20]),
        .I4(\u0/u12/X [24]),
        .I5(\u0/u12/X [19]),
        .O(\u0/out12 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__101
       (.I0(\u0/u12/X [29]),
        .I1(\u0/u12/X [28]),
        .I2(\u0/u12/X [27]),
        .I3(\u0/u12/X [26]),
        .I4(\u0/u12/X [30]),
        .I5(\u0/u12/X [25]),
        .O(\u0/out12 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__102
       (.I0(\u0/u12/X [5]),
        .I1(\u0/u12/X [4]),
        .I2(\u0/u12/X [3]),
        .I3(\u0/u12/X [2]),
        .I4(\u0/u12/X [6]),
        .I5(\u0/u12/X [1]),
        .O(\u0/out12 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__103
       (.I0(\u0/u13/X [41]),
        .I1(\u0/u13/X [40]),
        .I2(\u0/u13/X [39]),
        .I3(\u0/u13/X [38]),
        .I4(\u0/u13/X [42]),
        .I5(\u0/u13/X [37]),
        .O(\u0/out13 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__104
       (.I0(\u0/u13/X [17]),
        .I1(\u0/u13/X [16]),
        .I2(\u0/u13/X [15]),
        .I3(\u0/u13/X [14]),
        .I4(\u0/u13/X [18]),
        .I5(\u0/u13/X [13]),
        .O(\u0/out13 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__105
       (.I0(\u0/u13/X [35]),
        .I1(\u0/u13/X [34]),
        .I2(\u0/u13/X [33]),
        .I3(\u0/u13/X [32]),
        .I4(\u0/u13/X [36]),
        .I5(\u0/u13/X [31]),
        .O(\u0/out13 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__106
       (.I0(\u0/u13/X [11]),
        .I1(\u0/u13/X [10]),
        .I2(\u0/u13/X [9]),
        .I3(\u0/u13/X [8]),
        .I4(\u0/u13/X [12]),
        .I5(\u0/u13/X [7]),
        .O(\u0/out13 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__107
       (.I0(\u0/u13/X [47]),
        .I1(\u0/u13/X [46]),
        .I2(\u0/u13/X [45]),
        .I3(\u0/u13/X [44]),
        .I4(\u0/u13/X [48]),
        .I5(\u0/u13/X [43]),
        .O(\u0/out13 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__108
       (.I0(\u0/u13/X [23]),
        .I1(\u0/u13/X [22]),
        .I2(\u0/u13/X [21]),
        .I3(\u0/u13/X [20]),
        .I4(\u0/u13/X [24]),
        .I5(\u0/u13/X [19]),
        .O(\u0/out13 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__109
       (.I0(\u0/u13/X [29]),
        .I1(\u0/u13/X [28]),
        .I2(\u0/u13/X [27]),
        .I3(\u0/u13/X [26]),
        .I4(\u0/u13/X [30]),
        .I5(\u0/u13/X [25]),
        .O(\u0/out13 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__11
       (.I0(\u0/u1/X [47]),
        .I1(\u0/u1/X [46]),
        .I2(\u0/u1/X [45]),
        .I3(\u0/u1/X [44]),
        .I4(\u0/u1/X [48]),
        .I5(\u0/u1/X [43]),
        .O(\u0/out1 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__110
       (.I0(\u0/u13/X [5]),
        .I1(\u0/u13/X [4]),
        .I2(\u0/u13/X [3]),
        .I3(\u0/u13/X [2]),
        .I4(\u0/u13/X [6]),
        .I5(\u0/u13/X [1]),
        .O(\u0/out13 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__111
       (.I0(\u0/u14/X [41]),
        .I1(\u0/u14/X [40]),
        .I2(\u0/u14/X [39]),
        .I3(\u0/u14/X [38]),
        .I4(\u0/u14/X [42]),
        .I5(\u0/u14/X [37]),
        .O(\u0/out14 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__112
       (.I0(\u0/u14/X [17]),
        .I1(\u0/u14/X [16]),
        .I2(\u0/u14/X [15]),
        .I3(\u0/u14/X [14]),
        .I4(\u0/u14/X [18]),
        .I5(\u0/u14/X [13]),
        .O(\u0/out14 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__113
       (.I0(\u0/u14/X [35]),
        .I1(\u0/u14/X [34]),
        .I2(\u0/u14/X [33]),
        .I3(\u0/u14/X [32]),
        .I4(\u0/u14/X [36]),
        .I5(\u0/u14/X [31]),
        .O(\u0/out14 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__114
       (.I0(\u0/u14/X [11]),
        .I1(\u0/u14/X [10]),
        .I2(\u0/u14/X [9]),
        .I3(\u0/u14/X [8]),
        .I4(\u0/u14/X [12]),
        .I5(\u0/u14/X [7]),
        .O(\u0/out14 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__115
       (.I0(\u0/u14/X [47]),
        .I1(\u0/u14/X [46]),
        .I2(\u0/u14/X [45]),
        .I3(\u0/u14/X [44]),
        .I4(\u0/u14/X [48]),
        .I5(\u0/u14/X [43]),
        .O(\u0/out14 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__116
       (.I0(\u0/u14/X [23]),
        .I1(\u0/u14/X [22]),
        .I2(\u0/u14/X [21]),
        .I3(\u0/u14/X [20]),
        .I4(\u0/u14/X [24]),
        .I5(\u0/u14/X [19]),
        .O(\u0/out14 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__117
       (.I0(\u0/u14/X [29]),
        .I1(\u0/u14/X [28]),
        .I2(\u0/u14/X [27]),
        .I3(\u0/u14/X [26]),
        .I4(\u0/u14/X [30]),
        .I5(\u0/u14/X [25]),
        .O(\u0/out14 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__118
       (.I0(\u0/u14/X [5]),
        .I1(\u0/u14/X [4]),
        .I2(\u0/u14/X [3]),
        .I3(\u0/u14/X [2]),
        .I4(\u0/u14/X [6]),
        .I5(\u0/u14/X [1]),
        .O(\u0/out14 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__119
       (.I0(\u0/u15/X [41]),
        .I1(\u0/u15/X [40]),
        .I2(\u0/u15/X [39]),
        .I3(\u0/u15/X [38]),
        .I4(\u0/u15/X [42]),
        .I5(\u0/u15/X [37]),
        .O(\u0/out15 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__12
       (.I0(\u0/u1/X [23]),
        .I1(\u0/u1/X [22]),
        .I2(\u0/u1/X [21]),
        .I3(\u0/u1/X [20]),
        .I4(\u0/u1/X [24]),
        .I5(\u0/u1/X [19]),
        .O(\u0/out1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__120
       (.I0(\u0/u15/X [17]),
        .I1(\u0/u15/X [16]),
        .I2(\u0/u15/X [15]),
        .I3(\u0/u15/X [14]),
        .I4(\u0/u15/X [18]),
        .I5(\u0/u15/X [13]),
        .O(\u0/out15 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__121
       (.I0(\u0/u15/X [35]),
        .I1(\u0/u15/X [34]),
        .I2(\u0/u15/X [33]),
        .I3(\u0/u15/X [32]),
        .I4(\u0/u15/X [36]),
        .I5(\u0/u15/X [31]),
        .O(\u0/out15 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__122
       (.I0(\u0/u15/X [11]),
        .I1(\u0/u15/X [10]),
        .I2(\u0/u15/X [9]),
        .I3(\u0/u15/X [8]),
        .I4(\u0/u15/X [12]),
        .I5(\u0/u15/X [7]),
        .O(\u0/out15 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__123
       (.I0(\u0/u15/X [47]),
        .I1(\u0/u15/X [46]),
        .I2(\u0/u15/X [45]),
        .I3(\u0/u15/X [44]),
        .I4(\u0/u15/X [48]),
        .I5(\u0/u15/X [43]),
        .O(\u0/out15 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__124
       (.I0(\u0/u15/X [23]),
        .I1(\u0/u15/X [22]),
        .I2(\u0/u15/X [21]),
        .I3(\u0/u15/X [20]),
        .I4(\u0/u15/X [24]),
        .I5(\u0/u15/X [19]),
        .O(\u0/out15 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__125
       (.I0(\u0/u15/X [29]),
        .I1(\u0/u15/X [28]),
        .I2(\u0/u15/X [27]),
        .I3(\u0/u15/X [26]),
        .I4(\u0/u15/X [30]),
        .I5(\u0/u15/X [25]),
        .O(\u0/out15 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__126
       (.I0(\u0/u15/X [5]),
        .I1(\u0/u15/X [4]),
        .I2(\u0/u15/X [3]),
        .I3(\u0/u15/X [2]),
        .I4(\u0/u15/X [6]),
        .I5(\u0/u15/X [1]),
        .O(\u0/out15 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__127
       (.I0(\u1/u0/X [41]),
        .I1(\u1/u0/X [40]),
        .I2(\u1/u0/X [39]),
        .I3(\u1/u0/X [38]),
        .I4(\u1/u0/X [42]),
        .I5(\u1/u0/X [37]),
        .O(\u1/out0 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__128
       (.I0(\u1/u0/X [17]),
        .I1(\u1/u0/X [16]),
        .I2(\u1/u0/X [15]),
        .I3(\u1/u0/X [14]),
        .I4(\u1/u0/X [18]),
        .I5(\u1/u0/X [13]),
        .O(\u1/out0 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__129
       (.I0(\u1/u0/X [35]),
        .I1(\u1/u0/X [34]),
        .I2(\u1/u0/X [33]),
        .I3(\u1/u0/X [32]),
        .I4(\u1/u0/X [36]),
        .I5(\u1/u0/X [31]),
        .O(\u1/out0 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__13
       (.I0(\u0/u1/X [29]),
        .I1(\u0/u1/X [28]),
        .I2(\u0/u1/X [27]),
        .I3(\u0/u1/X [26]),
        .I4(\u0/u1/X [30]),
        .I5(\u0/u1/X [25]),
        .O(\u0/out1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__130
       (.I0(\u1/u0/X [11]),
        .I1(\u1/u0/X [10]),
        .I2(\u1/u0/X [9]),
        .I3(\u1/u0/X [8]),
        .I4(\u1/u0/X [12]),
        .I5(\u1/u0/X [7]),
        .O(\u1/out0 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__131
       (.I0(\u1/u0/X [47]),
        .I1(\u1/u0/X [46]),
        .I2(\u1/u0/X [45]),
        .I3(\u1/u0/X [44]),
        .I4(\u1/u0/X [48]),
        .I5(\u1/u0/X [43]),
        .O(\u1/out0 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__132
       (.I0(\u1/u0/X [23]),
        .I1(\u1/u0/X [22]),
        .I2(\u1/u0/X [21]),
        .I3(\u1/u0/X [20]),
        .I4(\u1/u0/X [24]),
        .I5(\u1/u0/X [19]),
        .O(\u1/out0 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__133
       (.I0(\u1/u0/X [29]),
        .I1(\u1/u0/X [28]),
        .I2(\u1/u0/X [27]),
        .I3(\u1/u0/X [26]),
        .I4(\u1/u0/X [30]),
        .I5(\u1/u0/X [25]),
        .O(\u1/out0 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__134
       (.I0(\u1/u0/X [5]),
        .I1(\u1/u0/X [4]),
        .I2(\u1/u0/X [3]),
        .I3(\u1/u0/X [2]),
        .I4(\u1/u0/X [6]),
        .I5(\u1/u0/X [1]),
        .O(\u1/out0 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__135
       (.I0(\u1/u1/X [41]),
        .I1(\u1/u1/X [40]),
        .I2(\u1/u1/X [39]),
        .I3(\u1/u1/X [38]),
        .I4(\u1/u1/X [42]),
        .I5(\u1/u1/X [37]),
        .O(\u1/out1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__136
       (.I0(\u1/u1/X [17]),
        .I1(\u1/u1/X [16]),
        .I2(\u1/u1/X [15]),
        .I3(\u1/u1/X [14]),
        .I4(\u1/u1/X [18]),
        .I5(\u1/u1/X [13]),
        .O(\u1/out1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__137
       (.I0(\u1/u1/X [35]),
        .I1(\u1/u1/X [34]),
        .I2(\u1/u1/X [33]),
        .I3(\u1/u1/X [32]),
        .I4(\u1/u1/X [36]),
        .I5(\u1/u1/X [31]),
        .O(\u1/out1 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__138
       (.I0(\u1/u1/X [11]),
        .I1(\u1/u1/X [10]),
        .I2(\u1/u1/X [9]),
        .I3(\u1/u1/X [8]),
        .I4(\u1/u1/X [12]),
        .I5(\u1/u1/X [7]),
        .O(\u1/out1 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__139
       (.I0(\u1/u1/X [47]),
        .I1(\u1/u1/X [46]),
        .I2(\u1/u1/X [45]),
        .I3(\u1/u1/X [44]),
        .I4(\u1/u1/X [48]),
        .I5(\u1/u1/X [43]),
        .O(\u1/out1 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__14
       (.I0(\u0/u1/X [5]),
        .I1(\u0/u1/X [4]),
        .I2(\u0/u1/X [3]),
        .I3(\u0/u1/X [2]),
        .I4(\u0/u1/X [6]),
        .I5(\u0/u1/X [1]),
        .O(\u0/out1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__140
       (.I0(\u1/u1/X [23]),
        .I1(\u1/u1/X [22]),
        .I2(\u1/u1/X [21]),
        .I3(\u1/u1/X [20]),
        .I4(\u1/u1/X [24]),
        .I5(\u1/u1/X [19]),
        .O(\u1/out1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__141
       (.I0(\u1/u1/X [29]),
        .I1(\u1/u1/X [28]),
        .I2(\u1/u1/X [27]),
        .I3(\u1/u1/X [26]),
        .I4(\u1/u1/X [30]),
        .I5(\u1/u1/X [25]),
        .O(\u1/out1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__142
       (.I0(\u1/u1/X [5]),
        .I1(\u1/u1/X [4]),
        .I2(\u1/u1/X [3]),
        .I3(\u1/u1/X [2]),
        .I4(\u1/u1/X [6]),
        .I5(\u1/u1/X [1]),
        .O(\u1/out1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__143
       (.I0(\u1/u2/X [41]),
        .I1(\u1/u2/X [40]),
        .I2(\u1/u2/X [39]),
        .I3(\u1/u2/X [38]),
        .I4(\u1/u2/X [42]),
        .I5(\u1/u2/X [37]),
        .O(\u1/out2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__144
       (.I0(\u1/u2/X [17]),
        .I1(\u1/u2/X [16]),
        .I2(\u1/u2/X [15]),
        .I3(\u1/u2/X [14]),
        .I4(\u1/u2/X [18]),
        .I5(\u1/u2/X [13]),
        .O(\u1/out2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__145
       (.I0(\u1/u2/X [35]),
        .I1(\u1/u2/X [34]),
        .I2(\u1/u2/X [33]),
        .I3(\u1/u2/X [32]),
        .I4(\u1/u2/X [36]),
        .I5(\u1/u2/X [31]),
        .O(\u1/out2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__146
       (.I0(\u1/u2/X [11]),
        .I1(\u1/u2/X [10]),
        .I2(\u1/u2/X [9]),
        .I3(\u1/u2/X [8]),
        .I4(\u1/u2/X [12]),
        .I5(\u1/u2/X [7]),
        .O(\u1/out2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__147
       (.I0(\u1/u2/X [47]),
        .I1(\u1/u2/X [46]),
        .I2(\u1/u2/X [45]),
        .I3(\u1/u2/X [44]),
        .I4(\u1/u2/X [48]),
        .I5(\u1/u2/X [43]),
        .O(\u1/out2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__148
       (.I0(\u1/u2/X [23]),
        .I1(\u1/u2/X [22]),
        .I2(\u1/u2/X [21]),
        .I3(\u1/u2/X [20]),
        .I4(\u1/u2/X [24]),
        .I5(\u1/u2/X [19]),
        .O(\u1/out2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__149
       (.I0(\u1/u2/X [29]),
        .I1(\u1/u2/X [28]),
        .I2(\u1/u2/X [27]),
        .I3(\u1/u2/X [26]),
        .I4(\u1/u2/X [30]),
        .I5(\u1/u2/X [25]),
        .O(\u1/out2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__15
       (.I0(\u0/u2/X [41]),
        .I1(\u0/u2/X [40]),
        .I2(\u0/u2/X [39]),
        .I3(\u0/u2/X [38]),
        .I4(\u0/u2/X [42]),
        .I5(\u0/u2/X [37]),
        .O(\u0/out2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__150
       (.I0(\u1/u2/X [5]),
        .I1(\u1/u2/X [4]),
        .I2(\u1/u2/X [3]),
        .I3(\u1/u2/X [2]),
        .I4(\u1/u2/X [6]),
        .I5(\u1/u2/X [1]),
        .O(\u1/out2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__151
       (.I0(\u1/u3/X [41]),
        .I1(\u1/u3/X [40]),
        .I2(\u1/u3/X [39]),
        .I3(\u1/u3/X [38]),
        .I4(\u1/u3/X [42]),
        .I5(\u1/u3/X [37]),
        .O(\u1/out3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__152
       (.I0(\u1/u3/X [17]),
        .I1(\u1/u3/X [16]),
        .I2(\u1/u3/X [15]),
        .I3(\u1/u3/X [14]),
        .I4(\u1/u3/X [18]),
        .I5(\u1/u3/X [13]),
        .O(\u1/out3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__153
       (.I0(\u1/u3/X [35]),
        .I1(\u1/u3/X [34]),
        .I2(\u1/u3/X [33]),
        .I3(\u1/u3/X [32]),
        .I4(\u1/u3/X [36]),
        .I5(\u1/u3/X [31]),
        .O(\u1/out3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__154
       (.I0(\u1/u3/X [11]),
        .I1(\u1/u3/X [10]),
        .I2(\u1/u3/X [9]),
        .I3(\u1/u3/X [8]),
        .I4(\u1/u3/X [12]),
        .I5(\u1/u3/X [7]),
        .O(\u1/out3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__155
       (.I0(\u1/u3/X [47]),
        .I1(\u1/u3/X [46]),
        .I2(\u1/u3/X [45]),
        .I3(\u1/u3/X [44]),
        .I4(\u1/u3/X [48]),
        .I5(\u1/u3/X [43]),
        .O(\u1/out3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__156
       (.I0(\u1/u3/X [23]),
        .I1(\u1/u3/X [22]),
        .I2(\u1/u3/X [21]),
        .I3(\u1/u3/X [20]),
        .I4(\u1/u3/X [24]),
        .I5(\u1/u3/X [19]),
        .O(\u1/out3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__157
       (.I0(\u1/u3/X [29]),
        .I1(\u1/u3/X [28]),
        .I2(\u1/u3/X [27]),
        .I3(\u1/u3/X [26]),
        .I4(\u1/u3/X [30]),
        .I5(\u1/u3/X [25]),
        .O(\u1/out3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__158
       (.I0(\u1/u3/X [5]),
        .I1(\u1/u3/X [4]),
        .I2(\u1/u3/X [3]),
        .I3(\u1/u3/X [2]),
        .I4(\u1/u3/X [6]),
        .I5(\u1/u3/X [1]),
        .O(\u1/out3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__159
       (.I0(\u1/u4/X [41]),
        .I1(\u1/u4/X [40]),
        .I2(\u1/u4/X [39]),
        .I3(\u1/u4/X [38]),
        .I4(\u1/u4/X [42]),
        .I5(\u1/u4/X [37]),
        .O(\u1/out4 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__16
       (.I0(\u0/u2/X [17]),
        .I1(\u0/u2/X [16]),
        .I2(\u0/u2/X [15]),
        .I3(\u0/u2/X [14]),
        .I4(\u0/u2/X [18]),
        .I5(\u0/u2/X [13]),
        .O(\u0/out2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__160
       (.I0(\u1/u4/X [17]),
        .I1(\u1/u4/X [16]),
        .I2(\u1/u4/X [15]),
        .I3(\u1/u4/X [14]),
        .I4(\u1/u4/X [18]),
        .I5(\u1/u4/X [13]),
        .O(\u1/out4 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__161
       (.I0(\u1/u4/X [35]),
        .I1(\u1/u4/X [34]),
        .I2(\u1/u4/X [33]),
        .I3(\u1/u4/X [32]),
        .I4(\u1/u4/X [36]),
        .I5(\u1/u4/X [31]),
        .O(\u1/out4 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__162
       (.I0(\u1/u4/X [11]),
        .I1(\u1/u4/X [10]),
        .I2(\u1/u4/X [9]),
        .I3(\u1/u4/X [8]),
        .I4(\u1/u4/X [12]),
        .I5(\u1/u4/X [7]),
        .O(\u1/out4 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__163
       (.I0(\u1/u4/X [47]),
        .I1(\u1/u4/X [46]),
        .I2(\u1/u4/X [45]),
        .I3(\u1/u4/X [44]),
        .I4(\u1/u4/X [48]),
        .I5(\u1/u4/X [43]),
        .O(\u1/out4 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__164
       (.I0(\u1/u4/X [23]),
        .I1(\u1/u4/X [22]),
        .I2(\u1/u4/X [21]),
        .I3(\u1/u4/X [20]),
        .I4(\u1/u4/X [24]),
        .I5(\u1/u4/X [19]),
        .O(\u1/out4 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__165
       (.I0(\u1/u4/X [29]),
        .I1(\u1/u4/X [28]),
        .I2(\u1/u4/X [27]),
        .I3(\u1/u4/X [26]),
        .I4(\u1/u4/X [30]),
        .I5(\u1/u4/X [25]),
        .O(\u1/out4 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__166
       (.I0(\u1/u4/X [5]),
        .I1(\u1/u4/X [4]),
        .I2(\u1/u4/X [3]),
        .I3(\u1/u4/X [2]),
        .I4(\u1/u4/X [6]),
        .I5(\u1/u4/X [1]),
        .O(\u1/out4 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__167
       (.I0(\u1/u5/X [41]),
        .I1(\u1/u5/X [40]),
        .I2(\u1/u5/X [39]),
        .I3(\u1/u5/X [38]),
        .I4(\u1/u5/X [42]),
        .I5(\u1/u5/X [37]),
        .O(\u1/out5 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__168
       (.I0(\u1/u5/X [17]),
        .I1(\u1/u5/X [16]),
        .I2(\u1/u5/X [15]),
        .I3(\u1/u5/X [14]),
        .I4(\u1/u5/X [18]),
        .I5(\u1/u5/X [13]),
        .O(\u1/out5 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__169
       (.I0(\u1/u5/X [35]),
        .I1(\u1/u5/X [34]),
        .I2(\u1/u5/X [33]),
        .I3(\u1/u5/X [32]),
        .I4(\u1/u5/X [36]),
        .I5(\u1/u5/X [31]),
        .O(\u1/out5 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__17
       (.I0(\u0/u2/X [35]),
        .I1(\u0/u2/X [34]),
        .I2(\u0/u2/X [33]),
        .I3(\u0/u2/X [32]),
        .I4(\u0/u2/X [36]),
        .I5(\u0/u2/X [31]),
        .O(\u0/out2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__170
       (.I0(\u1/u5/X [11]),
        .I1(\u1/u5/X [10]),
        .I2(\u1/u5/X [9]),
        .I3(\u1/u5/X [8]),
        .I4(\u1/u5/X [12]),
        .I5(\u1/u5/X [7]),
        .O(\u1/out5 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__171
       (.I0(\u1/u5/X [47]),
        .I1(\u1/u5/X [46]),
        .I2(\u1/u5/X [45]),
        .I3(\u1/u5/X [44]),
        .I4(\u1/u5/X [48]),
        .I5(\u1/u5/X [43]),
        .O(\u1/out5 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__172
       (.I0(\u1/u5/X [23]),
        .I1(\u1/u5/X [22]),
        .I2(\u1/u5/X [21]),
        .I3(\u1/u5/X [20]),
        .I4(\u1/u5/X [24]),
        .I5(\u1/u5/X [19]),
        .O(\u1/out5 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__173
       (.I0(\u1/u5/X [29]),
        .I1(\u1/u5/X [28]),
        .I2(\u1/u5/X [27]),
        .I3(\u1/u5/X [26]),
        .I4(\u1/u5/X [30]),
        .I5(\u1/u5/X [25]),
        .O(\u1/out5 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__174
       (.I0(\u1/u5/X [5]),
        .I1(\u1/u5/X [4]),
        .I2(\u1/u5/X [3]),
        .I3(\u1/u5/X [2]),
        .I4(\u1/u5/X [6]),
        .I5(\u1/u5/X [1]),
        .O(\u1/out5 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__175
       (.I0(\u1/u6/X [41]),
        .I1(\u1/u6/X [40]),
        .I2(\u1/u6/X [39]),
        .I3(\u1/u6/X [38]),
        .I4(\u1/u6/X [42]),
        .I5(\u1/u6/X [37]),
        .O(\u1/out6 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__176
       (.I0(\u1/u6/X [17]),
        .I1(\u1/u6/X [16]),
        .I2(\u1/u6/X [15]),
        .I3(\u1/u6/X [14]),
        .I4(\u1/u6/X [18]),
        .I5(\u1/u6/X [13]),
        .O(\u1/out6 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__177
       (.I0(\u1/u6/X [35]),
        .I1(\u1/u6/X [34]),
        .I2(\u1/u6/X [33]),
        .I3(\u1/u6/X [32]),
        .I4(\u1/u6/X [36]),
        .I5(\u1/u6/X [31]),
        .O(\u1/out6 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__178
       (.I0(\u1/u6/X [11]),
        .I1(\u1/u6/X [10]),
        .I2(\u1/u6/X [9]),
        .I3(\u1/u6/X [8]),
        .I4(\u1/u6/X [12]),
        .I5(\u1/u6/X [7]),
        .O(\u1/out6 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__179
       (.I0(\u1/u6/X [47]),
        .I1(\u1/u6/X [46]),
        .I2(\u1/u6/X [45]),
        .I3(\u1/u6/X [44]),
        .I4(\u1/u6/X [48]),
        .I5(\u1/u6/X [43]),
        .O(\u1/out6 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__18
       (.I0(\u0/u2/X [11]),
        .I1(\u0/u2/X [10]),
        .I2(\u0/u2/X [9]),
        .I3(\u0/u2/X [8]),
        .I4(\u0/u2/X [12]),
        .I5(\u0/u2/X [7]),
        .O(\u0/out2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__180
       (.I0(\u1/u6/X [23]),
        .I1(\u1/u6/X [22]),
        .I2(\u1/u6/X [21]),
        .I3(\u1/u6/X [20]),
        .I4(\u1/u6/X [24]),
        .I5(\u1/u6/X [19]),
        .O(\u1/out6 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__181
       (.I0(\u1/u6/X [29]),
        .I1(\u1/u6/X [28]),
        .I2(\u1/u6/X [27]),
        .I3(\u1/u6/X [26]),
        .I4(\u1/u6/X [30]),
        .I5(\u1/u6/X [25]),
        .O(\u1/out6 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__182
       (.I0(\u1/u6/X [5]),
        .I1(\u1/u6/X [4]),
        .I2(\u1/u6/X [3]),
        .I3(\u1/u6/X [2]),
        .I4(\u1/u6/X [6]),
        .I5(\u1/u6/X [1]),
        .O(\u1/out6 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__183
       (.I0(\u1/u7/X [41]),
        .I1(\u1/u7/X [40]),
        .I2(\u1/u7/X [39]),
        .I3(\u1/u7/X [38]),
        .I4(\u1/u7/X [42]),
        .I5(\u1/u7/X [37]),
        .O(\u1/out7 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__184
       (.I0(\u1/u7/X [17]),
        .I1(\u1/u7/X [16]),
        .I2(\u1/u7/X [15]),
        .I3(\u1/u7/X [14]),
        .I4(\u1/u7/X [18]),
        .I5(\u1/u7/X [13]),
        .O(\u1/out7 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__185
       (.I0(\u1/u7/X [35]),
        .I1(\u1/u7/X [34]),
        .I2(\u1/u7/X [33]),
        .I3(\u1/u7/X [32]),
        .I4(\u1/u7/X [36]),
        .I5(\u1/u7/X [31]),
        .O(\u1/out7 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__186
       (.I0(\u1/u7/X [11]),
        .I1(\u1/u7/X [10]),
        .I2(\u1/u7/X [9]),
        .I3(\u1/u7/X [8]),
        .I4(\u1/u7/X [12]),
        .I5(\u1/u7/X [7]),
        .O(\u1/out7 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__187
       (.I0(\u1/u7/X [47]),
        .I1(\u1/u7/X [46]),
        .I2(\u1/u7/X [45]),
        .I3(\u1/u7/X [44]),
        .I4(\u1/u7/X [48]),
        .I5(\u1/u7/X [43]),
        .O(\u1/out7 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__188
       (.I0(\u1/u7/X [23]),
        .I1(\u1/u7/X [22]),
        .I2(\u1/u7/X [21]),
        .I3(\u1/u7/X [20]),
        .I4(\u1/u7/X [24]),
        .I5(\u1/u7/X [19]),
        .O(\u1/out7 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__189
       (.I0(\u1/u7/X [29]),
        .I1(\u1/u7/X [28]),
        .I2(\u1/u7/X [27]),
        .I3(\u1/u7/X [26]),
        .I4(\u1/u7/X [30]),
        .I5(\u1/u7/X [25]),
        .O(\u1/out7 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__19
       (.I0(\u0/u2/X [47]),
        .I1(\u0/u2/X [46]),
        .I2(\u0/u2/X [45]),
        .I3(\u0/u2/X [44]),
        .I4(\u0/u2/X [48]),
        .I5(\u0/u2/X [43]),
        .O(\u0/out2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__190
       (.I0(\u1/u7/X [5]),
        .I1(\u1/u7/X [4]),
        .I2(\u1/u7/X [3]),
        .I3(\u1/u7/X [2]),
        .I4(\u1/u7/X [6]),
        .I5(\u1/u7/X [1]),
        .O(\u1/out7 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__191
       (.I0(\u1/u8/X [41]),
        .I1(\u1/u8/X [40]),
        .I2(\u1/u8/X [39]),
        .I3(\u1/u8/X [38]),
        .I4(\u1/u8/X [42]),
        .I5(\u1/u8/X [37]),
        .O(\u1/out8 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__192
       (.I0(\u1/u8/X [17]),
        .I1(\u1/u8/X [16]),
        .I2(\u1/u8/X [15]),
        .I3(\u1/u8/X [14]),
        .I4(\u1/u8/X [18]),
        .I5(\u1/u8/X [13]),
        .O(\u1/out8 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__193
       (.I0(\u1/u8/X [35]),
        .I1(\u1/u8/X [34]),
        .I2(\u1/u8/X [33]),
        .I3(\u1/u8/X [32]),
        .I4(\u1/u8/X [36]),
        .I5(\u1/u8/X [31]),
        .O(\u1/out8 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__194
       (.I0(\u1/u8/X [11]),
        .I1(\u1/u8/X [10]),
        .I2(\u1/u8/X [9]),
        .I3(\u1/u8/X [8]),
        .I4(\u1/u8/X [12]),
        .I5(\u1/u8/X [7]),
        .O(\u1/out8 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__195
       (.I0(\u1/u8/X [47]),
        .I1(\u1/u8/X [46]),
        .I2(\u1/u8/X [45]),
        .I3(\u1/u8/X [44]),
        .I4(\u1/u8/X [48]),
        .I5(\u1/u8/X [43]),
        .O(\u1/out8 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__196
       (.I0(\u1/u8/X [23]),
        .I1(\u1/u8/X [22]),
        .I2(\u1/u8/X [21]),
        .I3(\u1/u8/X [20]),
        .I4(\u1/u8/X [24]),
        .I5(\u1/u8/X [19]),
        .O(\u1/out8 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__197
       (.I0(\u1/u8/X [29]),
        .I1(\u1/u8/X [28]),
        .I2(\u1/u8/X [27]),
        .I3(\u1/u8/X [26]),
        .I4(\u1/u8/X [30]),
        .I5(\u1/u8/X [25]),
        .O(\u1/out8 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__198
       (.I0(\u1/u8/X [5]),
        .I1(\u1/u8/X [4]),
        .I2(\u1/u8/X [3]),
        .I3(\u1/u8/X [2]),
        .I4(\u1/u8/X [6]),
        .I5(\u1/u8/X [1]),
        .O(\u1/out8 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__199
       (.I0(\u1/u9/X [41]),
        .I1(\u1/u9/X [40]),
        .I2(\u1/u9/X [39]),
        .I3(\u1/u9/X [38]),
        .I4(\u1/u9/X [42]),
        .I5(\u1/u9/X [37]),
        .O(\u1/out9 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__2
       (.I0(\u0/u0/X [11]),
        .I1(\u0/u0/X [10]),
        .I2(\u0/u0/X [9]),
        .I3(\u0/u0/X [8]),
        .I4(\u0/u0/X [12]),
        .I5(\u0/u0/X [7]),
        .O(\u0/out0 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__20
       (.I0(\u0/u2/X [23]),
        .I1(\u0/u2/X [22]),
        .I2(\u0/u2/X [21]),
        .I3(\u0/u2/X [20]),
        .I4(\u0/u2/X [24]),
        .I5(\u0/u2/X [19]),
        .O(\u0/out2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__200
       (.I0(\u1/u9/X [17]),
        .I1(\u1/u9/X [16]),
        .I2(\u1/u9/X [15]),
        .I3(\u1/u9/X [14]),
        .I4(\u1/u9/X [18]),
        .I5(\u1/u9/X [13]),
        .O(\u1/out9 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__201
       (.I0(\u1/u9/X [35]),
        .I1(\u1/u9/X [34]),
        .I2(\u1/u9/X [33]),
        .I3(\u1/u9/X [32]),
        .I4(\u1/u9/X [36]),
        .I5(\u1/u9/X [31]),
        .O(\u1/out9 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__202
       (.I0(\u1/u9/X [11]),
        .I1(\u1/u9/X [10]),
        .I2(\u1/u9/X [9]),
        .I3(\u1/u9/X [8]),
        .I4(\u1/u9/X [12]),
        .I5(\u1/u9/X [7]),
        .O(\u1/out9 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__203
       (.I0(\u1/u9/X [47]),
        .I1(\u1/u9/X [46]),
        .I2(\u1/u9/X [45]),
        .I3(\u1/u9/X [44]),
        .I4(\u1/u9/X [48]),
        .I5(\u1/u9/X [43]),
        .O(\u1/out9 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__204
       (.I0(\u1/u9/X [23]),
        .I1(\u1/u9/X [22]),
        .I2(\u1/u9/X [21]),
        .I3(\u1/u9/X [20]),
        .I4(\u1/u9/X [24]),
        .I5(\u1/u9/X [19]),
        .O(\u1/out9 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__205
       (.I0(\u1/u9/X [29]),
        .I1(\u1/u9/X [28]),
        .I2(\u1/u9/X [27]),
        .I3(\u1/u9/X [26]),
        .I4(\u1/u9/X [30]),
        .I5(\u1/u9/X [25]),
        .O(\u1/out9 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__206
       (.I0(\u1/u9/X [5]),
        .I1(\u1/u9/X [4]),
        .I2(\u1/u9/X [3]),
        .I3(\u1/u9/X [2]),
        .I4(\u1/u9/X [6]),
        .I5(\u1/u9/X [1]),
        .O(\u1/out9 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__207
       (.I0(\u1/u10/X [41]),
        .I1(\u1/u10/X [40]),
        .I2(\u1/u10/X [39]),
        .I3(\u1/u10/X [38]),
        .I4(\u1/u10/X [42]),
        .I5(\u1/u10/X [37]),
        .O(\u1/out10 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__208
       (.I0(\u1/u10/X [17]),
        .I1(\u1/u10/X [16]),
        .I2(\u1/u10/X [15]),
        .I3(\u1/u10/X [14]),
        .I4(\u1/u10/X [18]),
        .I5(\u1/u10/X [13]),
        .O(\u1/out10 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__209
       (.I0(\u1/u10/X [35]),
        .I1(\u1/u10/X [34]),
        .I2(\u1/u10/X [33]),
        .I3(\u1/u10/X [32]),
        .I4(\u1/u10/X [36]),
        .I5(\u1/u10/X [31]),
        .O(\u1/out10 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__21
       (.I0(\u0/u2/X [29]),
        .I1(\u0/u2/X [28]),
        .I2(\u0/u2/X [27]),
        .I3(\u0/u2/X [26]),
        .I4(\u0/u2/X [30]),
        .I5(\u0/u2/X [25]),
        .O(\u0/out2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__210
       (.I0(\u1/u10/X [11]),
        .I1(\u1/u10/X [10]),
        .I2(\u1/u10/X [9]),
        .I3(\u1/u10/X [8]),
        .I4(\u1/u10/X [12]),
        .I5(\u1/u10/X [7]),
        .O(\u1/out10 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__211
       (.I0(\u1/u10/X [47]),
        .I1(\u1/u10/X [46]),
        .I2(\u1/u10/X [45]),
        .I3(\u1/u10/X [44]),
        .I4(\u1/u10/X [48]),
        .I5(\u1/u10/X [43]),
        .O(\u1/out10 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__212
       (.I0(\u1/u10/X [23]),
        .I1(\u1/u10/X [22]),
        .I2(\u1/u10/X [21]),
        .I3(\u1/u10/X [20]),
        .I4(\u1/u10/X [24]),
        .I5(\u1/u10/X [19]),
        .O(\u1/out10 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__213
       (.I0(\u1/u10/X [29]),
        .I1(\u1/u10/X [28]),
        .I2(\u1/u10/X [27]),
        .I3(\u1/u10/X [26]),
        .I4(\u1/u10/X [30]),
        .I5(\u1/u10/X [25]),
        .O(\u1/out10 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__214
       (.I0(\u1/u10/X [5]),
        .I1(\u1/u10/X [4]),
        .I2(\u1/u10/X [3]),
        .I3(\u1/u10/X [2]),
        .I4(\u1/u10/X [6]),
        .I5(\u1/u10/X [1]),
        .O(\u1/out10 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__215
       (.I0(\u1/u11/X [41]),
        .I1(\u1/u11/X [40]),
        .I2(\u1/u11/X [39]),
        .I3(\u1/u11/X [38]),
        .I4(\u1/u11/X [42]),
        .I5(\u1/u11/X [37]),
        .O(\u1/out11 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__216
       (.I0(\u1/u11/X [17]),
        .I1(\u1/u11/X [16]),
        .I2(\u1/u11/X [15]),
        .I3(\u1/u11/X [14]),
        .I4(\u1/u11/X [18]),
        .I5(\u1/u11/X [13]),
        .O(\u1/out11 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__217
       (.I0(\u1/u11/X [35]),
        .I1(\u1/u11/X [34]),
        .I2(\u1/u11/X [33]),
        .I3(\u1/u11/X [32]),
        .I4(\u1/u11/X [36]),
        .I5(\u1/u11/X [31]),
        .O(\u1/out11 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__218
       (.I0(\u1/u11/X [11]),
        .I1(\u1/u11/X [10]),
        .I2(\u1/u11/X [9]),
        .I3(\u1/u11/X [8]),
        .I4(\u1/u11/X [12]),
        .I5(\u1/u11/X [7]),
        .O(\u1/out11 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__219
       (.I0(\u1/u11/X [47]),
        .I1(\u1/u11/X [46]),
        .I2(\u1/u11/X [45]),
        .I3(\u1/u11/X [44]),
        .I4(\u1/u11/X [48]),
        .I5(\u1/u11/X [43]),
        .O(\u1/out11 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__22
       (.I0(\u0/u2/X [5]),
        .I1(\u0/u2/X [4]),
        .I2(\u0/u2/X [3]),
        .I3(\u0/u2/X [2]),
        .I4(\u0/u2/X [6]),
        .I5(\u0/u2/X [1]),
        .O(\u0/out2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__220
       (.I0(\u1/u11/X [23]),
        .I1(\u1/u11/X [22]),
        .I2(\u1/u11/X [21]),
        .I3(\u1/u11/X [20]),
        .I4(\u1/u11/X [24]),
        .I5(\u1/u11/X [19]),
        .O(\u1/out11 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__221
       (.I0(\u1/u11/X [29]),
        .I1(\u1/u11/X [28]),
        .I2(\u1/u11/X [27]),
        .I3(\u1/u11/X [26]),
        .I4(\u1/u11/X [30]),
        .I5(\u1/u11/X [25]),
        .O(\u1/out11 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__222
       (.I0(\u1/u11/X [5]),
        .I1(\u1/u11/X [4]),
        .I2(\u1/u11/X [3]),
        .I3(\u1/u11/X [2]),
        .I4(\u1/u11/X [6]),
        .I5(\u1/u11/X [1]),
        .O(\u1/out11 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__223
       (.I0(\u1/u12/X [41]),
        .I1(\u1/u12/X [40]),
        .I2(\u1/u12/X [39]),
        .I3(\u1/u12/X [38]),
        .I4(\u1/u12/X [42]),
        .I5(\u1/u12/X [37]),
        .O(\u1/out12 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__224
       (.I0(\u1/u12/X [17]),
        .I1(\u1/u12/X [16]),
        .I2(\u1/u12/X [15]),
        .I3(\u1/u12/X [14]),
        .I4(\u1/u12/X [18]),
        .I5(\u1/u12/X [13]),
        .O(\u1/out12 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__225
       (.I0(\u1/u12/X [35]),
        .I1(\u1/u12/X [34]),
        .I2(\u1/u12/X [33]),
        .I3(\u1/u12/X [32]),
        .I4(\u1/u12/X [36]),
        .I5(\u1/u12/X [31]),
        .O(\u1/out12 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__226
       (.I0(\u1/u12/X [11]),
        .I1(\u1/u12/X [10]),
        .I2(\u1/u12/X [9]),
        .I3(\u1/u12/X [8]),
        .I4(\u1/u12/X [12]),
        .I5(\u1/u12/X [7]),
        .O(\u1/out12 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__227
       (.I0(\u1/u12/X [47]),
        .I1(\u1/u12/X [46]),
        .I2(\u1/u12/X [45]),
        .I3(\u1/u12/X [44]),
        .I4(\u1/u12/X [48]),
        .I5(\u1/u12/X [43]),
        .O(\u1/out12 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__228
       (.I0(\u1/u12/X [23]),
        .I1(\u1/u12/X [22]),
        .I2(\u1/u12/X [21]),
        .I3(\u1/u12/X [20]),
        .I4(\u1/u12/X [24]),
        .I5(\u1/u12/X [19]),
        .O(\u1/out12 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__229
       (.I0(\u1/u12/X [29]),
        .I1(\u1/u12/X [28]),
        .I2(\u1/u12/X [27]),
        .I3(\u1/u12/X [26]),
        .I4(\u1/u12/X [30]),
        .I5(\u1/u12/X [25]),
        .O(\u1/out12 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__23
       (.I0(\u0/u3/X [41]),
        .I1(\u0/u3/X [40]),
        .I2(\u0/u3/X [39]),
        .I3(\u0/u3/X [38]),
        .I4(\u0/u3/X [42]),
        .I5(\u0/u3/X [37]),
        .O(\u0/out3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__230
       (.I0(\u1/u12/X [5]),
        .I1(\u1/u12/X [4]),
        .I2(\u1/u12/X [3]),
        .I3(\u1/u12/X [2]),
        .I4(\u1/u12/X [6]),
        .I5(\u1/u12/X [1]),
        .O(\u1/out12 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__231
       (.I0(\u1/u13/X [41]),
        .I1(\u1/u13/X [40]),
        .I2(\u1/u13/X [39]),
        .I3(\u1/u13/X [38]),
        .I4(\u1/u13/X [42]),
        .I5(\u1/u13/X [37]),
        .O(\u1/out13 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__232
       (.I0(\u1/u13/X [17]),
        .I1(\u1/u13/X [16]),
        .I2(\u1/u13/X [15]),
        .I3(\u1/u13/X [14]),
        .I4(\u1/u13/X [18]),
        .I5(\u1/u13/X [13]),
        .O(\u1/out13 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__233
       (.I0(\u1/u13/X [35]),
        .I1(\u1/u13/X [34]),
        .I2(\u1/u13/X [33]),
        .I3(\u1/u13/X [32]),
        .I4(\u1/u13/X [36]),
        .I5(\u1/u13/X [31]),
        .O(\u1/out13 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__234
       (.I0(\u1/u13/X [11]),
        .I1(\u1/u13/X [10]),
        .I2(\u1/u13/X [9]),
        .I3(\u1/u13/X [8]),
        .I4(\u1/u13/X [12]),
        .I5(\u1/u13/X [7]),
        .O(\u1/out13 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__235
       (.I0(\u1/u13/X [47]),
        .I1(\u1/u13/X [46]),
        .I2(\u1/u13/X [45]),
        .I3(\u1/u13/X [44]),
        .I4(\u1/u13/X [48]),
        .I5(\u1/u13/X [43]),
        .O(\u1/out13 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__236
       (.I0(\u1/u13/X [23]),
        .I1(\u1/u13/X [22]),
        .I2(\u1/u13/X [21]),
        .I3(\u1/u13/X [20]),
        .I4(\u1/u13/X [24]),
        .I5(\u1/u13/X [19]),
        .O(\u1/out13 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__237
       (.I0(\u1/u13/X [29]),
        .I1(\u1/u13/X [28]),
        .I2(\u1/u13/X [27]),
        .I3(\u1/u13/X [26]),
        .I4(\u1/u13/X [30]),
        .I5(\u1/u13/X [25]),
        .O(\u1/out13 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__238
       (.I0(\u1/u13/X [5]),
        .I1(\u1/u13/X [4]),
        .I2(\u1/u13/X [3]),
        .I3(\u1/u13/X [2]),
        .I4(\u1/u13/X [6]),
        .I5(\u1/u13/X [1]),
        .O(\u1/out13 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__239
       (.I0(\u1/u14/X [41]),
        .I1(\u1/u14/X [40]),
        .I2(\u1/u14/X [39]),
        .I3(\u1/u14/X [38]),
        .I4(\u1/u14/X [42]),
        .I5(\u1/u14/X [37]),
        .O(\u1/out14 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__24
       (.I0(\u0/u3/X [17]),
        .I1(\u0/u3/X [16]),
        .I2(\u0/u3/X [15]),
        .I3(\u0/u3/X [14]),
        .I4(\u0/u3/X [18]),
        .I5(\u0/u3/X [13]),
        .O(\u0/out3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__240
       (.I0(\u1/u14/X [17]),
        .I1(\u1/u14/X [16]),
        .I2(\u1/u14/X [15]),
        .I3(\u1/u14/X [14]),
        .I4(\u1/u14/X [18]),
        .I5(\u1/u14/X [13]),
        .O(\u1/out14 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__241
       (.I0(\u1/u14/X [35]),
        .I1(\u1/u14/X [34]),
        .I2(\u1/u14/X [33]),
        .I3(\u1/u14/X [32]),
        .I4(\u1/u14/X [36]),
        .I5(\u1/u14/X [31]),
        .O(\u1/out14 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__242
       (.I0(\u1/u14/X [11]),
        .I1(\u1/u14/X [10]),
        .I2(\u1/u14/X [9]),
        .I3(\u1/u14/X [8]),
        .I4(\u1/u14/X [12]),
        .I5(\u1/u14/X [7]),
        .O(\u1/out14 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__243
       (.I0(\u1/u14/X [47]),
        .I1(\u1/u14/X [46]),
        .I2(\u1/u14/X [45]),
        .I3(\u1/u14/X [44]),
        .I4(\u1/u14/X [48]),
        .I5(\u1/u14/X [43]),
        .O(\u1/out14 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__244
       (.I0(\u1/u14/X [23]),
        .I1(\u1/u14/X [22]),
        .I2(\u1/u14/X [21]),
        .I3(\u1/u14/X [20]),
        .I4(\u1/u14/X [24]),
        .I5(\u1/u14/X [19]),
        .O(\u1/out14 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__245
       (.I0(\u1/u14/X [29]),
        .I1(\u1/u14/X [28]),
        .I2(\u1/u14/X [27]),
        .I3(\u1/u14/X [26]),
        .I4(\u1/u14/X [30]),
        .I5(\u1/u14/X [25]),
        .O(\u1/out14 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__246
       (.I0(\u1/u14/X [5]),
        .I1(\u1/u14/X [4]),
        .I2(\u1/u14/X [3]),
        .I3(\u1/u14/X [2]),
        .I4(\u1/u14/X [6]),
        .I5(\u1/u14/X [1]),
        .O(\u1/out14 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__247
       (.I0(\u1/u15/X [41]),
        .I1(\u1/u15/X [40]),
        .I2(\u1/u15/X [39]),
        .I3(\u1/u15/X [38]),
        .I4(\u1/u15/X [42]),
        .I5(\u1/u15/X [37]),
        .O(\u1/out15 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__248
       (.I0(\u1/u15/X [17]),
        .I1(\u1/u15/X [16]),
        .I2(\u1/u15/X [15]),
        .I3(\u1/u15/X [14]),
        .I4(\u1/u15/X [18]),
        .I5(\u1/u15/X [13]),
        .O(\u1/out15 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__249
       (.I0(\u1/u15/X [35]),
        .I1(\u1/u15/X [34]),
        .I2(\u1/u15/X [33]),
        .I3(\u1/u15/X [32]),
        .I4(\u1/u15/X [36]),
        .I5(\u1/u15/X [31]),
        .O(\u1/out15 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__25
       (.I0(\u0/u3/X [35]),
        .I1(\u0/u3/X [34]),
        .I2(\u0/u3/X [33]),
        .I3(\u0/u3/X [32]),
        .I4(\u0/u3/X [36]),
        .I5(\u0/u3/X [31]),
        .O(\u0/out3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__250
       (.I0(\u1/u15/X [11]),
        .I1(\u1/u15/X [10]),
        .I2(\u1/u15/X [9]),
        .I3(\u1/u15/X [8]),
        .I4(\u1/u15/X [12]),
        .I5(\u1/u15/X [7]),
        .O(\u1/out15 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__251
       (.I0(\u1/u15/X [47]),
        .I1(\u1/u15/X [46]),
        .I2(\u1/u15/X [45]),
        .I3(\u1/u15/X [44]),
        .I4(\u1/u15/X [48]),
        .I5(\u1/u15/X [43]),
        .O(\u1/out15 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__252
       (.I0(\u1/u15/X [23]),
        .I1(\u1/u15/X [22]),
        .I2(\u1/u15/X [21]),
        .I3(\u1/u15/X [20]),
        .I4(\u1/u15/X [24]),
        .I5(\u1/u15/X [19]),
        .O(\u1/out15 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__253
       (.I0(\u1/u15/X [29]),
        .I1(\u1/u15/X [28]),
        .I2(\u1/u15/X [27]),
        .I3(\u1/u15/X [26]),
        .I4(\u1/u15/X [30]),
        .I5(\u1/u15/X [25]),
        .O(\u1/out15 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__254
       (.I0(\u1/u15/X [5]),
        .I1(\u1/u15/X [4]),
        .I2(\u1/u15/X [3]),
        .I3(\u1/u15/X [2]),
        .I4(\u1/u15/X [6]),
        .I5(\u1/u15/X [1]),
        .O(\u1/out15 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__255
       (.I0(\u2/u0/X [41]),
        .I1(\u2/u0/X [40]),
        .I2(\u2/u0/X [39]),
        .I3(\u2/u0/X [38]),
        .I4(\u2/u0/X [42]),
        .I5(\u2/u0/X [37]),
        .O(\u2/out0 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__256
       (.I0(\u2/u0/X [17]),
        .I1(\u2/u0/X [16]),
        .I2(\u2/u0/X [15]),
        .I3(\u2/u0/X [14]),
        .I4(\u2/u0/X [18]),
        .I5(\u2/u0/X [13]),
        .O(\u2/out0 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__257
       (.I0(\u2/u0/X [35]),
        .I1(\u2/u0/X [34]),
        .I2(\u2/u0/X [33]),
        .I3(\u2/u0/X [32]),
        .I4(\u2/u0/X [36]),
        .I5(\u2/u0/X [31]),
        .O(\u2/out0 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__258
       (.I0(\u2/u0/X [11]),
        .I1(\u2/u0/X [10]),
        .I2(\u2/u0/X [9]),
        .I3(\u2/u0/X [8]),
        .I4(\u2/u0/X [12]),
        .I5(\u2/u0/X [7]),
        .O(\u2/out0 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__259
       (.I0(\u2/u0/X [47]),
        .I1(\u2/u0/X [46]),
        .I2(\u2/u0/X [45]),
        .I3(\u2/u0/X [44]),
        .I4(\u2/u0/X [48]),
        .I5(\u2/u0/X [43]),
        .O(\u2/out0 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__26
       (.I0(\u0/u3/X [11]),
        .I1(\u0/u3/X [10]),
        .I2(\u0/u3/X [9]),
        .I3(\u0/u3/X [8]),
        .I4(\u0/u3/X [12]),
        .I5(\u0/u3/X [7]),
        .O(\u0/out3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__260
       (.I0(\u2/u0/X [23]),
        .I1(\u2/u0/X [22]),
        .I2(\u2/u0/X [21]),
        .I3(\u2/u0/X [20]),
        .I4(\u2/u0/X [24]),
        .I5(\u2/u0/X [19]),
        .O(\u2/out0 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__261
       (.I0(\u2/u0/X [29]),
        .I1(\u2/u0/X [28]),
        .I2(\u2/u0/X [27]),
        .I3(\u2/u0/X [26]),
        .I4(\u2/u0/X [30]),
        .I5(\u2/u0/X [25]),
        .O(\u2/out0 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__262
       (.I0(\u2/u0/X [5]),
        .I1(\u2/u0/X [4]),
        .I2(\u2/u0/X [3]),
        .I3(\u2/u0/X [2]),
        .I4(\u2/u0/X [6]),
        .I5(\u2/u0/X [1]),
        .O(\u2/out0 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__263
       (.I0(\u2/u1/X [41]),
        .I1(\u2/u1/X [40]),
        .I2(\u2/u1/X [39]),
        .I3(\u2/u1/X [38]),
        .I4(\u2/u1/X [42]),
        .I5(\u2/u1/X [37]),
        .O(\u2/out1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__264
       (.I0(\u2/u1/X [17]),
        .I1(\u2/u1/X [16]),
        .I2(\u2/u1/X [15]),
        .I3(\u2/u1/X [14]),
        .I4(\u2/u1/X [18]),
        .I5(\u2/u1/X [13]),
        .O(\u2/out1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__265
       (.I0(\u2/u1/X [35]),
        .I1(\u2/u1/X [34]),
        .I2(\u2/u1/X [33]),
        .I3(\u2/u1/X [32]),
        .I4(\u2/u1/X [36]),
        .I5(\u2/u1/X [31]),
        .O(\u2/out1 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__266
       (.I0(\u2/u1/X [11]),
        .I1(\u2/u1/X [10]),
        .I2(\u2/u1/X [9]),
        .I3(\u2/u1/X [8]),
        .I4(\u2/u1/X [12]),
        .I5(\u2/u1/X [7]),
        .O(\u2/out1 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__267
       (.I0(\u2/u1/X [47]),
        .I1(\u2/u1/X [46]),
        .I2(\u2/u1/X [45]),
        .I3(\u2/u1/X [44]),
        .I4(\u2/u1/X [48]),
        .I5(\u2/u1/X [43]),
        .O(\u2/out1 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__268
       (.I0(\u2/u1/X [23]),
        .I1(\u2/u1/X [22]),
        .I2(\u2/u1/X [21]),
        .I3(\u2/u1/X [20]),
        .I4(\u2/u1/X [24]),
        .I5(\u2/u1/X [19]),
        .O(\u2/out1 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__269
       (.I0(\u2/u1/X [29]),
        .I1(\u2/u1/X [28]),
        .I2(\u2/u1/X [27]),
        .I3(\u2/u1/X [26]),
        .I4(\u2/u1/X [30]),
        .I5(\u2/u1/X [25]),
        .O(\u2/out1 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__27
       (.I0(\u0/u3/X [47]),
        .I1(\u0/u3/X [46]),
        .I2(\u0/u3/X [45]),
        .I3(\u0/u3/X [44]),
        .I4(\u0/u3/X [48]),
        .I5(\u0/u3/X [43]),
        .O(\u0/out3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__270
       (.I0(\u2/u1/X [5]),
        .I1(\u2/u1/X [4]),
        .I2(\u2/u1/X [3]),
        .I3(\u2/u1/X [2]),
        .I4(\u2/u1/X [6]),
        .I5(\u2/u1/X [1]),
        .O(\u2/out1 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__271
       (.I0(\u2/u2/X [41]),
        .I1(\u2/u2/X [40]),
        .I2(\u2/u2/X [39]),
        .I3(\u2/u2/X [38]),
        .I4(\u2/u2/X [42]),
        .I5(\u2/u2/X [37]),
        .O(\u2/out2 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__272
       (.I0(\u2/u2/X [17]),
        .I1(\u2/u2/X [16]),
        .I2(\u2/u2/X [15]),
        .I3(\u2/u2/X [14]),
        .I4(\u2/u2/X [18]),
        .I5(\u2/u2/X [13]),
        .O(\u2/out2 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__273
       (.I0(\u2/u2/X [35]),
        .I1(\u2/u2/X [34]),
        .I2(\u2/u2/X [33]),
        .I3(\u2/u2/X [32]),
        .I4(\u2/u2/X [36]),
        .I5(\u2/u2/X [31]),
        .O(\u2/out2 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__274
       (.I0(\u2/u2/X [11]),
        .I1(\u2/u2/X [10]),
        .I2(\u2/u2/X [9]),
        .I3(\u2/u2/X [8]),
        .I4(\u2/u2/X [12]),
        .I5(\u2/u2/X [7]),
        .O(\u2/out2 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__275
       (.I0(\u2/u2/X [47]),
        .I1(\u2/u2/X [46]),
        .I2(\u2/u2/X [45]),
        .I3(\u2/u2/X [44]),
        .I4(\u2/u2/X [48]),
        .I5(\u2/u2/X [43]),
        .O(\u2/out2 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__276
       (.I0(\u2/u2/X [23]),
        .I1(\u2/u2/X [22]),
        .I2(\u2/u2/X [21]),
        .I3(\u2/u2/X [20]),
        .I4(\u2/u2/X [24]),
        .I5(\u2/u2/X [19]),
        .O(\u2/out2 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__277
       (.I0(\u2/u2/X [29]),
        .I1(\u2/u2/X [28]),
        .I2(\u2/u2/X [27]),
        .I3(\u2/u2/X [26]),
        .I4(\u2/u2/X [30]),
        .I5(\u2/u2/X [25]),
        .O(\u2/out2 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__278
       (.I0(\u2/u2/X [5]),
        .I1(\u2/u2/X [4]),
        .I2(\u2/u2/X [3]),
        .I3(\u2/u2/X [2]),
        .I4(\u2/u2/X [6]),
        .I5(\u2/u2/X [1]),
        .O(\u2/out2 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__279
       (.I0(\u2/u3/X [41]),
        .I1(\u2/u3/X [40]),
        .I2(\u2/u3/X [39]),
        .I3(\u2/u3/X [38]),
        .I4(\u2/u3/X [42]),
        .I5(\u2/u3/X [37]),
        .O(\u2/out3 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__28
       (.I0(\u0/u3/X [23]),
        .I1(\u0/u3/X [22]),
        .I2(\u0/u3/X [21]),
        .I3(\u0/u3/X [20]),
        .I4(\u0/u3/X [24]),
        .I5(\u0/u3/X [19]),
        .O(\u0/out3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__280
       (.I0(\u2/u3/X [17]),
        .I1(\u2/u3/X [16]),
        .I2(\u2/u3/X [15]),
        .I3(\u2/u3/X [14]),
        .I4(\u2/u3/X [18]),
        .I5(\u2/u3/X [13]),
        .O(\u2/out3 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__281
       (.I0(\u2/u3/X [35]),
        .I1(\u2/u3/X [34]),
        .I2(\u2/u3/X [33]),
        .I3(\u2/u3/X [32]),
        .I4(\u2/u3/X [36]),
        .I5(\u2/u3/X [31]),
        .O(\u2/out3 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__282
       (.I0(\u2/u3/X [11]),
        .I1(\u2/u3/X [10]),
        .I2(\u2/u3/X [9]),
        .I3(\u2/u3/X [8]),
        .I4(\u2/u3/X [12]),
        .I5(\u2/u3/X [7]),
        .O(\u2/out3 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__283
       (.I0(\u2/u3/X [47]),
        .I1(\u2/u3/X [46]),
        .I2(\u2/u3/X [45]),
        .I3(\u2/u3/X [44]),
        .I4(\u2/u3/X [48]),
        .I5(\u2/u3/X [43]),
        .O(\u2/out3 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__284
       (.I0(\u2/u3/X [23]),
        .I1(\u2/u3/X [22]),
        .I2(\u2/u3/X [21]),
        .I3(\u2/u3/X [20]),
        .I4(\u2/u3/X [24]),
        .I5(\u2/u3/X [19]),
        .O(\u2/out3 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__285
       (.I0(\u2/u3/X [29]),
        .I1(\u2/u3/X [28]),
        .I2(\u2/u3/X [27]),
        .I3(\u2/u3/X [26]),
        .I4(\u2/u3/X [30]),
        .I5(\u2/u3/X [25]),
        .O(\u2/out3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__286
       (.I0(\u2/u3/X [5]),
        .I1(\u2/u3/X [4]),
        .I2(\u2/u3/X [3]),
        .I3(\u2/u3/X [2]),
        .I4(\u2/u3/X [6]),
        .I5(\u2/u3/X [1]),
        .O(\u2/out3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__287
       (.I0(\u2/u4/X [41]),
        .I1(\u2/u4/X [40]),
        .I2(\u2/u4/X [39]),
        .I3(\u2/u4/X [38]),
        .I4(\u2/u4/X [42]),
        .I5(\u2/u4/X [37]),
        .O(\u2/out4 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__288
       (.I0(\u2/u4/X [17]),
        .I1(\u2/u4/X [16]),
        .I2(\u2/u4/X [15]),
        .I3(\u2/u4/X [14]),
        .I4(\u2/u4/X [18]),
        .I5(\u2/u4/X [13]),
        .O(\u2/out4 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__289
       (.I0(\u2/u4/X [35]),
        .I1(\u2/u4/X [34]),
        .I2(\u2/u4/X [33]),
        .I3(\u2/u4/X [32]),
        .I4(\u2/u4/X [36]),
        .I5(\u2/u4/X [31]),
        .O(\u2/out4 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__29
       (.I0(\u0/u3/X [29]),
        .I1(\u0/u3/X [28]),
        .I2(\u0/u3/X [27]),
        .I3(\u0/u3/X [26]),
        .I4(\u0/u3/X [30]),
        .I5(\u0/u3/X [25]),
        .O(\u0/out3 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__290
       (.I0(\u2/u4/X [11]),
        .I1(\u2/u4/X [10]),
        .I2(\u2/u4/X [9]),
        .I3(\u2/u4/X [8]),
        .I4(\u2/u4/X [12]),
        .I5(\u2/u4/X [7]),
        .O(\u2/out4 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__291
       (.I0(\u2/u4/X [47]),
        .I1(\u2/u4/X [46]),
        .I2(\u2/u4/X [45]),
        .I3(\u2/u4/X [44]),
        .I4(\u2/u4/X [48]),
        .I5(\u2/u4/X [43]),
        .O(\u2/out4 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__292
       (.I0(\u2/u4/X [23]),
        .I1(\u2/u4/X [22]),
        .I2(\u2/u4/X [21]),
        .I3(\u2/u4/X [20]),
        .I4(\u2/u4/X [24]),
        .I5(\u2/u4/X [19]),
        .O(\u2/out4 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__293
       (.I0(\u2/u4/X [29]),
        .I1(\u2/u4/X [28]),
        .I2(\u2/u4/X [27]),
        .I3(\u2/u4/X [26]),
        .I4(\u2/u4/X [30]),
        .I5(\u2/u4/X [25]),
        .O(\u2/out4 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__294
       (.I0(\u2/u4/X [5]),
        .I1(\u2/u4/X [4]),
        .I2(\u2/u4/X [3]),
        .I3(\u2/u4/X [2]),
        .I4(\u2/u4/X [6]),
        .I5(\u2/u4/X [1]),
        .O(\u2/out4 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__295
       (.I0(\u2/u5/X [41]),
        .I1(\u2/u5/X [40]),
        .I2(\u2/u5/X [39]),
        .I3(\u2/u5/X [38]),
        .I4(\u2/u5/X [42]),
        .I5(\u2/u5/X [37]),
        .O(\u2/out5 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__296
       (.I0(\u2/u5/X [17]),
        .I1(\u2/u5/X [16]),
        .I2(\u2/u5/X [15]),
        .I3(\u2/u5/X [14]),
        .I4(\u2/u5/X [18]),
        .I5(\u2/u5/X [13]),
        .O(\u2/out5 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__297
       (.I0(\u2/u5/X [35]),
        .I1(\u2/u5/X [34]),
        .I2(\u2/u5/X [33]),
        .I3(\u2/u5/X [32]),
        .I4(\u2/u5/X [36]),
        .I5(\u2/u5/X [31]),
        .O(\u2/out5 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__298
       (.I0(\u2/u5/X [11]),
        .I1(\u2/u5/X [10]),
        .I2(\u2/u5/X [9]),
        .I3(\u2/u5/X [8]),
        .I4(\u2/u5/X [12]),
        .I5(\u2/u5/X [7]),
        .O(\u2/out5 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__299
       (.I0(\u2/u5/X [47]),
        .I1(\u2/u5/X [46]),
        .I2(\u2/u5/X [45]),
        .I3(\u2/u5/X [44]),
        .I4(\u2/u5/X [48]),
        .I5(\u2/u5/X [43]),
        .O(\u2/out5 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__3
       (.I0(\u0/u0/X [47]),
        .I1(\u0/u0/X [46]),
        .I2(\u0/u0/X [45]),
        .I3(\u0/u0/X [44]),
        .I4(\u0/u0/X [48]),
        .I5(\u0/u0/X [43]),
        .O(\u0/out0 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__30
       (.I0(\u0/u3/X [5]),
        .I1(\u0/u3/X [4]),
        .I2(\u0/u3/X [3]),
        .I3(\u0/u3/X [2]),
        .I4(\u0/u3/X [6]),
        .I5(\u0/u3/X [1]),
        .O(\u0/out3 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__300
       (.I0(\u2/u5/X [23]),
        .I1(\u2/u5/X [22]),
        .I2(\u2/u5/X [21]),
        .I3(\u2/u5/X [20]),
        .I4(\u2/u5/X [24]),
        .I5(\u2/u5/X [19]),
        .O(\u2/out5 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__301
       (.I0(\u2/u5/X [29]),
        .I1(\u2/u5/X [28]),
        .I2(\u2/u5/X [27]),
        .I3(\u2/u5/X [26]),
        .I4(\u2/u5/X [30]),
        .I5(\u2/u5/X [25]),
        .O(\u2/out5 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__302
       (.I0(\u2/u5/X [5]),
        .I1(\u2/u5/X [4]),
        .I2(\u2/u5/X [3]),
        .I3(\u2/u5/X [2]),
        .I4(\u2/u5/X [6]),
        .I5(\u2/u5/X [1]),
        .O(\u2/out5 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__303
       (.I0(\u2/u6/X [41]),
        .I1(\u2/u6/X [40]),
        .I2(\u2/u6/X [39]),
        .I3(\u2/u6/X [38]),
        .I4(\u2/u6/X [42]),
        .I5(\u2/u6/X [37]),
        .O(\u2/out6 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__304
       (.I0(\u2/u6/X [17]),
        .I1(\u2/u6/X [16]),
        .I2(\u2/u6/X [15]),
        .I3(\u2/u6/X [14]),
        .I4(\u2/u6/X [18]),
        .I5(\u2/u6/X [13]),
        .O(\u2/out6 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__305
       (.I0(\u2/u6/X [35]),
        .I1(\u2/u6/X [34]),
        .I2(\u2/u6/X [33]),
        .I3(\u2/u6/X [32]),
        .I4(\u2/u6/X [36]),
        .I5(\u2/u6/X [31]),
        .O(\u2/out6 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__306
       (.I0(\u2/u6/X [11]),
        .I1(\u2/u6/X [10]),
        .I2(\u2/u6/X [9]),
        .I3(\u2/u6/X [8]),
        .I4(\u2/u6/X [12]),
        .I5(\u2/u6/X [7]),
        .O(\u2/out6 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__307
       (.I0(\u2/u6/X [47]),
        .I1(\u2/u6/X [46]),
        .I2(\u2/u6/X [45]),
        .I3(\u2/u6/X [44]),
        .I4(\u2/u6/X [48]),
        .I5(\u2/u6/X [43]),
        .O(\u2/out6 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__308
       (.I0(\u2/u6/X [23]),
        .I1(\u2/u6/X [22]),
        .I2(\u2/u6/X [21]),
        .I3(\u2/u6/X [20]),
        .I4(\u2/u6/X [24]),
        .I5(\u2/u6/X [19]),
        .O(\u2/out6 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__309
       (.I0(\u2/u6/X [29]),
        .I1(\u2/u6/X [28]),
        .I2(\u2/u6/X [27]),
        .I3(\u2/u6/X [26]),
        .I4(\u2/u6/X [30]),
        .I5(\u2/u6/X [25]),
        .O(\u2/out6 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__31
       (.I0(\u0/u4/X [41]),
        .I1(\u0/u4/X [40]),
        .I2(\u0/u4/X [39]),
        .I3(\u0/u4/X [38]),
        .I4(\u0/u4/X [42]),
        .I5(\u0/u4/X [37]),
        .O(\u0/out4 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__310
       (.I0(\u2/u6/X [5]),
        .I1(\u2/u6/X [4]),
        .I2(\u2/u6/X [3]),
        .I3(\u2/u6/X [2]),
        .I4(\u2/u6/X [6]),
        .I5(\u2/u6/X [1]),
        .O(\u2/out6 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__311
       (.I0(\u2/u7/X [41]),
        .I1(\u2/u7/X [40]),
        .I2(\u2/u7/X [39]),
        .I3(\u2/u7/X [38]),
        .I4(\u2/u7/X [42]),
        .I5(\u2/u7/X [37]),
        .O(\u2/out7 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__312
       (.I0(\u2/u7/X [17]),
        .I1(\u2/u7/X [16]),
        .I2(\u2/u7/X [15]),
        .I3(\u2/u7/X [14]),
        .I4(\u2/u7/X [18]),
        .I5(\u2/u7/X [13]),
        .O(\u2/out7 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__313
       (.I0(\u2/u7/X [35]),
        .I1(\u2/u7/X [34]),
        .I2(\u2/u7/X [33]),
        .I3(\u2/u7/X [32]),
        .I4(\u2/u7/X [36]),
        .I5(\u2/u7/X [31]),
        .O(\u2/out7 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__314
       (.I0(\u2/u7/X [11]),
        .I1(\u2/u7/X [10]),
        .I2(\u2/u7/X [9]),
        .I3(\u2/u7/X [8]),
        .I4(\u2/u7/X [12]),
        .I5(\u2/u7/X [7]),
        .O(\u2/out7 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__315
       (.I0(\u2/u7/X [47]),
        .I1(\u2/u7/X [46]),
        .I2(\u2/u7/X [45]),
        .I3(\u2/u7/X [44]),
        .I4(\u2/u7/X [48]),
        .I5(\u2/u7/X [43]),
        .O(\u2/out7 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__316
       (.I0(\u2/u7/X [23]),
        .I1(\u2/u7/X [22]),
        .I2(\u2/u7/X [21]),
        .I3(\u2/u7/X [20]),
        .I4(\u2/u7/X [24]),
        .I5(\u2/u7/X [19]),
        .O(\u2/out7 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__317
       (.I0(\u2/u7/X [29]),
        .I1(\u2/u7/X [28]),
        .I2(\u2/u7/X [27]),
        .I3(\u2/u7/X [26]),
        .I4(\u2/u7/X [30]),
        .I5(\u2/u7/X [25]),
        .O(\u2/out7 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__318
       (.I0(\u2/u7/X [5]),
        .I1(\u2/u7/X [4]),
        .I2(\u2/u7/X [3]),
        .I3(\u2/u7/X [2]),
        .I4(\u2/u7/X [6]),
        .I5(\u2/u7/X [1]),
        .O(\u2/out7 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__319
       (.I0(\u2/u8/X [41]),
        .I1(\u2/u8/X [40]),
        .I2(\u2/u8/X [39]),
        .I3(\u2/u8/X [38]),
        .I4(\u2/u8/X [42]),
        .I5(\u2/u8/X [37]),
        .O(\u2/out8 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__32
       (.I0(\u0/u4/X [17]),
        .I1(\u0/u4/X [16]),
        .I2(\u0/u4/X [15]),
        .I3(\u0/u4/X [14]),
        .I4(\u0/u4/X [18]),
        .I5(\u0/u4/X [13]),
        .O(\u0/out4 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__320
       (.I0(\u2/u8/X [17]),
        .I1(\u2/u8/X [16]),
        .I2(\u2/u8/X [15]),
        .I3(\u2/u8/X [14]),
        .I4(\u2/u8/X [18]),
        .I5(\u2/u8/X [13]),
        .O(\u2/out8 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__321
       (.I0(\u2/u8/X [35]),
        .I1(\u2/u8/X [34]),
        .I2(\u2/u8/X [33]),
        .I3(\u2/u8/X [32]),
        .I4(\u2/u8/X [36]),
        .I5(\u2/u8/X [31]),
        .O(\u2/out8 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__322
       (.I0(\u2/u8/X [11]),
        .I1(\u2/u8/X [10]),
        .I2(\u2/u8/X [9]),
        .I3(\u2/u8/X [8]),
        .I4(\u2/u8/X [12]),
        .I5(\u2/u8/X [7]),
        .O(\u2/out8 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__323
       (.I0(\u2/u8/X [47]),
        .I1(\u2/u8/X [46]),
        .I2(\u2/u8/X [45]),
        .I3(\u2/u8/X [44]),
        .I4(\u2/u8/X [48]),
        .I5(\u2/u8/X [43]),
        .O(\u2/out8 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__324
       (.I0(\u2/u8/X [23]),
        .I1(\u2/u8/X [22]),
        .I2(\u2/u8/X [21]),
        .I3(\u2/u8/X [20]),
        .I4(\u2/u8/X [24]),
        .I5(\u2/u8/X [19]),
        .O(\u2/out8 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__325
       (.I0(\u2/u8/X [29]),
        .I1(\u2/u8/X [28]),
        .I2(\u2/u8/X [27]),
        .I3(\u2/u8/X [26]),
        .I4(\u2/u8/X [30]),
        .I5(\u2/u8/X [25]),
        .O(\u2/out8 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__326
       (.I0(\u2/u8/X [5]),
        .I1(\u2/u8/X [4]),
        .I2(\u2/u8/X [3]),
        .I3(\u2/u8/X [2]),
        .I4(\u2/u8/X [6]),
        .I5(\u2/u8/X [1]),
        .O(\u2/out8 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__327
       (.I0(\u2/u9/X [41]),
        .I1(\u2/u9/X [40]),
        .I2(\u2/u9/X [39]),
        .I3(\u2/u9/X [38]),
        .I4(\u2/u9/X [42]),
        .I5(\u2/u9/X [37]),
        .O(\u2/out9 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__328
       (.I0(\u2/u9/X [17]),
        .I1(\u2/u9/X [16]),
        .I2(\u2/u9/X [15]),
        .I3(\u2/u9/X [14]),
        .I4(\u2/u9/X [18]),
        .I5(\u2/u9/X [13]),
        .O(\u2/out9 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__329
       (.I0(\u2/u9/X [35]),
        .I1(\u2/u9/X [34]),
        .I2(\u2/u9/X [33]),
        .I3(\u2/u9/X [32]),
        .I4(\u2/u9/X [36]),
        .I5(\u2/u9/X [31]),
        .O(\u2/out9 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__33
       (.I0(\u0/u4/X [35]),
        .I1(\u0/u4/X [34]),
        .I2(\u0/u4/X [33]),
        .I3(\u0/u4/X [32]),
        .I4(\u0/u4/X [36]),
        .I5(\u0/u4/X [31]),
        .O(\u0/out4 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__330
       (.I0(\u2/u9/X [11]),
        .I1(\u2/u9/X [10]),
        .I2(\u2/u9/X [9]),
        .I3(\u2/u9/X [8]),
        .I4(\u2/u9/X [12]),
        .I5(\u2/u9/X [7]),
        .O(\u2/out9 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__331
       (.I0(\u2/u9/X [47]),
        .I1(\u2/u9/X [46]),
        .I2(\u2/u9/X [45]),
        .I3(\u2/u9/X [44]),
        .I4(\u2/u9/X [48]),
        .I5(\u2/u9/X [43]),
        .O(\u2/out9 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__332
       (.I0(\u2/u9/X [23]),
        .I1(\u2/u9/X [22]),
        .I2(\u2/u9/X [21]),
        .I3(\u2/u9/X [20]),
        .I4(\u2/u9/X [24]),
        .I5(\u2/u9/X [19]),
        .O(\u2/out9 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__333
       (.I0(\u2/u9/X [29]),
        .I1(\u2/u9/X [28]),
        .I2(\u2/u9/X [27]),
        .I3(\u2/u9/X [26]),
        .I4(\u2/u9/X [30]),
        .I5(\u2/u9/X [25]),
        .O(\u2/out9 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__334
       (.I0(\u2/u9/X [5]),
        .I1(\u2/u9/X [4]),
        .I2(\u2/u9/X [3]),
        .I3(\u2/u9/X [2]),
        .I4(\u2/u9/X [6]),
        .I5(\u2/u9/X [1]),
        .O(\u2/out9 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__335
       (.I0(\u2/u10/X [41]),
        .I1(\u2/u10/X [40]),
        .I2(\u2/u10/X [39]),
        .I3(\u2/u10/X [38]),
        .I4(\u2/u10/X [42]),
        .I5(\u2/u10/X [37]),
        .O(\u2/out10 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__336
       (.I0(\u2/u10/X [17]),
        .I1(\u2/u10/X [16]),
        .I2(\u2/u10/X [15]),
        .I3(\u2/u10/X [14]),
        .I4(\u2/u10/X [18]),
        .I5(\u2/u10/X [13]),
        .O(\u2/out10 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__337
       (.I0(\u2/u10/X [35]),
        .I1(\u2/u10/X [34]),
        .I2(\u2/u10/X [33]),
        .I3(\u2/u10/X [32]),
        .I4(\u2/u10/X [36]),
        .I5(\u2/u10/X [31]),
        .O(\u2/out10 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__338
       (.I0(\u2/u10/X [11]),
        .I1(\u2/u10/X [10]),
        .I2(\u2/u10/X [9]),
        .I3(\u2/u10/X [8]),
        .I4(\u2/u10/X [12]),
        .I5(\u2/u10/X [7]),
        .O(\u2/out10 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__339
       (.I0(\u2/u10/X [47]),
        .I1(\u2/u10/X [46]),
        .I2(\u2/u10/X [45]),
        .I3(\u2/u10/X [44]),
        .I4(\u2/u10/X [48]),
        .I5(\u2/u10/X [43]),
        .O(\u2/out10 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__34
       (.I0(\u0/u4/X [11]),
        .I1(\u0/u4/X [10]),
        .I2(\u0/u4/X [9]),
        .I3(\u0/u4/X [8]),
        .I4(\u0/u4/X [12]),
        .I5(\u0/u4/X [7]),
        .O(\u0/out4 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__340
       (.I0(\u2/u10/X [23]),
        .I1(\u2/u10/X [22]),
        .I2(\u2/u10/X [21]),
        .I3(\u2/u10/X [20]),
        .I4(\u2/u10/X [24]),
        .I5(\u2/u10/X [19]),
        .O(\u2/out10 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__341
       (.I0(\u2/u10/X [29]),
        .I1(\u2/u10/X [28]),
        .I2(\u2/u10/X [27]),
        .I3(\u2/u10/X [26]),
        .I4(\u2/u10/X [30]),
        .I5(\u2/u10/X [25]),
        .O(\u2/out10 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__342
       (.I0(\u2/u10/X [5]),
        .I1(\u2/u10/X [4]),
        .I2(\u2/u10/X [3]),
        .I3(\u2/u10/X [2]),
        .I4(\u2/u10/X [6]),
        .I5(\u2/u10/X [1]),
        .O(\u2/out10 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__343
       (.I0(\u2/u11/X [41]),
        .I1(\u2/u11/X [40]),
        .I2(\u2/u11/X [39]),
        .I3(\u2/u11/X [38]),
        .I4(\u2/u11/X [42]),
        .I5(\u2/u11/X [37]),
        .O(\u2/out11 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__344
       (.I0(\u2/u11/X [17]),
        .I1(\u2/u11/X [16]),
        .I2(\u2/u11/X [15]),
        .I3(\u2/u11/X [14]),
        .I4(\u2/u11/X [18]),
        .I5(\u2/u11/X [13]),
        .O(\u2/out11 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__345
       (.I0(\u2/u11/X [35]),
        .I1(\u2/u11/X [34]),
        .I2(\u2/u11/X [33]),
        .I3(\u2/u11/X [32]),
        .I4(\u2/u11/X [36]),
        .I5(\u2/u11/X [31]),
        .O(\u2/out11 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__346
       (.I0(\u2/u11/X [11]),
        .I1(\u2/u11/X [10]),
        .I2(\u2/u11/X [9]),
        .I3(\u2/u11/X [8]),
        .I4(\u2/u11/X [12]),
        .I5(\u2/u11/X [7]),
        .O(\u2/out11 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__347
       (.I0(\u2/u11/X [47]),
        .I1(\u2/u11/X [46]),
        .I2(\u2/u11/X [45]),
        .I3(\u2/u11/X [44]),
        .I4(\u2/u11/X [48]),
        .I5(\u2/u11/X [43]),
        .O(\u2/out11 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__348
       (.I0(\u2/u11/X [23]),
        .I1(\u2/u11/X [22]),
        .I2(\u2/u11/X [21]),
        .I3(\u2/u11/X [20]),
        .I4(\u2/u11/X [24]),
        .I5(\u2/u11/X [19]),
        .O(\u2/out11 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__349
       (.I0(\u2/u11/X [29]),
        .I1(\u2/u11/X [28]),
        .I2(\u2/u11/X [27]),
        .I3(\u2/u11/X [26]),
        .I4(\u2/u11/X [30]),
        .I5(\u2/u11/X [25]),
        .O(\u2/out11 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__35
       (.I0(\u0/u4/X [47]),
        .I1(\u0/u4/X [46]),
        .I2(\u0/u4/X [45]),
        .I3(\u0/u4/X [44]),
        .I4(\u0/u4/X [48]),
        .I5(\u0/u4/X [43]),
        .O(\u0/out4 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__350
       (.I0(\u2/u11/X [5]),
        .I1(\u2/u11/X [4]),
        .I2(\u2/u11/X [3]),
        .I3(\u2/u11/X [2]),
        .I4(\u2/u11/X [6]),
        .I5(\u2/u11/X [1]),
        .O(\u2/out11 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__351
       (.I0(\u2/u12/X [41]),
        .I1(\u2/u12/X [40]),
        .I2(\u2/u12/X [39]),
        .I3(\u2/u12/X [38]),
        .I4(\u2/u12/X [42]),
        .I5(\u2/u12/X [37]),
        .O(\u2/out12 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__352
       (.I0(\u2/u12/X [17]),
        .I1(\u2/u12/X [16]),
        .I2(\u2/u12/X [15]),
        .I3(\u2/u12/X [14]),
        .I4(\u2/u12/X [18]),
        .I5(\u2/u12/X [13]),
        .O(\u2/out12 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__353
       (.I0(\u2/u12/X [35]),
        .I1(\u2/u12/X [34]),
        .I2(\u2/u12/X [33]),
        .I3(\u2/u12/X [32]),
        .I4(\u2/u12/X [36]),
        .I5(\u2/u12/X [31]),
        .O(\u2/out12 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__354
       (.I0(\u2/u12/X [11]),
        .I1(\u2/u12/X [10]),
        .I2(\u2/u12/X [9]),
        .I3(\u2/u12/X [8]),
        .I4(\u2/u12/X [12]),
        .I5(\u2/u12/X [7]),
        .O(\u2/out12 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__355
       (.I0(\u2/u12/X [47]),
        .I1(\u2/u12/X [46]),
        .I2(\u2/u12/X [45]),
        .I3(\u2/u12/X [44]),
        .I4(\u2/u12/X [48]),
        .I5(\u2/u12/X [43]),
        .O(\u2/out12 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__356
       (.I0(\u2/u12/X [23]),
        .I1(\u2/u12/X [22]),
        .I2(\u2/u12/X [21]),
        .I3(\u2/u12/X [20]),
        .I4(\u2/u12/X [24]),
        .I5(\u2/u12/X [19]),
        .O(\u2/out12 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__357
       (.I0(\u2/u12/X [29]),
        .I1(\u2/u12/X [28]),
        .I2(\u2/u12/X [27]),
        .I3(\u2/u12/X [26]),
        .I4(\u2/u12/X [30]),
        .I5(\u2/u12/X [25]),
        .O(\u2/out12 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__358
       (.I0(\u2/u12/X [5]),
        .I1(\u2/u12/X [4]),
        .I2(\u2/u12/X [3]),
        .I3(\u2/u12/X [2]),
        .I4(\u2/u12/X [6]),
        .I5(\u2/u12/X [1]),
        .O(\u2/out12 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__359
       (.I0(\u2/u13/X [41]),
        .I1(\u2/u13/X [40]),
        .I2(\u2/u13/X [39]),
        .I3(\u2/u13/X [38]),
        .I4(\u2/u13/X [42]),
        .I5(\u2/u13/X [37]),
        .O(\u2/out13 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__36
       (.I0(\u0/u4/X [23]),
        .I1(\u0/u4/X [22]),
        .I2(\u0/u4/X [21]),
        .I3(\u0/u4/X [20]),
        .I4(\u0/u4/X [24]),
        .I5(\u0/u4/X [19]),
        .O(\u0/out4 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__360
       (.I0(\u2/u13/X [17]),
        .I1(\u2/u13/X [16]),
        .I2(\u2/u13/X [15]),
        .I3(\u2/u13/X [14]),
        .I4(\u2/u13/X [18]),
        .I5(\u2/u13/X [13]),
        .O(\u2/out13 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__361
       (.I0(\u2/u13/X [35]),
        .I1(\u2/u13/X [34]),
        .I2(\u2/u13/X [33]),
        .I3(\u2/u13/X [32]),
        .I4(\u2/u13/X [36]),
        .I5(\u2/u13/X [31]),
        .O(\u2/out13 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__362
       (.I0(\u2/u13/X [11]),
        .I1(\u2/u13/X [10]),
        .I2(\u2/u13/X [9]),
        .I3(\u2/u13/X [8]),
        .I4(\u2/u13/X [12]),
        .I5(\u2/u13/X [7]),
        .O(\u2/out13 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__363
       (.I0(\u2/u13/X [47]),
        .I1(\u2/u13/X [46]),
        .I2(\u2/u13/X [45]),
        .I3(\u2/u13/X [44]),
        .I4(\u2/u13/X [48]),
        .I5(\u2/u13/X [43]),
        .O(\u2/out13 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__364
       (.I0(\u2/u13/X [23]),
        .I1(\u2/u13/X [22]),
        .I2(\u2/u13/X [21]),
        .I3(\u2/u13/X [20]),
        .I4(\u2/u13/X [24]),
        .I5(\u2/u13/X [19]),
        .O(\u2/out13 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__365
       (.I0(\u2/u13/X [29]),
        .I1(\u2/u13/X [28]),
        .I2(\u2/u13/X [27]),
        .I3(\u2/u13/X [26]),
        .I4(\u2/u13/X [30]),
        .I5(\u2/u13/X [25]),
        .O(\u2/out13 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__366
       (.I0(\u2/u13/X [5]),
        .I1(\u2/u13/X [4]),
        .I2(\u2/u13/X [3]),
        .I3(\u2/u13/X [2]),
        .I4(\u2/u13/X [6]),
        .I5(\u2/u13/X [1]),
        .O(\u2/out13 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__367
       (.I0(\u2/u14/X [41]),
        .I1(\u2/u14/X [40]),
        .I2(\u2/u14/X [39]),
        .I3(\u2/u14/X [38]),
        .I4(\u2/u14/X [42]),
        .I5(\u2/u14/X [37]),
        .O(\u2/out14 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__368
       (.I0(\u2/u14/X [17]),
        .I1(\u2/u14/X [16]),
        .I2(\u2/u14/X [15]),
        .I3(\u2/u14/X [14]),
        .I4(\u2/u14/X [18]),
        .I5(\u2/u14/X [13]),
        .O(\u2/out14 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__369
       (.I0(\u2/u14/X [35]),
        .I1(\u2/u14/X [34]),
        .I2(\u2/u14/X [33]),
        .I3(\u2/u14/X [32]),
        .I4(\u2/u14/X [36]),
        .I5(\u2/u14/X [31]),
        .O(\u2/out14 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__37
       (.I0(\u0/u4/X [29]),
        .I1(\u0/u4/X [28]),
        .I2(\u0/u4/X [27]),
        .I3(\u0/u4/X [26]),
        .I4(\u0/u4/X [30]),
        .I5(\u0/u4/X [25]),
        .O(\u0/out4 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__370
       (.I0(\u2/u14/X [11]),
        .I1(\u2/u14/X [10]),
        .I2(\u2/u14/X [9]),
        .I3(\u2/u14/X [8]),
        .I4(\u2/u14/X [12]),
        .I5(\u2/u14/X [7]),
        .O(\u2/out14 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__371
       (.I0(\u2/u14/X [47]),
        .I1(\u2/u14/X [46]),
        .I2(\u2/u14/X [45]),
        .I3(\u2/u14/X [44]),
        .I4(\u2/u14/X [48]),
        .I5(\u2/u14/X [43]),
        .O(\u2/out14 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__372
       (.I0(\u2/u14/X [23]),
        .I1(\u2/u14/X [22]),
        .I2(\u2/u14/X [21]),
        .I3(\u2/u14/X [20]),
        .I4(\u2/u14/X [24]),
        .I5(\u2/u14/X [19]),
        .O(\u2/out14 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__373
       (.I0(\u2/u14/X [29]),
        .I1(\u2/u14/X [28]),
        .I2(\u2/u14/X [27]),
        .I3(\u2/u14/X [26]),
        .I4(\u2/u14/X [30]),
        .I5(\u2/u14/X [25]),
        .O(\u2/out14 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__374
       (.I0(\u2/u14/X [5]),
        .I1(\u2/u14/X [4]),
        .I2(\u2/u14/X [3]),
        .I3(\u2/u14/X [2]),
        .I4(\u2/u14/X [6]),
        .I5(\u2/u14/X [1]),
        .O(\u2/out14 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__375
       (.I0(\u2/u15/X [41]),
        .I1(\u2/u15/X [40]),
        .I2(\u2/u15/X [39]),
        .I3(\u2/u15/X [38]),
        .I4(\u2/u15/X [42]),
        .I5(\u2/u15/X [37]),
        .O(\u2/out15 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__376
       (.I0(\u2/u15/X [17]),
        .I1(\u2/u15/X [16]),
        .I2(\u2/u15/X [15]),
        .I3(\u2/u15/X [14]),
        .I4(\u2/u15/X [18]),
        .I5(\u2/u15/X [13]),
        .O(\u2/out15 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__377
       (.I0(\u2/u15/X [35]),
        .I1(\u2/u15/X [34]),
        .I2(\u2/u15/X [33]),
        .I3(\u2/u15/X [32]),
        .I4(\u2/u15/X [36]),
        .I5(\u2/u15/X [31]),
        .O(\u2/out15 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__378
       (.I0(\u2/u15/X [11]),
        .I1(\u2/u15/X [10]),
        .I2(\u2/u15/X [9]),
        .I3(\u2/u15/X [8]),
        .I4(\u2/u15/X [12]),
        .I5(\u2/u15/X [7]),
        .O(\u2/out15 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__379
       (.I0(\u2/u15/X [47]),
        .I1(\u2/u15/X [46]),
        .I2(\u2/u15/X [45]),
        .I3(\u2/u15/X [44]),
        .I4(\u2/u15/X [48]),
        .I5(\u2/u15/X [43]),
        .O(\u2/out15 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__38
       (.I0(\u0/u4/X [5]),
        .I1(\u0/u4/X [4]),
        .I2(\u0/u4/X [3]),
        .I3(\u0/u4/X [2]),
        .I4(\u0/u4/X [6]),
        .I5(\u0/u4/X [1]),
        .O(\u0/out4 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__380
       (.I0(\u2/u15/X [23]),
        .I1(\u2/u15/X [22]),
        .I2(\u2/u15/X [21]),
        .I3(\u2/u15/X [20]),
        .I4(\u2/u15/X [24]),
        .I5(\u2/u15/X [19]),
        .O(\u2/out15 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__381
       (.I0(\u2/u15/X [29]),
        .I1(\u2/u15/X [28]),
        .I2(\u2/u15/X [27]),
        .I3(\u2/u15/X [26]),
        .I4(\u2/u15/X [30]),
        .I5(\u2/u15/X [25]),
        .O(\u2/out15 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__382
       (.I0(\u2/u15/X [5]),
        .I1(\u2/u15/X [4]),
        .I2(\u2/u15/X [3]),
        .I3(\u2/u15/X [2]),
        .I4(\u2/u15/X [6]),
        .I5(\u2/u15/X [1]),
        .O(\u2/out15 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__39
       (.I0(\u0/u5/X [41]),
        .I1(\u0/u5/X [40]),
        .I2(\u0/u5/X [39]),
        .I3(\u0/u5/X [38]),
        .I4(\u0/u5/X [42]),
        .I5(\u0/u5/X [37]),
        .O(\u0/out5 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__4
       (.I0(\u0/u0/X [23]),
        .I1(\u0/u0/X [22]),
        .I2(\u0/u0/X [21]),
        .I3(\u0/u0/X [20]),
        .I4(\u0/u0/X [24]),
        .I5(\u0/u0/X [19]),
        .O(\u0/out0 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__40
       (.I0(\u0/u5/X [17]),
        .I1(\u0/u5/X [16]),
        .I2(\u0/u5/X [15]),
        .I3(\u0/u5/X [14]),
        .I4(\u0/u5/X [18]),
        .I5(\u0/u5/X [13]),
        .O(\u0/out5 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__41
       (.I0(\u0/u5/X [35]),
        .I1(\u0/u5/X [34]),
        .I2(\u0/u5/X [33]),
        .I3(\u0/u5/X [32]),
        .I4(\u0/u5/X [36]),
        .I5(\u0/u5/X [31]),
        .O(\u0/out5 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__42
       (.I0(\u0/u5/X [11]),
        .I1(\u0/u5/X [10]),
        .I2(\u0/u5/X [9]),
        .I3(\u0/u5/X [8]),
        .I4(\u0/u5/X [12]),
        .I5(\u0/u5/X [7]),
        .O(\u0/out5 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__43
       (.I0(\u0/u5/X [47]),
        .I1(\u0/u5/X [46]),
        .I2(\u0/u5/X [45]),
        .I3(\u0/u5/X [44]),
        .I4(\u0/u5/X [48]),
        .I5(\u0/u5/X [43]),
        .O(\u0/out5 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__44
       (.I0(\u0/u5/X [23]),
        .I1(\u0/u5/X [22]),
        .I2(\u0/u5/X [21]),
        .I3(\u0/u5/X [20]),
        .I4(\u0/u5/X [24]),
        .I5(\u0/u5/X [19]),
        .O(\u0/out5 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__45
       (.I0(\u0/u5/X [29]),
        .I1(\u0/u5/X [28]),
        .I2(\u0/u5/X [27]),
        .I3(\u0/u5/X [26]),
        .I4(\u0/u5/X [30]),
        .I5(\u0/u5/X [25]),
        .O(\u0/out5 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__46
       (.I0(\u0/u5/X [5]),
        .I1(\u0/u5/X [4]),
        .I2(\u0/u5/X [3]),
        .I3(\u0/u5/X [2]),
        .I4(\u0/u5/X [6]),
        .I5(\u0/u5/X [1]),
        .O(\u0/out5 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__47
       (.I0(\u0/u6/X [41]),
        .I1(\u0/u6/X [40]),
        .I2(\u0/u6/X [39]),
        .I3(\u0/u6/X [38]),
        .I4(\u0/u6/X [42]),
        .I5(\u0/u6/X [37]),
        .O(\u0/out6 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__48
       (.I0(\u0/u6/X [17]),
        .I1(\u0/u6/X [16]),
        .I2(\u0/u6/X [15]),
        .I3(\u0/u6/X [14]),
        .I4(\u0/u6/X [18]),
        .I5(\u0/u6/X [13]),
        .O(\u0/out6 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__49
       (.I0(\u0/u6/X [35]),
        .I1(\u0/u6/X [34]),
        .I2(\u0/u6/X [33]),
        .I3(\u0/u6/X [32]),
        .I4(\u0/u6/X [36]),
        .I5(\u0/u6/X [31]),
        .O(\u0/out6 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__5
       (.I0(\u0/u0/X [29]),
        .I1(\u0/u0/X [28]),
        .I2(\u0/u0/X [27]),
        .I3(\u0/u0/X [26]),
        .I4(\u0/u0/X [30]),
        .I5(\u0/u0/X [25]),
        .O(\u0/out0 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__50
       (.I0(\u0/u6/X [11]),
        .I1(\u0/u6/X [10]),
        .I2(\u0/u6/X [9]),
        .I3(\u0/u6/X [8]),
        .I4(\u0/u6/X [12]),
        .I5(\u0/u6/X [7]),
        .O(\u0/out6 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__51
       (.I0(\u0/u6/X [47]),
        .I1(\u0/u6/X [46]),
        .I2(\u0/u6/X [45]),
        .I3(\u0/u6/X [44]),
        .I4(\u0/u6/X [48]),
        .I5(\u0/u6/X [43]),
        .O(\u0/out6 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__52
       (.I0(\u0/u6/X [23]),
        .I1(\u0/u6/X [22]),
        .I2(\u0/u6/X [21]),
        .I3(\u0/u6/X [20]),
        .I4(\u0/u6/X [24]),
        .I5(\u0/u6/X [19]),
        .O(\u0/out6 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__53
       (.I0(\u0/u6/X [29]),
        .I1(\u0/u6/X [28]),
        .I2(\u0/u6/X [27]),
        .I3(\u0/u6/X [26]),
        .I4(\u0/u6/X [30]),
        .I5(\u0/u6/X [25]),
        .O(\u0/out6 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__54
       (.I0(\u0/u6/X [5]),
        .I1(\u0/u6/X [4]),
        .I2(\u0/u6/X [3]),
        .I3(\u0/u6/X [2]),
        .I4(\u0/u6/X [6]),
        .I5(\u0/u6/X [1]),
        .O(\u0/out6 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__55
       (.I0(\u0/u7/X [41]),
        .I1(\u0/u7/X [40]),
        .I2(\u0/u7/X [39]),
        .I3(\u0/u7/X [38]),
        .I4(\u0/u7/X [42]),
        .I5(\u0/u7/X [37]),
        .O(\u0/out7 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__56
       (.I0(\u0/u7/X [17]),
        .I1(\u0/u7/X [16]),
        .I2(\u0/u7/X [15]),
        .I3(\u0/u7/X [14]),
        .I4(\u0/u7/X [18]),
        .I5(\u0/u7/X [13]),
        .O(\u0/out7 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__57
       (.I0(\u0/u7/X [35]),
        .I1(\u0/u7/X [34]),
        .I2(\u0/u7/X [33]),
        .I3(\u0/u7/X [32]),
        .I4(\u0/u7/X [36]),
        .I5(\u0/u7/X [31]),
        .O(\u0/out7 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__58
       (.I0(\u0/u7/X [11]),
        .I1(\u0/u7/X [10]),
        .I2(\u0/u7/X [9]),
        .I3(\u0/u7/X [8]),
        .I4(\u0/u7/X [12]),
        .I5(\u0/u7/X [7]),
        .O(\u0/out7 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__59
       (.I0(\u0/u7/X [47]),
        .I1(\u0/u7/X [46]),
        .I2(\u0/u7/X [45]),
        .I3(\u0/u7/X [44]),
        .I4(\u0/u7/X [48]),
        .I5(\u0/u7/X [43]),
        .O(\u0/out7 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__6
       (.I0(\u0/u0/X [5]),
        .I1(\u0/u0/X [4]),
        .I2(\u0/u0/X [3]),
        .I3(\u0/u0/X [2]),
        .I4(\u0/u0/X [6]),
        .I5(\u0/u0/X [1]),
        .O(\u0/out0 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__60
       (.I0(\u0/u7/X [23]),
        .I1(\u0/u7/X [22]),
        .I2(\u0/u7/X [21]),
        .I3(\u0/u7/X [20]),
        .I4(\u0/u7/X [24]),
        .I5(\u0/u7/X [19]),
        .O(\u0/out7 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__61
       (.I0(\u0/u7/X [29]),
        .I1(\u0/u7/X [28]),
        .I2(\u0/u7/X [27]),
        .I3(\u0/u7/X [26]),
        .I4(\u0/u7/X [30]),
        .I5(\u0/u7/X [25]),
        .O(\u0/out7 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__62
       (.I0(\u0/u7/X [5]),
        .I1(\u0/u7/X [4]),
        .I2(\u0/u7/X [3]),
        .I3(\u0/u7/X [2]),
        .I4(\u0/u7/X [6]),
        .I5(\u0/u7/X [1]),
        .O(\u0/out7 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__63
       (.I0(\u0/u8/X [41]),
        .I1(\u0/u8/X [40]),
        .I2(\u0/u8/X [39]),
        .I3(\u0/u8/X [38]),
        .I4(\u0/u8/X [42]),
        .I5(\u0/u8/X [37]),
        .O(\u0/out8 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__64
       (.I0(\u0/u8/X [17]),
        .I1(\u0/u8/X [16]),
        .I2(\u0/u8/X [15]),
        .I3(\u0/u8/X [14]),
        .I4(\u0/u8/X [18]),
        .I5(\u0/u8/X [13]),
        .O(\u0/out8 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__65
       (.I0(\u0/u8/X [35]),
        .I1(\u0/u8/X [34]),
        .I2(\u0/u8/X [33]),
        .I3(\u0/u8/X [32]),
        .I4(\u0/u8/X [36]),
        .I5(\u0/u8/X [31]),
        .O(\u0/out8 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__66
       (.I0(\u0/u8/X [11]),
        .I1(\u0/u8/X [10]),
        .I2(\u0/u8/X [9]),
        .I3(\u0/u8/X [8]),
        .I4(\u0/u8/X [12]),
        .I5(\u0/u8/X [7]),
        .O(\u0/out8 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__67
       (.I0(\u0/u8/X [47]),
        .I1(\u0/u8/X [46]),
        .I2(\u0/u8/X [45]),
        .I3(\u0/u8/X [44]),
        .I4(\u0/u8/X [48]),
        .I5(\u0/u8/X [43]),
        .O(\u0/out8 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__68
       (.I0(\u0/u8/X [23]),
        .I1(\u0/u8/X [22]),
        .I2(\u0/u8/X [21]),
        .I3(\u0/u8/X [20]),
        .I4(\u0/u8/X [24]),
        .I5(\u0/u8/X [19]),
        .O(\u0/out8 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__69
       (.I0(\u0/u8/X [29]),
        .I1(\u0/u8/X [28]),
        .I2(\u0/u8/X [27]),
        .I3(\u0/u8/X [26]),
        .I4(\u0/u8/X [30]),
        .I5(\u0/u8/X [25]),
        .O(\u0/out8 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__7
       (.I0(\u0/u1/X [41]),
        .I1(\u0/u1/X [40]),
        .I2(\u0/u1/X [39]),
        .I3(\u0/u1/X [38]),
        .I4(\u0/u1/X [42]),
        .I5(\u0/u1/X [37]),
        .O(\u0/out1 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__70
       (.I0(\u0/u8/X [5]),
        .I1(\u0/u8/X [4]),
        .I2(\u0/u8/X [3]),
        .I3(\u0/u8/X [2]),
        .I4(\u0/u8/X [6]),
        .I5(\u0/u8/X [1]),
        .O(\u0/out8 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__71
       (.I0(\u0/u9/X [41]),
        .I1(\u0/u9/X [40]),
        .I2(\u0/u9/X [39]),
        .I3(\u0/u9/X [38]),
        .I4(\u0/u9/X [42]),
        .I5(\u0/u9/X [37]),
        .O(\u0/out9 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__72
       (.I0(\u0/u9/X [17]),
        .I1(\u0/u9/X [16]),
        .I2(\u0/u9/X [15]),
        .I3(\u0/u9/X [14]),
        .I4(\u0/u9/X [18]),
        .I5(\u0/u9/X [13]),
        .O(\u0/out9 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__73
       (.I0(\u0/u9/X [35]),
        .I1(\u0/u9/X [34]),
        .I2(\u0/u9/X [33]),
        .I3(\u0/u9/X [32]),
        .I4(\u0/u9/X [36]),
        .I5(\u0/u9/X [31]),
        .O(\u0/out9 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__74
       (.I0(\u0/u9/X [11]),
        .I1(\u0/u9/X [10]),
        .I2(\u0/u9/X [9]),
        .I3(\u0/u9/X [8]),
        .I4(\u0/u9/X [12]),
        .I5(\u0/u9/X [7]),
        .O(\u0/out9 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__75
       (.I0(\u0/u9/X [47]),
        .I1(\u0/u9/X [46]),
        .I2(\u0/u9/X [45]),
        .I3(\u0/u9/X [44]),
        .I4(\u0/u9/X [48]),
        .I5(\u0/u9/X [43]),
        .O(\u0/out9 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__76
       (.I0(\u0/u9/X [23]),
        .I1(\u0/u9/X [22]),
        .I2(\u0/u9/X [21]),
        .I3(\u0/u9/X [20]),
        .I4(\u0/u9/X [24]),
        .I5(\u0/u9/X [19]),
        .O(\u0/out9 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__77
       (.I0(\u0/u9/X [29]),
        .I1(\u0/u9/X [28]),
        .I2(\u0/u9/X [27]),
        .I3(\u0/u9/X [26]),
        .I4(\u0/u9/X [30]),
        .I5(\u0/u9/X [25]),
        .O(\u0/out9 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__78
       (.I0(\u0/u9/X [5]),
        .I1(\u0/u9/X [4]),
        .I2(\u0/u9/X [3]),
        .I3(\u0/u9/X [2]),
        .I4(\u0/u9/X [6]),
        .I5(\u0/u9/X [1]),
        .O(\u0/out9 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__79
       (.I0(\u0/u10/X [41]),
        .I1(\u0/u10/X [40]),
        .I2(\u0/u10/X [39]),
        .I3(\u0/u10/X [38]),
        .I4(\u0/u10/X [42]),
        .I5(\u0/u10/X [37]),
        .O(\u0/out10 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__8
       (.I0(\u0/u1/X [17]),
        .I1(\u0/u1/X [16]),
        .I2(\u0/u1/X [15]),
        .I3(\u0/u1/X [14]),
        .I4(\u0/u1/X [18]),
        .I5(\u0/u1/X [13]),
        .O(\u0/out1 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__80
       (.I0(\u0/u10/X [17]),
        .I1(\u0/u10/X [16]),
        .I2(\u0/u10/X [15]),
        .I3(\u0/u10/X [14]),
        .I4(\u0/u10/X [18]),
        .I5(\u0/u10/X [13]),
        .O(\u0/out10 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__81
       (.I0(\u0/u10/X [35]),
        .I1(\u0/u10/X [34]),
        .I2(\u0/u10/X [33]),
        .I3(\u0/u10/X [32]),
        .I4(\u0/u10/X [36]),
        .I5(\u0/u10/X [31]),
        .O(\u0/out10 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__82
       (.I0(\u0/u10/X [11]),
        .I1(\u0/u10/X [10]),
        .I2(\u0/u10/X [9]),
        .I3(\u0/u10/X [8]),
        .I4(\u0/u10/X [12]),
        .I5(\u0/u10/X [7]),
        .O(\u0/out10 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__83
       (.I0(\u0/u10/X [47]),
        .I1(\u0/u10/X [46]),
        .I2(\u0/u10/X [45]),
        .I3(\u0/u10/X [44]),
        .I4(\u0/u10/X [48]),
        .I5(\u0/u10/X [43]),
        .O(\u0/out10 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__84
       (.I0(\u0/u10/X [23]),
        .I1(\u0/u10/X [22]),
        .I2(\u0/u10/X [21]),
        .I3(\u0/u10/X [20]),
        .I4(\u0/u10/X [24]),
        .I5(\u0/u10/X [19]),
        .O(\u0/out10 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__85
       (.I0(\u0/u10/X [29]),
        .I1(\u0/u10/X [28]),
        .I2(\u0/u10/X [27]),
        .I3(\u0/u10/X [26]),
        .I4(\u0/u10/X [30]),
        .I5(\u0/u10/X [25]),
        .O(\u0/out10 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__86
       (.I0(\u0/u10/X [5]),
        .I1(\u0/u10/X [4]),
        .I2(\u0/u10/X [3]),
        .I3(\u0/u10/X [2]),
        .I4(\u0/u10/X [6]),
        .I5(\u0/u10/X [1]),
        .O(\u0/out10 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__87
       (.I0(\u0/u11/X [41]),
        .I1(\u0/u11/X [40]),
        .I2(\u0/u11/X [39]),
        .I3(\u0/u11/X [38]),
        .I4(\u0/u11/X [42]),
        .I5(\u0/u11/X [37]),
        .O(\u0/out11 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__88
       (.I0(\u0/u11/X [17]),
        .I1(\u0/u11/X [16]),
        .I2(\u0/u11/X [15]),
        .I3(\u0/u11/X [14]),
        .I4(\u0/u11/X [18]),
        .I5(\u0/u11/X [13]),
        .O(\u0/out11 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__89
       (.I0(\u0/u11/X [35]),
        .I1(\u0/u11/X [34]),
        .I2(\u0/u11/X [33]),
        .I3(\u0/u11/X [32]),
        .I4(\u0/u11/X [36]),
        .I5(\u0/u11/X [31]),
        .O(\u0/out11 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__9
       (.I0(\u0/u1/X [35]),
        .I1(\u0/u1/X [34]),
        .I2(\u0/u1/X [33]),
        .I3(\u0/u1/X [32]),
        .I4(\u0/u1/X [36]),
        .I5(\u0/u1/X [31]),
        .O(\u0/out1 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__90
       (.I0(\u0/u11/X [11]),
        .I1(\u0/u11/X [10]),
        .I2(\u0/u11/X [9]),
        .I3(\u0/u11/X [8]),
        .I4(\u0/u11/X [12]),
        .I5(\u0/u11/X [7]),
        .O(\u0/out11 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__91
       (.I0(\u0/u11/X [47]),
        .I1(\u0/u11/X [46]),
        .I2(\u0/u11/X [45]),
        .I3(\u0/u11/X [44]),
        .I4(\u0/u11/X [48]),
        .I5(\u0/u11/X [43]),
        .O(\u0/out11 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB64A99D24B39E827)) 
    g0_b2__92
       (.I0(\u0/u11/X [23]),
        .I1(\u0/u11/X [22]),
        .I2(\u0/u11/X [21]),
        .I3(\u0/u11/X [20]),
        .I4(\u0/u11/X [24]),
        .I5(\u0/u11/X [19]),
        .O(\u0/out11 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h63AC9D6185795A96)) 
    g0_b2__93
       (.I0(\u0/u11/X [29]),
        .I1(\u0/u11/X [28]),
        .I2(\u0/u11/X [27]),
        .I3(\u0/u11/X [26]),
        .I4(\u0/u11/X [30]),
        .I5(\u0/u11/X [25]),
        .O(\u0/out11 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC9934B35265E9C27)) 
    g0_b2__94
       (.I0(\u0/u11/X [5]),
        .I1(\u0/u11/X [4]),
        .I2(\u0/u11/X [3]),
        .I3(\u0/u11/X [2]),
        .I4(\u0/u11/X [6]),
        .I5(\u0/u11/X [1]),
        .O(\u0/out11 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9AA526DAAD195A99)) 
    g0_b2__95
       (.I0(\u0/u12/X [41]),
        .I1(\u0/u12/X [40]),
        .I2(\u0/u12/X [39]),
        .I3(\u0/u12/X [38]),
        .I4(\u0/u12/X [42]),
        .I5(\u0/u12/X [37]),
        .O(\u0/out12 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA794D8275C632ED8)) 
    g0_b2__96
       (.I0(\u0/u12/X [17]),
        .I1(\u0/u12/X [16]),
        .I2(\u0/u12/X [15]),
        .I3(\u0/u12/X [14]),
        .I4(\u0/u12/X [18]),
        .I5(\u0/u12/X [13]),
        .O(\u0/out12 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A69A54E0DB67A49)) 
    g0_b2__97
       (.I0(\u0/u12/X [35]),
        .I1(\u0/u12/X [34]),
        .I2(\u0/u12/X [33]),
        .I3(\u0/u12/X [32]),
        .I4(\u0/u12/X [36]),
        .I5(\u0/u12/X [31]),
        .O(\u0/out12 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6E618D66919E5A99)) 
    g0_b2__98
       (.I0(\u0/u12/X [11]),
        .I1(\u0/u12/X [10]),
        .I2(\u0/u12/X [9]),
        .I3(\u0/u12/X [8]),
        .I4(\u0/u12/X [12]),
        .I5(\u0/u12/X [7]),
        .O(\u0/out12 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h639C5A6527C6D839)) 
    g0_b2__99
       (.I0(\u0/u12/X [47]),
        .I1(\u0/u12/X [46]),
        .I2(\u0/u12/X [45]),
        .I3(\u0/u12/X [44]),
        .I4(\u0/u12/X [48]),
        .I5(\u0/u12/X [43]),
        .O(\u0/out12 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3
       (.I0(\u0/u0/X [41]),
        .I1(\u0/u0/X [40]),
        .I2(\u0/u0/X [39]),
        .I3(\u0/u0/X [38]),
        .I4(\u0/u0/X [42]),
        .I5(\u0/u0/X [37]),
        .O(\u0/out0 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__0
       (.I0(\u0/u0/X [17]),
        .I1(\u0/u0/X [16]),
        .I2(\u0/u0/X [15]),
        .I3(\u0/u0/X [14]),
        .I4(\u0/u0/X [18]),
        .I5(\u0/u0/X [13]),
        .O(\u0/out0 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__1
       (.I0(\u0/u0/X [35]),
        .I1(\u0/u0/X [34]),
        .I2(\u0/u0/X [33]),
        .I3(\u0/u0/X [32]),
        .I4(\u0/u0/X [36]),
        .I5(\u0/u0/X [31]),
        .O(\u0/out0 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__10
       (.I0(\u0/u1/X [11]),
        .I1(\u0/u1/X [10]),
        .I2(\u0/u1/X [9]),
        .I3(\u0/u1/X [8]),
        .I4(\u0/u1/X [12]),
        .I5(\u0/u1/X [7]),
        .O(\u0/out1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__100
       (.I0(\u0/u12/X [23]),
        .I1(\u0/u12/X [22]),
        .I2(\u0/u12/X [21]),
        .I3(\u0/u12/X [20]),
        .I4(\u0/u12/X [24]),
        .I5(\u0/u12/X [19]),
        .O(\u0/out12 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__101
       (.I0(\u0/u12/X [29]),
        .I1(\u0/u12/X [28]),
        .I2(\u0/u12/X [27]),
        .I3(\u0/u12/X [26]),
        .I4(\u0/u12/X [30]),
        .I5(\u0/u12/X [25]),
        .O(\u0/out12 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__102
       (.I0(\u0/u12/X [5]),
        .I1(\u0/u12/X [4]),
        .I2(\u0/u12/X [3]),
        .I3(\u0/u12/X [2]),
        .I4(\u0/u12/X [6]),
        .I5(\u0/u12/X [1]),
        .O(\u0/out12 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__103
       (.I0(\u0/u13/X [41]),
        .I1(\u0/u13/X [40]),
        .I2(\u0/u13/X [39]),
        .I3(\u0/u13/X [38]),
        .I4(\u0/u13/X [42]),
        .I5(\u0/u13/X [37]),
        .O(\u0/out13 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__104
       (.I0(\u0/u13/X [17]),
        .I1(\u0/u13/X [16]),
        .I2(\u0/u13/X [15]),
        .I3(\u0/u13/X [14]),
        .I4(\u0/u13/X [18]),
        .I5(\u0/u13/X [13]),
        .O(\u0/out13 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__105
       (.I0(\u0/u13/X [35]),
        .I1(\u0/u13/X [34]),
        .I2(\u0/u13/X [33]),
        .I3(\u0/u13/X [32]),
        .I4(\u0/u13/X [36]),
        .I5(\u0/u13/X [31]),
        .O(\u0/out13 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__106
       (.I0(\u0/u13/X [11]),
        .I1(\u0/u13/X [10]),
        .I2(\u0/u13/X [9]),
        .I3(\u0/u13/X [8]),
        .I4(\u0/u13/X [12]),
        .I5(\u0/u13/X [7]),
        .O(\u0/out13 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__107
       (.I0(\u0/u13/X [47]),
        .I1(\u0/u13/X [46]),
        .I2(\u0/u13/X [45]),
        .I3(\u0/u13/X [44]),
        .I4(\u0/u13/X [48]),
        .I5(\u0/u13/X [43]),
        .O(\u0/out13 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__108
       (.I0(\u0/u13/X [23]),
        .I1(\u0/u13/X [22]),
        .I2(\u0/u13/X [21]),
        .I3(\u0/u13/X [20]),
        .I4(\u0/u13/X [24]),
        .I5(\u0/u13/X [19]),
        .O(\u0/out13 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__109
       (.I0(\u0/u13/X [29]),
        .I1(\u0/u13/X [28]),
        .I2(\u0/u13/X [27]),
        .I3(\u0/u13/X [26]),
        .I4(\u0/u13/X [30]),
        .I5(\u0/u13/X [25]),
        .O(\u0/out13 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__11
       (.I0(\u0/u1/X [47]),
        .I1(\u0/u1/X [46]),
        .I2(\u0/u1/X [45]),
        .I3(\u0/u1/X [44]),
        .I4(\u0/u1/X [48]),
        .I5(\u0/u1/X [43]),
        .O(\u0/out1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__110
       (.I0(\u0/u13/X [5]),
        .I1(\u0/u13/X [4]),
        .I2(\u0/u13/X [3]),
        .I3(\u0/u13/X [2]),
        .I4(\u0/u13/X [6]),
        .I5(\u0/u13/X [1]),
        .O(\u0/out13 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__111
       (.I0(\u0/u14/X [41]),
        .I1(\u0/u14/X [40]),
        .I2(\u0/u14/X [39]),
        .I3(\u0/u14/X [38]),
        .I4(\u0/u14/X [42]),
        .I5(\u0/u14/X [37]),
        .O(\u0/out14 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__112
       (.I0(\u0/u14/X [17]),
        .I1(\u0/u14/X [16]),
        .I2(\u0/u14/X [15]),
        .I3(\u0/u14/X [14]),
        .I4(\u0/u14/X [18]),
        .I5(\u0/u14/X [13]),
        .O(\u0/out14 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__113
       (.I0(\u0/u14/X [35]),
        .I1(\u0/u14/X [34]),
        .I2(\u0/u14/X [33]),
        .I3(\u0/u14/X [32]),
        .I4(\u0/u14/X [36]),
        .I5(\u0/u14/X [31]),
        .O(\u0/out14 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__114
       (.I0(\u0/u14/X [11]),
        .I1(\u0/u14/X [10]),
        .I2(\u0/u14/X [9]),
        .I3(\u0/u14/X [8]),
        .I4(\u0/u14/X [12]),
        .I5(\u0/u14/X [7]),
        .O(\u0/out14 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__115
       (.I0(\u0/u14/X [47]),
        .I1(\u0/u14/X [46]),
        .I2(\u0/u14/X [45]),
        .I3(\u0/u14/X [44]),
        .I4(\u0/u14/X [48]),
        .I5(\u0/u14/X [43]),
        .O(\u0/out14 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__116
       (.I0(\u0/u14/X [23]),
        .I1(\u0/u14/X [22]),
        .I2(\u0/u14/X [21]),
        .I3(\u0/u14/X [20]),
        .I4(\u0/u14/X [24]),
        .I5(\u0/u14/X [19]),
        .O(\u0/out14 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__117
       (.I0(\u0/u14/X [29]),
        .I1(\u0/u14/X [28]),
        .I2(\u0/u14/X [27]),
        .I3(\u0/u14/X [26]),
        .I4(\u0/u14/X [30]),
        .I5(\u0/u14/X [25]),
        .O(\u0/out14 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__118
       (.I0(\u0/u14/X [5]),
        .I1(\u0/u14/X [4]),
        .I2(\u0/u14/X [3]),
        .I3(\u0/u14/X [2]),
        .I4(\u0/u14/X [6]),
        .I5(\u0/u14/X [1]),
        .O(\u0/out14 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__119
       (.I0(\u0/u15/X [41]),
        .I1(\u0/u15/X [40]),
        .I2(\u0/u15/X [39]),
        .I3(\u0/u15/X [38]),
        .I4(\u0/u15/X [42]),
        .I5(\u0/u15/X [37]),
        .O(\u0/out15 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__12
       (.I0(\u0/u1/X [23]),
        .I1(\u0/u1/X [22]),
        .I2(\u0/u1/X [21]),
        .I3(\u0/u1/X [20]),
        .I4(\u0/u1/X [24]),
        .I5(\u0/u1/X [19]),
        .O(\u0/out1 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__120
       (.I0(\u0/u15/X [17]),
        .I1(\u0/u15/X [16]),
        .I2(\u0/u15/X [15]),
        .I3(\u0/u15/X [14]),
        .I4(\u0/u15/X [18]),
        .I5(\u0/u15/X [13]),
        .O(\u0/out15 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__121
       (.I0(\u0/u15/X [35]),
        .I1(\u0/u15/X [34]),
        .I2(\u0/u15/X [33]),
        .I3(\u0/u15/X [32]),
        .I4(\u0/u15/X [36]),
        .I5(\u0/u15/X [31]),
        .O(\u0/out15 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__122
       (.I0(\u0/u15/X [11]),
        .I1(\u0/u15/X [10]),
        .I2(\u0/u15/X [9]),
        .I3(\u0/u15/X [8]),
        .I4(\u0/u15/X [12]),
        .I5(\u0/u15/X [7]),
        .O(\u0/out15 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__123
       (.I0(\u0/u15/X [47]),
        .I1(\u0/u15/X [46]),
        .I2(\u0/u15/X [45]),
        .I3(\u0/u15/X [44]),
        .I4(\u0/u15/X [48]),
        .I5(\u0/u15/X [43]),
        .O(\u0/out15 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__124
       (.I0(\u0/u15/X [23]),
        .I1(\u0/u15/X [22]),
        .I2(\u0/u15/X [21]),
        .I3(\u0/u15/X [20]),
        .I4(\u0/u15/X [24]),
        .I5(\u0/u15/X [19]),
        .O(\u0/out15 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__125
       (.I0(\u0/u15/X [29]),
        .I1(\u0/u15/X [28]),
        .I2(\u0/u15/X [27]),
        .I3(\u0/u15/X [26]),
        .I4(\u0/u15/X [30]),
        .I5(\u0/u15/X [25]),
        .O(\u0/out15 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__126
       (.I0(\u0/u15/X [5]),
        .I1(\u0/u15/X [4]),
        .I2(\u0/u15/X [3]),
        .I3(\u0/u15/X [2]),
        .I4(\u0/u15/X [6]),
        .I5(\u0/u15/X [1]),
        .O(\u0/out15 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__127
       (.I0(\u1/u0/X [41]),
        .I1(\u1/u0/X [40]),
        .I2(\u1/u0/X [39]),
        .I3(\u1/u0/X [38]),
        .I4(\u1/u0/X [42]),
        .I5(\u1/u0/X [37]),
        .O(\u1/out0 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__128
       (.I0(\u1/u0/X [17]),
        .I1(\u1/u0/X [16]),
        .I2(\u1/u0/X [15]),
        .I3(\u1/u0/X [14]),
        .I4(\u1/u0/X [18]),
        .I5(\u1/u0/X [13]),
        .O(\u1/out0 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__129
       (.I0(\u1/u0/X [35]),
        .I1(\u1/u0/X [34]),
        .I2(\u1/u0/X [33]),
        .I3(\u1/u0/X [32]),
        .I4(\u1/u0/X [36]),
        .I5(\u1/u0/X [31]),
        .O(\u1/out0 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__13
       (.I0(\u0/u1/X [29]),
        .I1(\u0/u1/X [28]),
        .I2(\u0/u1/X [27]),
        .I3(\u0/u1/X [26]),
        .I4(\u0/u1/X [30]),
        .I5(\u0/u1/X [25]),
        .O(\u0/out1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__130
       (.I0(\u1/u0/X [11]),
        .I1(\u1/u0/X [10]),
        .I2(\u1/u0/X [9]),
        .I3(\u1/u0/X [8]),
        .I4(\u1/u0/X [12]),
        .I5(\u1/u0/X [7]),
        .O(\u1/out0 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__131
       (.I0(\u1/u0/X [47]),
        .I1(\u1/u0/X [46]),
        .I2(\u1/u0/X [45]),
        .I3(\u1/u0/X [44]),
        .I4(\u1/u0/X [48]),
        .I5(\u1/u0/X [43]),
        .O(\u1/out0 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__132
       (.I0(\u1/u0/X [23]),
        .I1(\u1/u0/X [22]),
        .I2(\u1/u0/X [21]),
        .I3(\u1/u0/X [20]),
        .I4(\u1/u0/X [24]),
        .I5(\u1/u0/X [19]),
        .O(\u1/out0 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__133
       (.I0(\u1/u0/X [29]),
        .I1(\u1/u0/X [28]),
        .I2(\u1/u0/X [27]),
        .I3(\u1/u0/X [26]),
        .I4(\u1/u0/X [30]),
        .I5(\u1/u0/X [25]),
        .O(\u1/out0 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__134
       (.I0(\u1/u0/X [5]),
        .I1(\u1/u0/X [4]),
        .I2(\u1/u0/X [3]),
        .I3(\u1/u0/X [2]),
        .I4(\u1/u0/X [6]),
        .I5(\u1/u0/X [1]),
        .O(\u1/out0 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__135
       (.I0(\u1/u1/X [41]),
        .I1(\u1/u1/X [40]),
        .I2(\u1/u1/X [39]),
        .I3(\u1/u1/X [38]),
        .I4(\u1/u1/X [42]),
        .I5(\u1/u1/X [37]),
        .O(\u1/out1 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__136
       (.I0(\u1/u1/X [17]),
        .I1(\u1/u1/X [16]),
        .I2(\u1/u1/X [15]),
        .I3(\u1/u1/X [14]),
        .I4(\u1/u1/X [18]),
        .I5(\u1/u1/X [13]),
        .O(\u1/out1 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__137
       (.I0(\u1/u1/X [35]),
        .I1(\u1/u1/X [34]),
        .I2(\u1/u1/X [33]),
        .I3(\u1/u1/X [32]),
        .I4(\u1/u1/X [36]),
        .I5(\u1/u1/X [31]),
        .O(\u1/out1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__138
       (.I0(\u1/u1/X [11]),
        .I1(\u1/u1/X [10]),
        .I2(\u1/u1/X [9]),
        .I3(\u1/u1/X [8]),
        .I4(\u1/u1/X [12]),
        .I5(\u1/u1/X [7]),
        .O(\u1/out1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__139
       (.I0(\u1/u1/X [47]),
        .I1(\u1/u1/X [46]),
        .I2(\u1/u1/X [45]),
        .I3(\u1/u1/X [44]),
        .I4(\u1/u1/X [48]),
        .I5(\u1/u1/X [43]),
        .O(\u1/out1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__14
       (.I0(\u0/u1/X [5]),
        .I1(\u0/u1/X [4]),
        .I2(\u0/u1/X [3]),
        .I3(\u0/u1/X [2]),
        .I4(\u0/u1/X [6]),
        .I5(\u0/u1/X [1]),
        .O(\u0/out1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__140
       (.I0(\u1/u1/X [23]),
        .I1(\u1/u1/X [22]),
        .I2(\u1/u1/X [21]),
        .I3(\u1/u1/X [20]),
        .I4(\u1/u1/X [24]),
        .I5(\u1/u1/X [19]),
        .O(\u1/out1 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__141
       (.I0(\u1/u1/X [29]),
        .I1(\u1/u1/X [28]),
        .I2(\u1/u1/X [27]),
        .I3(\u1/u1/X [26]),
        .I4(\u1/u1/X [30]),
        .I5(\u1/u1/X [25]),
        .O(\u1/out1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__142
       (.I0(\u1/u1/X [5]),
        .I1(\u1/u1/X [4]),
        .I2(\u1/u1/X [3]),
        .I3(\u1/u1/X [2]),
        .I4(\u1/u1/X [6]),
        .I5(\u1/u1/X [1]),
        .O(\u1/out1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__143
       (.I0(\u1/u2/X [41]),
        .I1(\u1/u2/X [40]),
        .I2(\u1/u2/X [39]),
        .I3(\u1/u2/X [38]),
        .I4(\u1/u2/X [42]),
        .I5(\u1/u2/X [37]),
        .O(\u1/out2 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__144
       (.I0(\u1/u2/X [17]),
        .I1(\u1/u2/X [16]),
        .I2(\u1/u2/X [15]),
        .I3(\u1/u2/X [14]),
        .I4(\u1/u2/X [18]),
        .I5(\u1/u2/X [13]),
        .O(\u1/out2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__145
       (.I0(\u1/u2/X [35]),
        .I1(\u1/u2/X [34]),
        .I2(\u1/u2/X [33]),
        .I3(\u1/u2/X [32]),
        .I4(\u1/u2/X [36]),
        .I5(\u1/u2/X [31]),
        .O(\u1/out2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__146
       (.I0(\u1/u2/X [11]),
        .I1(\u1/u2/X [10]),
        .I2(\u1/u2/X [9]),
        .I3(\u1/u2/X [8]),
        .I4(\u1/u2/X [12]),
        .I5(\u1/u2/X [7]),
        .O(\u1/out2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__147
       (.I0(\u1/u2/X [47]),
        .I1(\u1/u2/X [46]),
        .I2(\u1/u2/X [45]),
        .I3(\u1/u2/X [44]),
        .I4(\u1/u2/X [48]),
        .I5(\u1/u2/X [43]),
        .O(\u1/out2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__148
       (.I0(\u1/u2/X [23]),
        .I1(\u1/u2/X [22]),
        .I2(\u1/u2/X [21]),
        .I3(\u1/u2/X [20]),
        .I4(\u1/u2/X [24]),
        .I5(\u1/u2/X [19]),
        .O(\u1/out2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__149
       (.I0(\u1/u2/X [29]),
        .I1(\u1/u2/X [28]),
        .I2(\u1/u2/X [27]),
        .I3(\u1/u2/X [26]),
        .I4(\u1/u2/X [30]),
        .I5(\u1/u2/X [25]),
        .O(\u1/out2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__15
       (.I0(\u0/u2/X [41]),
        .I1(\u0/u2/X [40]),
        .I2(\u0/u2/X [39]),
        .I3(\u0/u2/X [38]),
        .I4(\u0/u2/X [42]),
        .I5(\u0/u2/X [37]),
        .O(\u0/out2 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__150
       (.I0(\u1/u2/X [5]),
        .I1(\u1/u2/X [4]),
        .I2(\u1/u2/X [3]),
        .I3(\u1/u2/X [2]),
        .I4(\u1/u2/X [6]),
        .I5(\u1/u2/X [1]),
        .O(\u1/out2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__151
       (.I0(\u1/u3/X [41]),
        .I1(\u1/u3/X [40]),
        .I2(\u1/u3/X [39]),
        .I3(\u1/u3/X [38]),
        .I4(\u1/u3/X [42]),
        .I5(\u1/u3/X [37]),
        .O(\u1/out3 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__152
       (.I0(\u1/u3/X [17]),
        .I1(\u1/u3/X [16]),
        .I2(\u1/u3/X [15]),
        .I3(\u1/u3/X [14]),
        .I4(\u1/u3/X [18]),
        .I5(\u1/u3/X [13]),
        .O(\u1/out3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__153
       (.I0(\u1/u3/X [35]),
        .I1(\u1/u3/X [34]),
        .I2(\u1/u3/X [33]),
        .I3(\u1/u3/X [32]),
        .I4(\u1/u3/X [36]),
        .I5(\u1/u3/X [31]),
        .O(\u1/out3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__154
       (.I0(\u1/u3/X [11]),
        .I1(\u1/u3/X [10]),
        .I2(\u1/u3/X [9]),
        .I3(\u1/u3/X [8]),
        .I4(\u1/u3/X [12]),
        .I5(\u1/u3/X [7]),
        .O(\u1/out3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__155
       (.I0(\u1/u3/X [47]),
        .I1(\u1/u3/X [46]),
        .I2(\u1/u3/X [45]),
        .I3(\u1/u3/X [44]),
        .I4(\u1/u3/X [48]),
        .I5(\u1/u3/X [43]),
        .O(\u1/out3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__156
       (.I0(\u1/u3/X [23]),
        .I1(\u1/u3/X [22]),
        .I2(\u1/u3/X [21]),
        .I3(\u1/u3/X [20]),
        .I4(\u1/u3/X [24]),
        .I5(\u1/u3/X [19]),
        .O(\u1/out3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__157
       (.I0(\u1/u3/X [29]),
        .I1(\u1/u3/X [28]),
        .I2(\u1/u3/X [27]),
        .I3(\u1/u3/X [26]),
        .I4(\u1/u3/X [30]),
        .I5(\u1/u3/X [25]),
        .O(\u1/out3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__158
       (.I0(\u1/u3/X [5]),
        .I1(\u1/u3/X [4]),
        .I2(\u1/u3/X [3]),
        .I3(\u1/u3/X [2]),
        .I4(\u1/u3/X [6]),
        .I5(\u1/u3/X [1]),
        .O(\u1/out3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__159
       (.I0(\u1/u4/X [41]),
        .I1(\u1/u4/X [40]),
        .I2(\u1/u4/X [39]),
        .I3(\u1/u4/X [38]),
        .I4(\u1/u4/X [42]),
        .I5(\u1/u4/X [37]),
        .O(\u1/out4 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__16
       (.I0(\u0/u2/X [17]),
        .I1(\u0/u2/X [16]),
        .I2(\u0/u2/X [15]),
        .I3(\u0/u2/X [14]),
        .I4(\u0/u2/X [18]),
        .I5(\u0/u2/X [13]),
        .O(\u0/out2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__160
       (.I0(\u1/u4/X [17]),
        .I1(\u1/u4/X [16]),
        .I2(\u1/u4/X [15]),
        .I3(\u1/u4/X [14]),
        .I4(\u1/u4/X [18]),
        .I5(\u1/u4/X [13]),
        .O(\u1/out4 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__161
       (.I0(\u1/u4/X [35]),
        .I1(\u1/u4/X [34]),
        .I2(\u1/u4/X [33]),
        .I3(\u1/u4/X [32]),
        .I4(\u1/u4/X [36]),
        .I5(\u1/u4/X [31]),
        .O(\u1/out4 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__162
       (.I0(\u1/u4/X [11]),
        .I1(\u1/u4/X [10]),
        .I2(\u1/u4/X [9]),
        .I3(\u1/u4/X [8]),
        .I4(\u1/u4/X [12]),
        .I5(\u1/u4/X [7]),
        .O(\u1/out4 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__163
       (.I0(\u1/u4/X [47]),
        .I1(\u1/u4/X [46]),
        .I2(\u1/u4/X [45]),
        .I3(\u1/u4/X [44]),
        .I4(\u1/u4/X [48]),
        .I5(\u1/u4/X [43]),
        .O(\u1/out4 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__164
       (.I0(\u1/u4/X [23]),
        .I1(\u1/u4/X [22]),
        .I2(\u1/u4/X [21]),
        .I3(\u1/u4/X [20]),
        .I4(\u1/u4/X [24]),
        .I5(\u1/u4/X [19]),
        .O(\u1/out4 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__165
       (.I0(\u1/u4/X [29]),
        .I1(\u1/u4/X [28]),
        .I2(\u1/u4/X [27]),
        .I3(\u1/u4/X [26]),
        .I4(\u1/u4/X [30]),
        .I5(\u1/u4/X [25]),
        .O(\u1/out4 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__166
       (.I0(\u1/u4/X [5]),
        .I1(\u1/u4/X [4]),
        .I2(\u1/u4/X [3]),
        .I3(\u1/u4/X [2]),
        .I4(\u1/u4/X [6]),
        .I5(\u1/u4/X [1]),
        .O(\u1/out4 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__167
       (.I0(\u1/u5/X [41]),
        .I1(\u1/u5/X [40]),
        .I2(\u1/u5/X [39]),
        .I3(\u1/u5/X [38]),
        .I4(\u1/u5/X [42]),
        .I5(\u1/u5/X [37]),
        .O(\u1/out5 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__168
       (.I0(\u1/u5/X [17]),
        .I1(\u1/u5/X [16]),
        .I2(\u1/u5/X [15]),
        .I3(\u1/u5/X [14]),
        .I4(\u1/u5/X [18]),
        .I5(\u1/u5/X [13]),
        .O(\u1/out5 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__169
       (.I0(\u1/u5/X [35]),
        .I1(\u1/u5/X [34]),
        .I2(\u1/u5/X [33]),
        .I3(\u1/u5/X [32]),
        .I4(\u1/u5/X [36]),
        .I5(\u1/u5/X [31]),
        .O(\u1/out5 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__17
       (.I0(\u0/u2/X [35]),
        .I1(\u0/u2/X [34]),
        .I2(\u0/u2/X [33]),
        .I3(\u0/u2/X [32]),
        .I4(\u0/u2/X [36]),
        .I5(\u0/u2/X [31]),
        .O(\u0/out2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__170
       (.I0(\u1/u5/X [11]),
        .I1(\u1/u5/X [10]),
        .I2(\u1/u5/X [9]),
        .I3(\u1/u5/X [8]),
        .I4(\u1/u5/X [12]),
        .I5(\u1/u5/X [7]),
        .O(\u1/out5 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__171
       (.I0(\u1/u5/X [47]),
        .I1(\u1/u5/X [46]),
        .I2(\u1/u5/X [45]),
        .I3(\u1/u5/X [44]),
        .I4(\u1/u5/X [48]),
        .I5(\u1/u5/X [43]),
        .O(\u1/out5 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__172
       (.I0(\u1/u5/X [23]),
        .I1(\u1/u5/X [22]),
        .I2(\u1/u5/X [21]),
        .I3(\u1/u5/X [20]),
        .I4(\u1/u5/X [24]),
        .I5(\u1/u5/X [19]),
        .O(\u1/out5 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__173
       (.I0(\u1/u5/X [29]),
        .I1(\u1/u5/X [28]),
        .I2(\u1/u5/X [27]),
        .I3(\u1/u5/X [26]),
        .I4(\u1/u5/X [30]),
        .I5(\u1/u5/X [25]),
        .O(\u1/out5 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__174
       (.I0(\u1/u5/X [5]),
        .I1(\u1/u5/X [4]),
        .I2(\u1/u5/X [3]),
        .I3(\u1/u5/X [2]),
        .I4(\u1/u5/X [6]),
        .I5(\u1/u5/X [1]),
        .O(\u1/out5 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__175
       (.I0(\u1/u6/X [41]),
        .I1(\u1/u6/X [40]),
        .I2(\u1/u6/X [39]),
        .I3(\u1/u6/X [38]),
        .I4(\u1/u6/X [42]),
        .I5(\u1/u6/X [37]),
        .O(\u1/out6 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__176
       (.I0(\u1/u6/X [17]),
        .I1(\u1/u6/X [16]),
        .I2(\u1/u6/X [15]),
        .I3(\u1/u6/X [14]),
        .I4(\u1/u6/X [18]),
        .I5(\u1/u6/X [13]),
        .O(\u1/out6 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__177
       (.I0(\u1/u6/X [35]),
        .I1(\u1/u6/X [34]),
        .I2(\u1/u6/X [33]),
        .I3(\u1/u6/X [32]),
        .I4(\u1/u6/X [36]),
        .I5(\u1/u6/X [31]),
        .O(\u1/out6 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__178
       (.I0(\u1/u6/X [11]),
        .I1(\u1/u6/X [10]),
        .I2(\u1/u6/X [9]),
        .I3(\u1/u6/X [8]),
        .I4(\u1/u6/X [12]),
        .I5(\u1/u6/X [7]),
        .O(\u1/out6 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__179
       (.I0(\u1/u6/X [47]),
        .I1(\u1/u6/X [46]),
        .I2(\u1/u6/X [45]),
        .I3(\u1/u6/X [44]),
        .I4(\u1/u6/X [48]),
        .I5(\u1/u6/X [43]),
        .O(\u1/out6 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__18
       (.I0(\u0/u2/X [11]),
        .I1(\u0/u2/X [10]),
        .I2(\u0/u2/X [9]),
        .I3(\u0/u2/X [8]),
        .I4(\u0/u2/X [12]),
        .I5(\u0/u2/X [7]),
        .O(\u0/out2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__180
       (.I0(\u1/u6/X [23]),
        .I1(\u1/u6/X [22]),
        .I2(\u1/u6/X [21]),
        .I3(\u1/u6/X [20]),
        .I4(\u1/u6/X [24]),
        .I5(\u1/u6/X [19]),
        .O(\u1/out6 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__181
       (.I0(\u1/u6/X [29]),
        .I1(\u1/u6/X [28]),
        .I2(\u1/u6/X [27]),
        .I3(\u1/u6/X [26]),
        .I4(\u1/u6/X [30]),
        .I5(\u1/u6/X [25]),
        .O(\u1/out6 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__182
       (.I0(\u1/u6/X [5]),
        .I1(\u1/u6/X [4]),
        .I2(\u1/u6/X [3]),
        .I3(\u1/u6/X [2]),
        .I4(\u1/u6/X [6]),
        .I5(\u1/u6/X [1]),
        .O(\u1/out6 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__183
       (.I0(\u1/u7/X [41]),
        .I1(\u1/u7/X [40]),
        .I2(\u1/u7/X [39]),
        .I3(\u1/u7/X [38]),
        .I4(\u1/u7/X [42]),
        .I5(\u1/u7/X [37]),
        .O(\u1/out7 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__184
       (.I0(\u1/u7/X [17]),
        .I1(\u1/u7/X [16]),
        .I2(\u1/u7/X [15]),
        .I3(\u1/u7/X [14]),
        .I4(\u1/u7/X [18]),
        .I5(\u1/u7/X [13]),
        .O(\u1/out7 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__185
       (.I0(\u1/u7/X [35]),
        .I1(\u1/u7/X [34]),
        .I2(\u1/u7/X [33]),
        .I3(\u1/u7/X [32]),
        .I4(\u1/u7/X [36]),
        .I5(\u1/u7/X [31]),
        .O(\u1/out7 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__186
       (.I0(\u1/u7/X [11]),
        .I1(\u1/u7/X [10]),
        .I2(\u1/u7/X [9]),
        .I3(\u1/u7/X [8]),
        .I4(\u1/u7/X [12]),
        .I5(\u1/u7/X [7]),
        .O(\u1/out7 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__187
       (.I0(\u1/u7/X [47]),
        .I1(\u1/u7/X [46]),
        .I2(\u1/u7/X [45]),
        .I3(\u1/u7/X [44]),
        .I4(\u1/u7/X [48]),
        .I5(\u1/u7/X [43]),
        .O(\u1/out7 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__188
       (.I0(\u1/u7/X [23]),
        .I1(\u1/u7/X [22]),
        .I2(\u1/u7/X [21]),
        .I3(\u1/u7/X [20]),
        .I4(\u1/u7/X [24]),
        .I5(\u1/u7/X [19]),
        .O(\u1/out7 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__189
       (.I0(\u1/u7/X [29]),
        .I1(\u1/u7/X [28]),
        .I2(\u1/u7/X [27]),
        .I3(\u1/u7/X [26]),
        .I4(\u1/u7/X [30]),
        .I5(\u1/u7/X [25]),
        .O(\u1/out7 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__19
       (.I0(\u0/u2/X [47]),
        .I1(\u0/u2/X [46]),
        .I2(\u0/u2/X [45]),
        .I3(\u0/u2/X [44]),
        .I4(\u0/u2/X [48]),
        .I5(\u0/u2/X [43]),
        .O(\u0/out2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__190
       (.I0(\u1/u7/X [5]),
        .I1(\u1/u7/X [4]),
        .I2(\u1/u7/X [3]),
        .I3(\u1/u7/X [2]),
        .I4(\u1/u7/X [6]),
        .I5(\u1/u7/X [1]),
        .O(\u1/out7 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__191
       (.I0(\u1/u8/X [41]),
        .I1(\u1/u8/X [40]),
        .I2(\u1/u8/X [39]),
        .I3(\u1/u8/X [38]),
        .I4(\u1/u8/X [42]),
        .I5(\u1/u8/X [37]),
        .O(\u1/out8 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__192
       (.I0(\u1/u8/X [17]),
        .I1(\u1/u8/X [16]),
        .I2(\u1/u8/X [15]),
        .I3(\u1/u8/X [14]),
        .I4(\u1/u8/X [18]),
        .I5(\u1/u8/X [13]),
        .O(\u1/out8 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__193
       (.I0(\u1/u8/X [35]),
        .I1(\u1/u8/X [34]),
        .I2(\u1/u8/X [33]),
        .I3(\u1/u8/X [32]),
        .I4(\u1/u8/X [36]),
        .I5(\u1/u8/X [31]),
        .O(\u1/out8 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__194
       (.I0(\u1/u8/X [11]),
        .I1(\u1/u8/X [10]),
        .I2(\u1/u8/X [9]),
        .I3(\u1/u8/X [8]),
        .I4(\u1/u8/X [12]),
        .I5(\u1/u8/X [7]),
        .O(\u1/out8 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__195
       (.I0(\u1/u8/X [47]),
        .I1(\u1/u8/X [46]),
        .I2(\u1/u8/X [45]),
        .I3(\u1/u8/X [44]),
        .I4(\u1/u8/X [48]),
        .I5(\u1/u8/X [43]),
        .O(\u1/out8 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__196
       (.I0(\u1/u8/X [23]),
        .I1(\u1/u8/X [22]),
        .I2(\u1/u8/X [21]),
        .I3(\u1/u8/X [20]),
        .I4(\u1/u8/X [24]),
        .I5(\u1/u8/X [19]),
        .O(\u1/out8 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__197
       (.I0(\u1/u8/X [29]),
        .I1(\u1/u8/X [28]),
        .I2(\u1/u8/X [27]),
        .I3(\u1/u8/X [26]),
        .I4(\u1/u8/X [30]),
        .I5(\u1/u8/X [25]),
        .O(\u1/out8 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__198
       (.I0(\u1/u8/X [5]),
        .I1(\u1/u8/X [4]),
        .I2(\u1/u8/X [3]),
        .I3(\u1/u8/X [2]),
        .I4(\u1/u8/X [6]),
        .I5(\u1/u8/X [1]),
        .O(\u1/out8 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__199
       (.I0(\u1/u9/X [41]),
        .I1(\u1/u9/X [40]),
        .I2(\u1/u9/X [39]),
        .I3(\u1/u9/X [38]),
        .I4(\u1/u9/X [42]),
        .I5(\u1/u9/X [37]),
        .O(\u1/out9 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__2
       (.I0(\u0/u0/X [11]),
        .I1(\u0/u0/X [10]),
        .I2(\u0/u0/X [9]),
        .I3(\u0/u0/X [8]),
        .I4(\u0/u0/X [12]),
        .I5(\u0/u0/X [7]),
        .O(\u0/out0 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__20
       (.I0(\u0/u2/X [23]),
        .I1(\u0/u2/X [22]),
        .I2(\u0/u2/X [21]),
        .I3(\u0/u2/X [20]),
        .I4(\u0/u2/X [24]),
        .I5(\u0/u2/X [19]),
        .O(\u0/out2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__200
       (.I0(\u1/u9/X [17]),
        .I1(\u1/u9/X [16]),
        .I2(\u1/u9/X [15]),
        .I3(\u1/u9/X [14]),
        .I4(\u1/u9/X [18]),
        .I5(\u1/u9/X [13]),
        .O(\u1/out9 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__201
       (.I0(\u1/u9/X [35]),
        .I1(\u1/u9/X [34]),
        .I2(\u1/u9/X [33]),
        .I3(\u1/u9/X [32]),
        .I4(\u1/u9/X [36]),
        .I5(\u1/u9/X [31]),
        .O(\u1/out9 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__202
       (.I0(\u1/u9/X [11]),
        .I1(\u1/u9/X [10]),
        .I2(\u1/u9/X [9]),
        .I3(\u1/u9/X [8]),
        .I4(\u1/u9/X [12]),
        .I5(\u1/u9/X [7]),
        .O(\u1/out9 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__203
       (.I0(\u1/u9/X [47]),
        .I1(\u1/u9/X [46]),
        .I2(\u1/u9/X [45]),
        .I3(\u1/u9/X [44]),
        .I4(\u1/u9/X [48]),
        .I5(\u1/u9/X [43]),
        .O(\u1/out9 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__204
       (.I0(\u1/u9/X [23]),
        .I1(\u1/u9/X [22]),
        .I2(\u1/u9/X [21]),
        .I3(\u1/u9/X [20]),
        .I4(\u1/u9/X [24]),
        .I5(\u1/u9/X [19]),
        .O(\u1/out9 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__205
       (.I0(\u1/u9/X [29]),
        .I1(\u1/u9/X [28]),
        .I2(\u1/u9/X [27]),
        .I3(\u1/u9/X [26]),
        .I4(\u1/u9/X [30]),
        .I5(\u1/u9/X [25]),
        .O(\u1/out9 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__206
       (.I0(\u1/u9/X [5]),
        .I1(\u1/u9/X [4]),
        .I2(\u1/u9/X [3]),
        .I3(\u1/u9/X [2]),
        .I4(\u1/u9/X [6]),
        .I5(\u1/u9/X [1]),
        .O(\u1/out9 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__207
       (.I0(\u1/u10/X [41]),
        .I1(\u1/u10/X [40]),
        .I2(\u1/u10/X [39]),
        .I3(\u1/u10/X [38]),
        .I4(\u1/u10/X [42]),
        .I5(\u1/u10/X [37]),
        .O(\u1/out10 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__208
       (.I0(\u1/u10/X [17]),
        .I1(\u1/u10/X [16]),
        .I2(\u1/u10/X [15]),
        .I3(\u1/u10/X [14]),
        .I4(\u1/u10/X [18]),
        .I5(\u1/u10/X [13]),
        .O(\u1/out10 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__209
       (.I0(\u1/u10/X [35]),
        .I1(\u1/u10/X [34]),
        .I2(\u1/u10/X [33]),
        .I3(\u1/u10/X [32]),
        .I4(\u1/u10/X [36]),
        .I5(\u1/u10/X [31]),
        .O(\u1/out10 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__21
       (.I0(\u0/u2/X [29]),
        .I1(\u0/u2/X [28]),
        .I2(\u0/u2/X [27]),
        .I3(\u0/u2/X [26]),
        .I4(\u0/u2/X [30]),
        .I5(\u0/u2/X [25]),
        .O(\u0/out2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__210
       (.I0(\u1/u10/X [11]),
        .I1(\u1/u10/X [10]),
        .I2(\u1/u10/X [9]),
        .I3(\u1/u10/X [8]),
        .I4(\u1/u10/X [12]),
        .I5(\u1/u10/X [7]),
        .O(\u1/out10 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__211
       (.I0(\u1/u10/X [47]),
        .I1(\u1/u10/X [46]),
        .I2(\u1/u10/X [45]),
        .I3(\u1/u10/X [44]),
        .I4(\u1/u10/X [48]),
        .I5(\u1/u10/X [43]),
        .O(\u1/out10 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__212
       (.I0(\u1/u10/X [23]),
        .I1(\u1/u10/X [22]),
        .I2(\u1/u10/X [21]),
        .I3(\u1/u10/X [20]),
        .I4(\u1/u10/X [24]),
        .I5(\u1/u10/X [19]),
        .O(\u1/out10 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__213
       (.I0(\u1/u10/X [29]),
        .I1(\u1/u10/X [28]),
        .I2(\u1/u10/X [27]),
        .I3(\u1/u10/X [26]),
        .I4(\u1/u10/X [30]),
        .I5(\u1/u10/X [25]),
        .O(\u1/out10 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__214
       (.I0(\u1/u10/X [5]),
        .I1(\u1/u10/X [4]),
        .I2(\u1/u10/X [3]),
        .I3(\u1/u10/X [2]),
        .I4(\u1/u10/X [6]),
        .I5(\u1/u10/X [1]),
        .O(\u1/out10 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__215
       (.I0(\u1/u11/X [41]),
        .I1(\u1/u11/X [40]),
        .I2(\u1/u11/X [39]),
        .I3(\u1/u11/X [38]),
        .I4(\u1/u11/X [42]),
        .I5(\u1/u11/X [37]),
        .O(\u1/out11 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__216
       (.I0(\u1/u11/X [17]),
        .I1(\u1/u11/X [16]),
        .I2(\u1/u11/X [15]),
        .I3(\u1/u11/X [14]),
        .I4(\u1/u11/X [18]),
        .I5(\u1/u11/X [13]),
        .O(\u1/out11 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__217
       (.I0(\u1/u11/X [35]),
        .I1(\u1/u11/X [34]),
        .I2(\u1/u11/X [33]),
        .I3(\u1/u11/X [32]),
        .I4(\u1/u11/X [36]),
        .I5(\u1/u11/X [31]),
        .O(\u1/out11 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__218
       (.I0(\u1/u11/X [11]),
        .I1(\u1/u11/X [10]),
        .I2(\u1/u11/X [9]),
        .I3(\u1/u11/X [8]),
        .I4(\u1/u11/X [12]),
        .I5(\u1/u11/X [7]),
        .O(\u1/out11 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__219
       (.I0(\u1/u11/X [47]),
        .I1(\u1/u11/X [46]),
        .I2(\u1/u11/X [45]),
        .I3(\u1/u11/X [44]),
        .I4(\u1/u11/X [48]),
        .I5(\u1/u11/X [43]),
        .O(\u1/out11 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__22
       (.I0(\u0/u2/X [5]),
        .I1(\u0/u2/X [4]),
        .I2(\u0/u2/X [3]),
        .I3(\u0/u2/X [2]),
        .I4(\u0/u2/X [6]),
        .I5(\u0/u2/X [1]),
        .O(\u0/out2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__220
       (.I0(\u1/u11/X [23]),
        .I1(\u1/u11/X [22]),
        .I2(\u1/u11/X [21]),
        .I3(\u1/u11/X [20]),
        .I4(\u1/u11/X [24]),
        .I5(\u1/u11/X [19]),
        .O(\u1/out11 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__221
       (.I0(\u1/u11/X [29]),
        .I1(\u1/u11/X [28]),
        .I2(\u1/u11/X [27]),
        .I3(\u1/u11/X [26]),
        .I4(\u1/u11/X [30]),
        .I5(\u1/u11/X [25]),
        .O(\u1/out11 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__222
       (.I0(\u1/u11/X [5]),
        .I1(\u1/u11/X [4]),
        .I2(\u1/u11/X [3]),
        .I3(\u1/u11/X [2]),
        .I4(\u1/u11/X [6]),
        .I5(\u1/u11/X [1]),
        .O(\u1/out11 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__223
       (.I0(\u1/u12/X [41]),
        .I1(\u1/u12/X [40]),
        .I2(\u1/u12/X [39]),
        .I3(\u1/u12/X [38]),
        .I4(\u1/u12/X [42]),
        .I5(\u1/u12/X [37]),
        .O(\u1/out12 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__224
       (.I0(\u1/u12/X [17]),
        .I1(\u1/u12/X [16]),
        .I2(\u1/u12/X [15]),
        .I3(\u1/u12/X [14]),
        .I4(\u1/u12/X [18]),
        .I5(\u1/u12/X [13]),
        .O(\u1/out12 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__225
       (.I0(\u1/u12/X [35]),
        .I1(\u1/u12/X [34]),
        .I2(\u1/u12/X [33]),
        .I3(\u1/u12/X [32]),
        .I4(\u1/u12/X [36]),
        .I5(\u1/u12/X [31]),
        .O(\u1/out12 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__226
       (.I0(\u1/u12/X [11]),
        .I1(\u1/u12/X [10]),
        .I2(\u1/u12/X [9]),
        .I3(\u1/u12/X [8]),
        .I4(\u1/u12/X [12]),
        .I5(\u1/u12/X [7]),
        .O(\u1/out12 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__227
       (.I0(\u1/u12/X [47]),
        .I1(\u1/u12/X [46]),
        .I2(\u1/u12/X [45]),
        .I3(\u1/u12/X [44]),
        .I4(\u1/u12/X [48]),
        .I5(\u1/u12/X [43]),
        .O(\u1/out12 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__228
       (.I0(\u1/u12/X [23]),
        .I1(\u1/u12/X [22]),
        .I2(\u1/u12/X [21]),
        .I3(\u1/u12/X [20]),
        .I4(\u1/u12/X [24]),
        .I5(\u1/u12/X [19]),
        .O(\u1/out12 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__229
       (.I0(\u1/u12/X [29]),
        .I1(\u1/u12/X [28]),
        .I2(\u1/u12/X [27]),
        .I3(\u1/u12/X [26]),
        .I4(\u1/u12/X [30]),
        .I5(\u1/u12/X [25]),
        .O(\u1/out12 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__23
       (.I0(\u0/u3/X [41]),
        .I1(\u0/u3/X [40]),
        .I2(\u0/u3/X [39]),
        .I3(\u0/u3/X [38]),
        .I4(\u0/u3/X [42]),
        .I5(\u0/u3/X [37]),
        .O(\u0/out3 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__230
       (.I0(\u1/u12/X [5]),
        .I1(\u1/u12/X [4]),
        .I2(\u1/u12/X [3]),
        .I3(\u1/u12/X [2]),
        .I4(\u1/u12/X [6]),
        .I5(\u1/u12/X [1]),
        .O(\u1/out12 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__231
       (.I0(\u1/u13/X [41]),
        .I1(\u1/u13/X [40]),
        .I2(\u1/u13/X [39]),
        .I3(\u1/u13/X [38]),
        .I4(\u1/u13/X [42]),
        .I5(\u1/u13/X [37]),
        .O(\u1/out13 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__232
       (.I0(\u1/u13/X [17]),
        .I1(\u1/u13/X [16]),
        .I2(\u1/u13/X [15]),
        .I3(\u1/u13/X [14]),
        .I4(\u1/u13/X [18]),
        .I5(\u1/u13/X [13]),
        .O(\u1/out13 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__233
       (.I0(\u1/u13/X [35]),
        .I1(\u1/u13/X [34]),
        .I2(\u1/u13/X [33]),
        .I3(\u1/u13/X [32]),
        .I4(\u1/u13/X [36]),
        .I5(\u1/u13/X [31]),
        .O(\u1/out13 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__234
       (.I0(\u1/u13/X [11]),
        .I1(\u1/u13/X [10]),
        .I2(\u1/u13/X [9]),
        .I3(\u1/u13/X [8]),
        .I4(\u1/u13/X [12]),
        .I5(\u1/u13/X [7]),
        .O(\u1/out13 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__235
       (.I0(\u1/u13/X [47]),
        .I1(\u1/u13/X [46]),
        .I2(\u1/u13/X [45]),
        .I3(\u1/u13/X [44]),
        .I4(\u1/u13/X [48]),
        .I5(\u1/u13/X [43]),
        .O(\u1/out13 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__236
       (.I0(\u1/u13/X [23]),
        .I1(\u1/u13/X [22]),
        .I2(\u1/u13/X [21]),
        .I3(\u1/u13/X [20]),
        .I4(\u1/u13/X [24]),
        .I5(\u1/u13/X [19]),
        .O(\u1/out13 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__237
       (.I0(\u1/u13/X [29]),
        .I1(\u1/u13/X [28]),
        .I2(\u1/u13/X [27]),
        .I3(\u1/u13/X [26]),
        .I4(\u1/u13/X [30]),
        .I5(\u1/u13/X [25]),
        .O(\u1/out13 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__238
       (.I0(\u1/u13/X [5]),
        .I1(\u1/u13/X [4]),
        .I2(\u1/u13/X [3]),
        .I3(\u1/u13/X [2]),
        .I4(\u1/u13/X [6]),
        .I5(\u1/u13/X [1]),
        .O(\u1/out13 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__239
       (.I0(\u1/u14/X [41]),
        .I1(\u1/u14/X [40]),
        .I2(\u1/u14/X [39]),
        .I3(\u1/u14/X [38]),
        .I4(\u1/u14/X [42]),
        .I5(\u1/u14/X [37]),
        .O(\u1/out14 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__24
       (.I0(\u0/u3/X [17]),
        .I1(\u0/u3/X [16]),
        .I2(\u0/u3/X [15]),
        .I3(\u0/u3/X [14]),
        .I4(\u0/u3/X [18]),
        .I5(\u0/u3/X [13]),
        .O(\u0/out3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__240
       (.I0(\u1/u14/X [17]),
        .I1(\u1/u14/X [16]),
        .I2(\u1/u14/X [15]),
        .I3(\u1/u14/X [14]),
        .I4(\u1/u14/X [18]),
        .I5(\u1/u14/X [13]),
        .O(\u1/out14 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__241
       (.I0(\u1/u14/X [35]),
        .I1(\u1/u14/X [34]),
        .I2(\u1/u14/X [33]),
        .I3(\u1/u14/X [32]),
        .I4(\u1/u14/X [36]),
        .I5(\u1/u14/X [31]),
        .O(\u1/out14 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__242
       (.I0(\u1/u14/X [11]),
        .I1(\u1/u14/X [10]),
        .I2(\u1/u14/X [9]),
        .I3(\u1/u14/X [8]),
        .I4(\u1/u14/X [12]),
        .I5(\u1/u14/X [7]),
        .O(\u1/out14 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__243
       (.I0(\u1/u14/X [47]),
        .I1(\u1/u14/X [46]),
        .I2(\u1/u14/X [45]),
        .I3(\u1/u14/X [44]),
        .I4(\u1/u14/X [48]),
        .I5(\u1/u14/X [43]),
        .O(\u1/out14 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__244
       (.I0(\u1/u14/X [23]),
        .I1(\u1/u14/X [22]),
        .I2(\u1/u14/X [21]),
        .I3(\u1/u14/X [20]),
        .I4(\u1/u14/X [24]),
        .I5(\u1/u14/X [19]),
        .O(\u1/out14 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__245
       (.I0(\u1/u14/X [29]),
        .I1(\u1/u14/X [28]),
        .I2(\u1/u14/X [27]),
        .I3(\u1/u14/X [26]),
        .I4(\u1/u14/X [30]),
        .I5(\u1/u14/X [25]),
        .O(\u1/out14 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__246
       (.I0(\u1/u14/X [5]),
        .I1(\u1/u14/X [4]),
        .I2(\u1/u14/X [3]),
        .I3(\u1/u14/X [2]),
        .I4(\u1/u14/X [6]),
        .I5(\u1/u14/X [1]),
        .O(\u1/out14 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__247
       (.I0(\u1/u15/X [41]),
        .I1(\u1/u15/X [40]),
        .I2(\u1/u15/X [39]),
        .I3(\u1/u15/X [38]),
        .I4(\u1/u15/X [42]),
        .I5(\u1/u15/X [37]),
        .O(\u1/out15 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__248
       (.I0(\u1/u15/X [17]),
        .I1(\u1/u15/X [16]),
        .I2(\u1/u15/X [15]),
        .I3(\u1/u15/X [14]),
        .I4(\u1/u15/X [18]),
        .I5(\u1/u15/X [13]),
        .O(\u1/out15 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__249
       (.I0(\u1/u15/X [35]),
        .I1(\u1/u15/X [34]),
        .I2(\u1/u15/X [33]),
        .I3(\u1/u15/X [32]),
        .I4(\u1/u15/X [36]),
        .I5(\u1/u15/X [31]),
        .O(\u1/out15 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__25
       (.I0(\u0/u3/X [35]),
        .I1(\u0/u3/X [34]),
        .I2(\u0/u3/X [33]),
        .I3(\u0/u3/X [32]),
        .I4(\u0/u3/X [36]),
        .I5(\u0/u3/X [31]),
        .O(\u0/out3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__250
       (.I0(\u1/u15/X [11]),
        .I1(\u1/u15/X [10]),
        .I2(\u1/u15/X [9]),
        .I3(\u1/u15/X [8]),
        .I4(\u1/u15/X [12]),
        .I5(\u1/u15/X [7]),
        .O(\u1/out15 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__251
       (.I0(\u1/u15/X [47]),
        .I1(\u1/u15/X [46]),
        .I2(\u1/u15/X [45]),
        .I3(\u1/u15/X [44]),
        .I4(\u1/u15/X [48]),
        .I5(\u1/u15/X [43]),
        .O(\u1/out15 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__252
       (.I0(\u1/u15/X [23]),
        .I1(\u1/u15/X [22]),
        .I2(\u1/u15/X [21]),
        .I3(\u1/u15/X [20]),
        .I4(\u1/u15/X [24]),
        .I5(\u1/u15/X [19]),
        .O(\u1/out15 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__253
       (.I0(\u1/u15/X [29]),
        .I1(\u1/u15/X [28]),
        .I2(\u1/u15/X [27]),
        .I3(\u1/u15/X [26]),
        .I4(\u1/u15/X [30]),
        .I5(\u1/u15/X [25]),
        .O(\u1/out15 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__254
       (.I0(\u1/u15/X [5]),
        .I1(\u1/u15/X [4]),
        .I2(\u1/u15/X [3]),
        .I3(\u1/u15/X [2]),
        .I4(\u1/u15/X [6]),
        .I5(\u1/u15/X [1]),
        .O(\u1/out15 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__255
       (.I0(\u2/u0/X [41]),
        .I1(\u2/u0/X [40]),
        .I2(\u2/u0/X [39]),
        .I3(\u2/u0/X [38]),
        .I4(\u2/u0/X [42]),
        .I5(\u2/u0/X [37]),
        .O(\u2/out0 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__256
       (.I0(\u2/u0/X [17]),
        .I1(\u2/u0/X [16]),
        .I2(\u2/u0/X [15]),
        .I3(\u2/u0/X [14]),
        .I4(\u2/u0/X [18]),
        .I5(\u2/u0/X [13]),
        .O(\u2/out0 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__257
       (.I0(\u2/u0/X [35]),
        .I1(\u2/u0/X [34]),
        .I2(\u2/u0/X [33]),
        .I3(\u2/u0/X [32]),
        .I4(\u2/u0/X [36]),
        .I5(\u2/u0/X [31]),
        .O(\u2/out0 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__258
       (.I0(\u2/u0/X [11]),
        .I1(\u2/u0/X [10]),
        .I2(\u2/u0/X [9]),
        .I3(\u2/u0/X [8]),
        .I4(\u2/u0/X [12]),
        .I5(\u2/u0/X [7]),
        .O(\u2/out0 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__259
       (.I0(\u2/u0/X [47]),
        .I1(\u2/u0/X [46]),
        .I2(\u2/u0/X [45]),
        .I3(\u2/u0/X [44]),
        .I4(\u2/u0/X [48]),
        .I5(\u2/u0/X [43]),
        .O(\u2/out0 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__26
       (.I0(\u0/u3/X [11]),
        .I1(\u0/u3/X [10]),
        .I2(\u0/u3/X [9]),
        .I3(\u0/u3/X [8]),
        .I4(\u0/u3/X [12]),
        .I5(\u0/u3/X [7]),
        .O(\u0/out3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__260
       (.I0(\u2/u0/X [23]),
        .I1(\u2/u0/X [22]),
        .I2(\u2/u0/X [21]),
        .I3(\u2/u0/X [20]),
        .I4(\u2/u0/X [24]),
        .I5(\u2/u0/X [19]),
        .O(\u2/out0 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__261
       (.I0(\u2/u0/X [29]),
        .I1(\u2/u0/X [28]),
        .I2(\u2/u0/X [27]),
        .I3(\u2/u0/X [26]),
        .I4(\u2/u0/X [30]),
        .I5(\u2/u0/X [25]),
        .O(\u2/out0 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__262
       (.I0(\u2/u0/X [5]),
        .I1(\u2/u0/X [4]),
        .I2(\u2/u0/X [3]),
        .I3(\u2/u0/X [2]),
        .I4(\u2/u0/X [6]),
        .I5(\u2/u0/X [1]),
        .O(\u2/out0 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__263
       (.I0(\u2/u1/X [41]),
        .I1(\u2/u1/X [40]),
        .I2(\u2/u1/X [39]),
        .I3(\u2/u1/X [38]),
        .I4(\u2/u1/X [42]),
        .I5(\u2/u1/X [37]),
        .O(\u2/out1 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__264
       (.I0(\u2/u1/X [17]),
        .I1(\u2/u1/X [16]),
        .I2(\u2/u1/X [15]),
        .I3(\u2/u1/X [14]),
        .I4(\u2/u1/X [18]),
        .I5(\u2/u1/X [13]),
        .O(\u2/out1 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__265
       (.I0(\u2/u1/X [35]),
        .I1(\u2/u1/X [34]),
        .I2(\u2/u1/X [33]),
        .I3(\u2/u1/X [32]),
        .I4(\u2/u1/X [36]),
        .I5(\u2/u1/X [31]),
        .O(\u2/out1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__266
       (.I0(\u2/u1/X [11]),
        .I1(\u2/u1/X [10]),
        .I2(\u2/u1/X [9]),
        .I3(\u2/u1/X [8]),
        .I4(\u2/u1/X [12]),
        .I5(\u2/u1/X [7]),
        .O(\u2/out1 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__267
       (.I0(\u2/u1/X [47]),
        .I1(\u2/u1/X [46]),
        .I2(\u2/u1/X [45]),
        .I3(\u2/u1/X [44]),
        .I4(\u2/u1/X [48]),
        .I5(\u2/u1/X [43]),
        .O(\u2/out1 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__268
       (.I0(\u2/u1/X [23]),
        .I1(\u2/u1/X [22]),
        .I2(\u2/u1/X [21]),
        .I3(\u2/u1/X [20]),
        .I4(\u2/u1/X [24]),
        .I5(\u2/u1/X [19]),
        .O(\u2/out1 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__269
       (.I0(\u2/u1/X [29]),
        .I1(\u2/u1/X [28]),
        .I2(\u2/u1/X [27]),
        .I3(\u2/u1/X [26]),
        .I4(\u2/u1/X [30]),
        .I5(\u2/u1/X [25]),
        .O(\u2/out1 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__27
       (.I0(\u0/u3/X [47]),
        .I1(\u0/u3/X [46]),
        .I2(\u0/u3/X [45]),
        .I3(\u0/u3/X [44]),
        .I4(\u0/u3/X [48]),
        .I5(\u0/u3/X [43]),
        .O(\u0/out3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__270
       (.I0(\u2/u1/X [5]),
        .I1(\u2/u1/X [4]),
        .I2(\u2/u1/X [3]),
        .I3(\u2/u1/X [2]),
        .I4(\u2/u1/X [6]),
        .I5(\u2/u1/X [1]),
        .O(\u2/out1 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__271
       (.I0(\u2/u2/X [41]),
        .I1(\u2/u2/X [40]),
        .I2(\u2/u2/X [39]),
        .I3(\u2/u2/X [38]),
        .I4(\u2/u2/X [42]),
        .I5(\u2/u2/X [37]),
        .O(\u2/out2 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__272
       (.I0(\u2/u2/X [17]),
        .I1(\u2/u2/X [16]),
        .I2(\u2/u2/X [15]),
        .I3(\u2/u2/X [14]),
        .I4(\u2/u2/X [18]),
        .I5(\u2/u2/X [13]),
        .O(\u2/out2 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__273
       (.I0(\u2/u2/X [35]),
        .I1(\u2/u2/X [34]),
        .I2(\u2/u2/X [33]),
        .I3(\u2/u2/X [32]),
        .I4(\u2/u2/X [36]),
        .I5(\u2/u2/X [31]),
        .O(\u2/out2 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__274
       (.I0(\u2/u2/X [11]),
        .I1(\u2/u2/X [10]),
        .I2(\u2/u2/X [9]),
        .I3(\u2/u2/X [8]),
        .I4(\u2/u2/X [12]),
        .I5(\u2/u2/X [7]),
        .O(\u2/out2 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__275
       (.I0(\u2/u2/X [47]),
        .I1(\u2/u2/X [46]),
        .I2(\u2/u2/X [45]),
        .I3(\u2/u2/X [44]),
        .I4(\u2/u2/X [48]),
        .I5(\u2/u2/X [43]),
        .O(\u2/out2 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__276
       (.I0(\u2/u2/X [23]),
        .I1(\u2/u2/X [22]),
        .I2(\u2/u2/X [21]),
        .I3(\u2/u2/X [20]),
        .I4(\u2/u2/X [24]),
        .I5(\u2/u2/X [19]),
        .O(\u2/out2 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__277
       (.I0(\u2/u2/X [29]),
        .I1(\u2/u2/X [28]),
        .I2(\u2/u2/X [27]),
        .I3(\u2/u2/X [26]),
        .I4(\u2/u2/X [30]),
        .I5(\u2/u2/X [25]),
        .O(\u2/out2 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__278
       (.I0(\u2/u2/X [5]),
        .I1(\u2/u2/X [4]),
        .I2(\u2/u2/X [3]),
        .I3(\u2/u2/X [2]),
        .I4(\u2/u2/X [6]),
        .I5(\u2/u2/X [1]),
        .O(\u2/out2 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__279
       (.I0(\u2/u3/X [41]),
        .I1(\u2/u3/X [40]),
        .I2(\u2/u3/X [39]),
        .I3(\u2/u3/X [38]),
        .I4(\u2/u3/X [42]),
        .I5(\u2/u3/X [37]),
        .O(\u2/out3 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__28
       (.I0(\u0/u3/X [23]),
        .I1(\u0/u3/X [22]),
        .I2(\u0/u3/X [21]),
        .I3(\u0/u3/X [20]),
        .I4(\u0/u3/X [24]),
        .I5(\u0/u3/X [19]),
        .O(\u0/out3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__280
       (.I0(\u2/u3/X [17]),
        .I1(\u2/u3/X [16]),
        .I2(\u2/u3/X [15]),
        .I3(\u2/u3/X [14]),
        .I4(\u2/u3/X [18]),
        .I5(\u2/u3/X [13]),
        .O(\u2/out3 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__281
       (.I0(\u2/u3/X [35]),
        .I1(\u2/u3/X [34]),
        .I2(\u2/u3/X [33]),
        .I3(\u2/u3/X [32]),
        .I4(\u2/u3/X [36]),
        .I5(\u2/u3/X [31]),
        .O(\u2/out3 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__282
       (.I0(\u2/u3/X [11]),
        .I1(\u2/u3/X [10]),
        .I2(\u2/u3/X [9]),
        .I3(\u2/u3/X [8]),
        .I4(\u2/u3/X [12]),
        .I5(\u2/u3/X [7]),
        .O(\u2/out3 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__283
       (.I0(\u2/u3/X [47]),
        .I1(\u2/u3/X [46]),
        .I2(\u2/u3/X [45]),
        .I3(\u2/u3/X [44]),
        .I4(\u2/u3/X [48]),
        .I5(\u2/u3/X [43]),
        .O(\u2/out3 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__284
       (.I0(\u2/u3/X [23]),
        .I1(\u2/u3/X [22]),
        .I2(\u2/u3/X [21]),
        .I3(\u2/u3/X [20]),
        .I4(\u2/u3/X [24]),
        .I5(\u2/u3/X [19]),
        .O(\u2/out3 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__285
       (.I0(\u2/u3/X [29]),
        .I1(\u2/u3/X [28]),
        .I2(\u2/u3/X [27]),
        .I3(\u2/u3/X [26]),
        .I4(\u2/u3/X [30]),
        .I5(\u2/u3/X [25]),
        .O(\u2/out3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__286
       (.I0(\u2/u3/X [5]),
        .I1(\u2/u3/X [4]),
        .I2(\u2/u3/X [3]),
        .I3(\u2/u3/X [2]),
        .I4(\u2/u3/X [6]),
        .I5(\u2/u3/X [1]),
        .O(\u2/out3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__287
       (.I0(\u2/u4/X [41]),
        .I1(\u2/u4/X [40]),
        .I2(\u2/u4/X [39]),
        .I3(\u2/u4/X [38]),
        .I4(\u2/u4/X [42]),
        .I5(\u2/u4/X [37]),
        .O(\u2/out4 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__288
       (.I0(\u2/u4/X [17]),
        .I1(\u2/u4/X [16]),
        .I2(\u2/u4/X [15]),
        .I3(\u2/u4/X [14]),
        .I4(\u2/u4/X [18]),
        .I5(\u2/u4/X [13]),
        .O(\u2/out4 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__289
       (.I0(\u2/u4/X [35]),
        .I1(\u2/u4/X [34]),
        .I2(\u2/u4/X [33]),
        .I3(\u2/u4/X [32]),
        .I4(\u2/u4/X [36]),
        .I5(\u2/u4/X [31]),
        .O(\u2/out4 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__29
       (.I0(\u0/u3/X [29]),
        .I1(\u0/u3/X [28]),
        .I2(\u0/u3/X [27]),
        .I3(\u0/u3/X [26]),
        .I4(\u0/u3/X [30]),
        .I5(\u0/u3/X [25]),
        .O(\u0/out3 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__290
       (.I0(\u2/u4/X [11]),
        .I1(\u2/u4/X [10]),
        .I2(\u2/u4/X [9]),
        .I3(\u2/u4/X [8]),
        .I4(\u2/u4/X [12]),
        .I5(\u2/u4/X [7]),
        .O(\u2/out4 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__291
       (.I0(\u2/u4/X [47]),
        .I1(\u2/u4/X [46]),
        .I2(\u2/u4/X [45]),
        .I3(\u2/u4/X [44]),
        .I4(\u2/u4/X [48]),
        .I5(\u2/u4/X [43]),
        .O(\u2/out4 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__292
       (.I0(\u2/u4/X [23]),
        .I1(\u2/u4/X [22]),
        .I2(\u2/u4/X [21]),
        .I3(\u2/u4/X [20]),
        .I4(\u2/u4/X [24]),
        .I5(\u2/u4/X [19]),
        .O(\u2/out4 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__293
       (.I0(\u2/u4/X [29]),
        .I1(\u2/u4/X [28]),
        .I2(\u2/u4/X [27]),
        .I3(\u2/u4/X [26]),
        .I4(\u2/u4/X [30]),
        .I5(\u2/u4/X [25]),
        .O(\u2/out4 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__294
       (.I0(\u2/u4/X [5]),
        .I1(\u2/u4/X [4]),
        .I2(\u2/u4/X [3]),
        .I3(\u2/u4/X [2]),
        .I4(\u2/u4/X [6]),
        .I5(\u2/u4/X [1]),
        .O(\u2/out4 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__295
       (.I0(\u2/u5/X [41]),
        .I1(\u2/u5/X [40]),
        .I2(\u2/u5/X [39]),
        .I3(\u2/u5/X [38]),
        .I4(\u2/u5/X [42]),
        .I5(\u2/u5/X [37]),
        .O(\u2/out5 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__296
       (.I0(\u2/u5/X [17]),
        .I1(\u2/u5/X [16]),
        .I2(\u2/u5/X [15]),
        .I3(\u2/u5/X [14]),
        .I4(\u2/u5/X [18]),
        .I5(\u2/u5/X [13]),
        .O(\u2/out5 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__297
       (.I0(\u2/u5/X [35]),
        .I1(\u2/u5/X [34]),
        .I2(\u2/u5/X [33]),
        .I3(\u2/u5/X [32]),
        .I4(\u2/u5/X [36]),
        .I5(\u2/u5/X [31]),
        .O(\u2/out5 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__298
       (.I0(\u2/u5/X [11]),
        .I1(\u2/u5/X [10]),
        .I2(\u2/u5/X [9]),
        .I3(\u2/u5/X [8]),
        .I4(\u2/u5/X [12]),
        .I5(\u2/u5/X [7]),
        .O(\u2/out5 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__299
       (.I0(\u2/u5/X [47]),
        .I1(\u2/u5/X [46]),
        .I2(\u2/u5/X [45]),
        .I3(\u2/u5/X [44]),
        .I4(\u2/u5/X [48]),
        .I5(\u2/u5/X [43]),
        .O(\u2/out5 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__3
       (.I0(\u0/u0/X [47]),
        .I1(\u0/u0/X [46]),
        .I2(\u0/u0/X [45]),
        .I3(\u0/u0/X [44]),
        .I4(\u0/u0/X [48]),
        .I5(\u0/u0/X [43]),
        .O(\u0/out0 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__30
       (.I0(\u0/u3/X [5]),
        .I1(\u0/u3/X [4]),
        .I2(\u0/u3/X [3]),
        .I3(\u0/u3/X [2]),
        .I4(\u0/u3/X [6]),
        .I5(\u0/u3/X [1]),
        .O(\u0/out3 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__300
       (.I0(\u2/u5/X [23]),
        .I1(\u2/u5/X [22]),
        .I2(\u2/u5/X [21]),
        .I3(\u2/u5/X [20]),
        .I4(\u2/u5/X [24]),
        .I5(\u2/u5/X [19]),
        .O(\u2/out5 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__301
       (.I0(\u2/u5/X [29]),
        .I1(\u2/u5/X [28]),
        .I2(\u2/u5/X [27]),
        .I3(\u2/u5/X [26]),
        .I4(\u2/u5/X [30]),
        .I5(\u2/u5/X [25]),
        .O(\u2/out5 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__302
       (.I0(\u2/u5/X [5]),
        .I1(\u2/u5/X [4]),
        .I2(\u2/u5/X [3]),
        .I3(\u2/u5/X [2]),
        .I4(\u2/u5/X [6]),
        .I5(\u2/u5/X [1]),
        .O(\u2/out5 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__303
       (.I0(\u2/u6/X [41]),
        .I1(\u2/u6/X [40]),
        .I2(\u2/u6/X [39]),
        .I3(\u2/u6/X [38]),
        .I4(\u2/u6/X [42]),
        .I5(\u2/u6/X [37]),
        .O(\u2/out6 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__304
       (.I0(\u2/u6/X [17]),
        .I1(\u2/u6/X [16]),
        .I2(\u2/u6/X [15]),
        .I3(\u2/u6/X [14]),
        .I4(\u2/u6/X [18]),
        .I5(\u2/u6/X [13]),
        .O(\u2/out6 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__305
       (.I0(\u2/u6/X [35]),
        .I1(\u2/u6/X [34]),
        .I2(\u2/u6/X [33]),
        .I3(\u2/u6/X [32]),
        .I4(\u2/u6/X [36]),
        .I5(\u2/u6/X [31]),
        .O(\u2/out6 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__306
       (.I0(\u2/u6/X [11]),
        .I1(\u2/u6/X [10]),
        .I2(\u2/u6/X [9]),
        .I3(\u2/u6/X [8]),
        .I4(\u2/u6/X [12]),
        .I5(\u2/u6/X [7]),
        .O(\u2/out6 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__307
       (.I0(\u2/u6/X [47]),
        .I1(\u2/u6/X [46]),
        .I2(\u2/u6/X [45]),
        .I3(\u2/u6/X [44]),
        .I4(\u2/u6/X [48]),
        .I5(\u2/u6/X [43]),
        .O(\u2/out6 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__308
       (.I0(\u2/u6/X [23]),
        .I1(\u2/u6/X [22]),
        .I2(\u2/u6/X [21]),
        .I3(\u2/u6/X [20]),
        .I4(\u2/u6/X [24]),
        .I5(\u2/u6/X [19]),
        .O(\u2/out6 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__309
       (.I0(\u2/u6/X [29]),
        .I1(\u2/u6/X [28]),
        .I2(\u2/u6/X [27]),
        .I3(\u2/u6/X [26]),
        .I4(\u2/u6/X [30]),
        .I5(\u2/u6/X [25]),
        .O(\u2/out6 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__31
       (.I0(\u0/u4/X [41]),
        .I1(\u0/u4/X [40]),
        .I2(\u0/u4/X [39]),
        .I3(\u0/u4/X [38]),
        .I4(\u0/u4/X [42]),
        .I5(\u0/u4/X [37]),
        .O(\u0/out4 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__310
       (.I0(\u2/u6/X [5]),
        .I1(\u2/u6/X [4]),
        .I2(\u2/u6/X [3]),
        .I3(\u2/u6/X [2]),
        .I4(\u2/u6/X [6]),
        .I5(\u2/u6/X [1]),
        .O(\u2/out6 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__311
       (.I0(\u2/u7/X [41]),
        .I1(\u2/u7/X [40]),
        .I2(\u2/u7/X [39]),
        .I3(\u2/u7/X [38]),
        .I4(\u2/u7/X [42]),
        .I5(\u2/u7/X [37]),
        .O(\u2/out7 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__312
       (.I0(\u2/u7/X [17]),
        .I1(\u2/u7/X [16]),
        .I2(\u2/u7/X [15]),
        .I3(\u2/u7/X [14]),
        .I4(\u2/u7/X [18]),
        .I5(\u2/u7/X [13]),
        .O(\u2/out7 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__313
       (.I0(\u2/u7/X [35]),
        .I1(\u2/u7/X [34]),
        .I2(\u2/u7/X [33]),
        .I3(\u2/u7/X [32]),
        .I4(\u2/u7/X [36]),
        .I5(\u2/u7/X [31]),
        .O(\u2/out7 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__314
       (.I0(\u2/u7/X [11]),
        .I1(\u2/u7/X [10]),
        .I2(\u2/u7/X [9]),
        .I3(\u2/u7/X [8]),
        .I4(\u2/u7/X [12]),
        .I5(\u2/u7/X [7]),
        .O(\u2/out7 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__315
       (.I0(\u2/u7/X [47]),
        .I1(\u2/u7/X [46]),
        .I2(\u2/u7/X [45]),
        .I3(\u2/u7/X [44]),
        .I4(\u2/u7/X [48]),
        .I5(\u2/u7/X [43]),
        .O(\u2/out7 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__316
       (.I0(\u2/u7/X [23]),
        .I1(\u2/u7/X [22]),
        .I2(\u2/u7/X [21]),
        .I3(\u2/u7/X [20]),
        .I4(\u2/u7/X [24]),
        .I5(\u2/u7/X [19]),
        .O(\u2/out7 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__317
       (.I0(\u2/u7/X [29]),
        .I1(\u2/u7/X [28]),
        .I2(\u2/u7/X [27]),
        .I3(\u2/u7/X [26]),
        .I4(\u2/u7/X [30]),
        .I5(\u2/u7/X [25]),
        .O(\u2/out7 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__318
       (.I0(\u2/u7/X [5]),
        .I1(\u2/u7/X [4]),
        .I2(\u2/u7/X [3]),
        .I3(\u2/u7/X [2]),
        .I4(\u2/u7/X [6]),
        .I5(\u2/u7/X [1]),
        .O(\u2/out7 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__319
       (.I0(\u2/u8/X [41]),
        .I1(\u2/u8/X [40]),
        .I2(\u2/u8/X [39]),
        .I3(\u2/u8/X [38]),
        .I4(\u2/u8/X [42]),
        .I5(\u2/u8/X [37]),
        .O(\u2/out8 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__32
       (.I0(\u0/u4/X [17]),
        .I1(\u0/u4/X [16]),
        .I2(\u0/u4/X [15]),
        .I3(\u0/u4/X [14]),
        .I4(\u0/u4/X [18]),
        .I5(\u0/u4/X [13]),
        .O(\u0/out4 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__320
       (.I0(\u2/u8/X [17]),
        .I1(\u2/u8/X [16]),
        .I2(\u2/u8/X [15]),
        .I3(\u2/u8/X [14]),
        .I4(\u2/u8/X [18]),
        .I5(\u2/u8/X [13]),
        .O(\u2/out8 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__321
       (.I0(\u2/u8/X [35]),
        .I1(\u2/u8/X [34]),
        .I2(\u2/u8/X [33]),
        .I3(\u2/u8/X [32]),
        .I4(\u2/u8/X [36]),
        .I5(\u2/u8/X [31]),
        .O(\u2/out8 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__322
       (.I0(\u2/u8/X [11]),
        .I1(\u2/u8/X [10]),
        .I2(\u2/u8/X [9]),
        .I3(\u2/u8/X [8]),
        .I4(\u2/u8/X [12]),
        .I5(\u2/u8/X [7]),
        .O(\u2/out8 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__323
       (.I0(\u2/u8/X [47]),
        .I1(\u2/u8/X [46]),
        .I2(\u2/u8/X [45]),
        .I3(\u2/u8/X [44]),
        .I4(\u2/u8/X [48]),
        .I5(\u2/u8/X [43]),
        .O(\u2/out8 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__324
       (.I0(\u2/u8/X [23]),
        .I1(\u2/u8/X [22]),
        .I2(\u2/u8/X [21]),
        .I3(\u2/u8/X [20]),
        .I4(\u2/u8/X [24]),
        .I5(\u2/u8/X [19]),
        .O(\u2/out8 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__325
       (.I0(\u2/u8/X [29]),
        .I1(\u2/u8/X [28]),
        .I2(\u2/u8/X [27]),
        .I3(\u2/u8/X [26]),
        .I4(\u2/u8/X [30]),
        .I5(\u2/u8/X [25]),
        .O(\u2/out8 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__326
       (.I0(\u2/u8/X [5]),
        .I1(\u2/u8/X [4]),
        .I2(\u2/u8/X [3]),
        .I3(\u2/u8/X [2]),
        .I4(\u2/u8/X [6]),
        .I5(\u2/u8/X [1]),
        .O(\u2/out8 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__327
       (.I0(\u2/u9/X [41]),
        .I1(\u2/u9/X [40]),
        .I2(\u2/u9/X [39]),
        .I3(\u2/u9/X [38]),
        .I4(\u2/u9/X [42]),
        .I5(\u2/u9/X [37]),
        .O(\u2/out9 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__328
       (.I0(\u2/u9/X [17]),
        .I1(\u2/u9/X [16]),
        .I2(\u2/u9/X [15]),
        .I3(\u2/u9/X [14]),
        .I4(\u2/u9/X [18]),
        .I5(\u2/u9/X [13]),
        .O(\u2/out9 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__329
       (.I0(\u2/u9/X [35]),
        .I1(\u2/u9/X [34]),
        .I2(\u2/u9/X [33]),
        .I3(\u2/u9/X [32]),
        .I4(\u2/u9/X [36]),
        .I5(\u2/u9/X [31]),
        .O(\u2/out9 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__33
       (.I0(\u0/u4/X [35]),
        .I1(\u0/u4/X [34]),
        .I2(\u0/u4/X [33]),
        .I3(\u0/u4/X [32]),
        .I4(\u0/u4/X [36]),
        .I5(\u0/u4/X [31]),
        .O(\u0/out4 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__330
       (.I0(\u2/u9/X [11]),
        .I1(\u2/u9/X [10]),
        .I2(\u2/u9/X [9]),
        .I3(\u2/u9/X [8]),
        .I4(\u2/u9/X [12]),
        .I5(\u2/u9/X [7]),
        .O(\u2/out9 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__331
       (.I0(\u2/u9/X [47]),
        .I1(\u2/u9/X [46]),
        .I2(\u2/u9/X [45]),
        .I3(\u2/u9/X [44]),
        .I4(\u2/u9/X [48]),
        .I5(\u2/u9/X [43]),
        .O(\u2/out9 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__332
       (.I0(\u2/u9/X [23]),
        .I1(\u2/u9/X [22]),
        .I2(\u2/u9/X [21]),
        .I3(\u2/u9/X [20]),
        .I4(\u2/u9/X [24]),
        .I5(\u2/u9/X [19]),
        .O(\u2/out9 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__333
       (.I0(\u2/u9/X [29]),
        .I1(\u2/u9/X [28]),
        .I2(\u2/u9/X [27]),
        .I3(\u2/u9/X [26]),
        .I4(\u2/u9/X [30]),
        .I5(\u2/u9/X [25]),
        .O(\u2/out9 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__334
       (.I0(\u2/u9/X [5]),
        .I1(\u2/u9/X [4]),
        .I2(\u2/u9/X [3]),
        .I3(\u2/u9/X [2]),
        .I4(\u2/u9/X [6]),
        .I5(\u2/u9/X [1]),
        .O(\u2/out9 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__335
       (.I0(\u2/u10/X [41]),
        .I1(\u2/u10/X [40]),
        .I2(\u2/u10/X [39]),
        .I3(\u2/u10/X [38]),
        .I4(\u2/u10/X [42]),
        .I5(\u2/u10/X [37]),
        .O(\u2/out10 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__336
       (.I0(\u2/u10/X [17]),
        .I1(\u2/u10/X [16]),
        .I2(\u2/u10/X [15]),
        .I3(\u2/u10/X [14]),
        .I4(\u2/u10/X [18]),
        .I5(\u2/u10/X [13]),
        .O(\u2/out10 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__337
       (.I0(\u2/u10/X [35]),
        .I1(\u2/u10/X [34]),
        .I2(\u2/u10/X [33]),
        .I3(\u2/u10/X [32]),
        .I4(\u2/u10/X [36]),
        .I5(\u2/u10/X [31]),
        .O(\u2/out10 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__338
       (.I0(\u2/u10/X [11]),
        .I1(\u2/u10/X [10]),
        .I2(\u2/u10/X [9]),
        .I3(\u2/u10/X [8]),
        .I4(\u2/u10/X [12]),
        .I5(\u2/u10/X [7]),
        .O(\u2/out10 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__339
       (.I0(\u2/u10/X [47]),
        .I1(\u2/u10/X [46]),
        .I2(\u2/u10/X [45]),
        .I3(\u2/u10/X [44]),
        .I4(\u2/u10/X [48]),
        .I5(\u2/u10/X [43]),
        .O(\u2/out10 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__34
       (.I0(\u0/u4/X [11]),
        .I1(\u0/u4/X [10]),
        .I2(\u0/u4/X [9]),
        .I3(\u0/u4/X [8]),
        .I4(\u0/u4/X [12]),
        .I5(\u0/u4/X [7]),
        .O(\u0/out4 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__340
       (.I0(\u2/u10/X [23]),
        .I1(\u2/u10/X [22]),
        .I2(\u2/u10/X [21]),
        .I3(\u2/u10/X [20]),
        .I4(\u2/u10/X [24]),
        .I5(\u2/u10/X [19]),
        .O(\u2/out10 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__341
       (.I0(\u2/u10/X [29]),
        .I1(\u2/u10/X [28]),
        .I2(\u2/u10/X [27]),
        .I3(\u2/u10/X [26]),
        .I4(\u2/u10/X [30]),
        .I5(\u2/u10/X [25]),
        .O(\u2/out10 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__342
       (.I0(\u2/u10/X [5]),
        .I1(\u2/u10/X [4]),
        .I2(\u2/u10/X [3]),
        .I3(\u2/u10/X [2]),
        .I4(\u2/u10/X [6]),
        .I5(\u2/u10/X [1]),
        .O(\u2/out10 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__343
       (.I0(\u2/u11/X [41]),
        .I1(\u2/u11/X [40]),
        .I2(\u2/u11/X [39]),
        .I3(\u2/u11/X [38]),
        .I4(\u2/u11/X [42]),
        .I5(\u2/u11/X [37]),
        .O(\u2/out11 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__344
       (.I0(\u2/u11/X [17]),
        .I1(\u2/u11/X [16]),
        .I2(\u2/u11/X [15]),
        .I3(\u2/u11/X [14]),
        .I4(\u2/u11/X [18]),
        .I5(\u2/u11/X [13]),
        .O(\u2/out11 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__345
       (.I0(\u2/u11/X [35]),
        .I1(\u2/u11/X [34]),
        .I2(\u2/u11/X [33]),
        .I3(\u2/u11/X [32]),
        .I4(\u2/u11/X [36]),
        .I5(\u2/u11/X [31]),
        .O(\u2/out11 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__346
       (.I0(\u2/u11/X [11]),
        .I1(\u2/u11/X [10]),
        .I2(\u2/u11/X [9]),
        .I3(\u2/u11/X [8]),
        .I4(\u2/u11/X [12]),
        .I5(\u2/u11/X [7]),
        .O(\u2/out11 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__347
       (.I0(\u2/u11/X [47]),
        .I1(\u2/u11/X [46]),
        .I2(\u2/u11/X [45]),
        .I3(\u2/u11/X [44]),
        .I4(\u2/u11/X [48]),
        .I5(\u2/u11/X [43]),
        .O(\u2/out11 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__348
       (.I0(\u2/u11/X [23]),
        .I1(\u2/u11/X [22]),
        .I2(\u2/u11/X [21]),
        .I3(\u2/u11/X [20]),
        .I4(\u2/u11/X [24]),
        .I5(\u2/u11/X [19]),
        .O(\u2/out11 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__349
       (.I0(\u2/u11/X [29]),
        .I1(\u2/u11/X [28]),
        .I2(\u2/u11/X [27]),
        .I3(\u2/u11/X [26]),
        .I4(\u2/u11/X [30]),
        .I5(\u2/u11/X [25]),
        .O(\u2/out11 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__35
       (.I0(\u0/u4/X [47]),
        .I1(\u0/u4/X [46]),
        .I2(\u0/u4/X [45]),
        .I3(\u0/u4/X [44]),
        .I4(\u0/u4/X [48]),
        .I5(\u0/u4/X [43]),
        .O(\u0/out4 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__350
       (.I0(\u2/u11/X [5]),
        .I1(\u2/u11/X [4]),
        .I2(\u2/u11/X [3]),
        .I3(\u2/u11/X [2]),
        .I4(\u2/u11/X [6]),
        .I5(\u2/u11/X [1]),
        .O(\u2/out11 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__351
       (.I0(\u2/u12/X [41]),
        .I1(\u2/u12/X [40]),
        .I2(\u2/u12/X [39]),
        .I3(\u2/u12/X [38]),
        .I4(\u2/u12/X [42]),
        .I5(\u2/u12/X [37]),
        .O(\u2/out12 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__352
       (.I0(\u2/u12/X [17]),
        .I1(\u2/u12/X [16]),
        .I2(\u2/u12/X [15]),
        .I3(\u2/u12/X [14]),
        .I4(\u2/u12/X [18]),
        .I5(\u2/u12/X [13]),
        .O(\u2/out12 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__353
       (.I0(\u2/u12/X [35]),
        .I1(\u2/u12/X [34]),
        .I2(\u2/u12/X [33]),
        .I3(\u2/u12/X [32]),
        .I4(\u2/u12/X [36]),
        .I5(\u2/u12/X [31]),
        .O(\u2/out12 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__354
       (.I0(\u2/u12/X [11]),
        .I1(\u2/u12/X [10]),
        .I2(\u2/u12/X [9]),
        .I3(\u2/u12/X [8]),
        .I4(\u2/u12/X [12]),
        .I5(\u2/u12/X [7]),
        .O(\u2/out12 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__355
       (.I0(\u2/u12/X [47]),
        .I1(\u2/u12/X [46]),
        .I2(\u2/u12/X [45]),
        .I3(\u2/u12/X [44]),
        .I4(\u2/u12/X [48]),
        .I5(\u2/u12/X [43]),
        .O(\u2/out12 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__356
       (.I0(\u2/u12/X [23]),
        .I1(\u2/u12/X [22]),
        .I2(\u2/u12/X [21]),
        .I3(\u2/u12/X [20]),
        .I4(\u2/u12/X [24]),
        .I5(\u2/u12/X [19]),
        .O(\u2/out12 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__357
       (.I0(\u2/u12/X [29]),
        .I1(\u2/u12/X [28]),
        .I2(\u2/u12/X [27]),
        .I3(\u2/u12/X [26]),
        .I4(\u2/u12/X [30]),
        .I5(\u2/u12/X [25]),
        .O(\u2/out12 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__358
       (.I0(\u2/u12/X [5]),
        .I1(\u2/u12/X [4]),
        .I2(\u2/u12/X [3]),
        .I3(\u2/u12/X [2]),
        .I4(\u2/u12/X [6]),
        .I5(\u2/u12/X [1]),
        .O(\u2/out12 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__359
       (.I0(\u2/u13/X [41]),
        .I1(\u2/u13/X [40]),
        .I2(\u2/u13/X [39]),
        .I3(\u2/u13/X [38]),
        .I4(\u2/u13/X [42]),
        .I5(\u2/u13/X [37]),
        .O(\u2/out13 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__36
       (.I0(\u0/u4/X [23]),
        .I1(\u0/u4/X [22]),
        .I2(\u0/u4/X [21]),
        .I3(\u0/u4/X [20]),
        .I4(\u0/u4/X [24]),
        .I5(\u0/u4/X [19]),
        .O(\u0/out4 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__360
       (.I0(\u2/u13/X [17]),
        .I1(\u2/u13/X [16]),
        .I2(\u2/u13/X [15]),
        .I3(\u2/u13/X [14]),
        .I4(\u2/u13/X [18]),
        .I5(\u2/u13/X [13]),
        .O(\u2/out13 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__361
       (.I0(\u2/u13/X [35]),
        .I1(\u2/u13/X [34]),
        .I2(\u2/u13/X [33]),
        .I3(\u2/u13/X [32]),
        .I4(\u2/u13/X [36]),
        .I5(\u2/u13/X [31]),
        .O(\u2/out13 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__362
       (.I0(\u2/u13/X [11]),
        .I1(\u2/u13/X [10]),
        .I2(\u2/u13/X [9]),
        .I3(\u2/u13/X [8]),
        .I4(\u2/u13/X [12]),
        .I5(\u2/u13/X [7]),
        .O(\u2/out13 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__363
       (.I0(\u2/u13/X [47]),
        .I1(\u2/u13/X [46]),
        .I2(\u2/u13/X [45]),
        .I3(\u2/u13/X [44]),
        .I4(\u2/u13/X [48]),
        .I5(\u2/u13/X [43]),
        .O(\u2/out13 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__364
       (.I0(\u2/u13/X [23]),
        .I1(\u2/u13/X [22]),
        .I2(\u2/u13/X [21]),
        .I3(\u2/u13/X [20]),
        .I4(\u2/u13/X [24]),
        .I5(\u2/u13/X [19]),
        .O(\u2/out13 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__365
       (.I0(\u2/u13/X [29]),
        .I1(\u2/u13/X [28]),
        .I2(\u2/u13/X [27]),
        .I3(\u2/u13/X [26]),
        .I4(\u2/u13/X [30]),
        .I5(\u2/u13/X [25]),
        .O(\u2/out13 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__366
       (.I0(\u2/u13/X [5]),
        .I1(\u2/u13/X [4]),
        .I2(\u2/u13/X [3]),
        .I3(\u2/u13/X [2]),
        .I4(\u2/u13/X [6]),
        .I5(\u2/u13/X [1]),
        .O(\u2/out13 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__367
       (.I0(\u2/u14/X [41]),
        .I1(\u2/u14/X [40]),
        .I2(\u2/u14/X [39]),
        .I3(\u2/u14/X [38]),
        .I4(\u2/u14/X [42]),
        .I5(\u2/u14/X [37]),
        .O(\u2/out14 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__368
       (.I0(\u2/u14/X [17]),
        .I1(\u2/u14/X [16]),
        .I2(\u2/u14/X [15]),
        .I3(\u2/u14/X [14]),
        .I4(\u2/u14/X [18]),
        .I5(\u2/u14/X [13]),
        .O(\u2/out14 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__369
       (.I0(\u2/u14/X [35]),
        .I1(\u2/u14/X [34]),
        .I2(\u2/u14/X [33]),
        .I3(\u2/u14/X [32]),
        .I4(\u2/u14/X [36]),
        .I5(\u2/u14/X [31]),
        .O(\u2/out14 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__37
       (.I0(\u0/u4/X [29]),
        .I1(\u0/u4/X [28]),
        .I2(\u0/u4/X [27]),
        .I3(\u0/u4/X [26]),
        .I4(\u0/u4/X [30]),
        .I5(\u0/u4/X [25]),
        .O(\u0/out4 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__370
       (.I0(\u2/u14/X [11]),
        .I1(\u2/u14/X [10]),
        .I2(\u2/u14/X [9]),
        .I3(\u2/u14/X [8]),
        .I4(\u2/u14/X [12]),
        .I5(\u2/u14/X [7]),
        .O(\u2/out14 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__371
       (.I0(\u2/u14/X [47]),
        .I1(\u2/u14/X [46]),
        .I2(\u2/u14/X [45]),
        .I3(\u2/u14/X [44]),
        .I4(\u2/u14/X [48]),
        .I5(\u2/u14/X [43]),
        .O(\u2/out14 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__372
       (.I0(\u2/u14/X [23]),
        .I1(\u2/u14/X [22]),
        .I2(\u2/u14/X [21]),
        .I3(\u2/u14/X [20]),
        .I4(\u2/u14/X [24]),
        .I5(\u2/u14/X [19]),
        .O(\u2/out14 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__373
       (.I0(\u2/u14/X [29]),
        .I1(\u2/u14/X [28]),
        .I2(\u2/u14/X [27]),
        .I3(\u2/u14/X [26]),
        .I4(\u2/u14/X [30]),
        .I5(\u2/u14/X [25]),
        .O(\u2/out14 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__374
       (.I0(\u2/u14/X [5]),
        .I1(\u2/u14/X [4]),
        .I2(\u2/u14/X [3]),
        .I3(\u2/u14/X [2]),
        .I4(\u2/u14/X [6]),
        .I5(\u2/u14/X [1]),
        .O(\u2/out14 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__375
       (.I0(\u2/u15/X [41]),
        .I1(\u2/u15/X [40]),
        .I2(\u2/u15/X [39]),
        .I3(\u2/u15/X [38]),
        .I4(\u2/u15/X [42]),
        .I5(\u2/u15/X [37]),
        .O(\u2/out15 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__376
       (.I0(\u2/u15/X [17]),
        .I1(\u2/u15/X [16]),
        .I2(\u2/u15/X [15]),
        .I3(\u2/u15/X [14]),
        .I4(\u2/u15/X [18]),
        .I5(\u2/u15/X [13]),
        .O(\u2/out15 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__377
       (.I0(\u2/u15/X [35]),
        .I1(\u2/u15/X [34]),
        .I2(\u2/u15/X [33]),
        .I3(\u2/u15/X [32]),
        .I4(\u2/u15/X [36]),
        .I5(\u2/u15/X [31]),
        .O(\u2/out15 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__378
       (.I0(\u2/u15/X [11]),
        .I1(\u2/u15/X [10]),
        .I2(\u2/u15/X [9]),
        .I3(\u2/u15/X [8]),
        .I4(\u2/u15/X [12]),
        .I5(\u2/u15/X [7]),
        .O(\u2/out15 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__379
       (.I0(\u2/u15/X [47]),
        .I1(\u2/u15/X [46]),
        .I2(\u2/u15/X [45]),
        .I3(\u2/u15/X [44]),
        .I4(\u2/u15/X [48]),
        .I5(\u2/u15/X [43]),
        .O(\u2/out15 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__38
       (.I0(\u0/u4/X [5]),
        .I1(\u0/u4/X [4]),
        .I2(\u0/u4/X [3]),
        .I3(\u0/u4/X [2]),
        .I4(\u0/u4/X [6]),
        .I5(\u0/u4/X [1]),
        .O(\u0/out4 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__380
       (.I0(\u2/u15/X [23]),
        .I1(\u2/u15/X [22]),
        .I2(\u2/u15/X [21]),
        .I3(\u2/u15/X [20]),
        .I4(\u2/u15/X [24]),
        .I5(\u2/u15/X [19]),
        .O(\u2/out15 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__381
       (.I0(\u2/u15/X [29]),
        .I1(\u2/u15/X [28]),
        .I2(\u2/u15/X [27]),
        .I3(\u2/u15/X [26]),
        .I4(\u2/u15/X [30]),
        .I5(\u2/u15/X [25]),
        .O(\u2/out15 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__382
       (.I0(\u2/u15/X [5]),
        .I1(\u2/u15/X [4]),
        .I2(\u2/u15/X [3]),
        .I3(\u2/u15/X [2]),
        .I4(\u2/u15/X [6]),
        .I5(\u2/u15/X [1]),
        .O(\u2/out15 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__39
       (.I0(\u0/u5/X [41]),
        .I1(\u0/u5/X [40]),
        .I2(\u0/u5/X [39]),
        .I3(\u0/u5/X [38]),
        .I4(\u0/u5/X [42]),
        .I5(\u0/u5/X [37]),
        .O(\u0/out5 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__4
       (.I0(\u0/u0/X [23]),
        .I1(\u0/u0/X [22]),
        .I2(\u0/u0/X [21]),
        .I3(\u0/u0/X [20]),
        .I4(\u0/u0/X [24]),
        .I5(\u0/u0/X [19]),
        .O(\u0/out0 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__40
       (.I0(\u0/u5/X [17]),
        .I1(\u0/u5/X [16]),
        .I2(\u0/u5/X [15]),
        .I3(\u0/u5/X [14]),
        .I4(\u0/u5/X [18]),
        .I5(\u0/u5/X [13]),
        .O(\u0/out5 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__41
       (.I0(\u0/u5/X [35]),
        .I1(\u0/u5/X [34]),
        .I2(\u0/u5/X [33]),
        .I3(\u0/u5/X [32]),
        .I4(\u0/u5/X [36]),
        .I5(\u0/u5/X [31]),
        .O(\u0/out5 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__42
       (.I0(\u0/u5/X [11]),
        .I1(\u0/u5/X [10]),
        .I2(\u0/u5/X [9]),
        .I3(\u0/u5/X [8]),
        .I4(\u0/u5/X [12]),
        .I5(\u0/u5/X [7]),
        .O(\u0/out5 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__43
       (.I0(\u0/u5/X [47]),
        .I1(\u0/u5/X [46]),
        .I2(\u0/u5/X [45]),
        .I3(\u0/u5/X [44]),
        .I4(\u0/u5/X [48]),
        .I5(\u0/u5/X [43]),
        .O(\u0/out5 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__44
       (.I0(\u0/u5/X [23]),
        .I1(\u0/u5/X [22]),
        .I2(\u0/u5/X [21]),
        .I3(\u0/u5/X [20]),
        .I4(\u0/u5/X [24]),
        .I5(\u0/u5/X [19]),
        .O(\u0/out5 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__45
       (.I0(\u0/u5/X [29]),
        .I1(\u0/u5/X [28]),
        .I2(\u0/u5/X [27]),
        .I3(\u0/u5/X [26]),
        .I4(\u0/u5/X [30]),
        .I5(\u0/u5/X [25]),
        .O(\u0/out5 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__46
       (.I0(\u0/u5/X [5]),
        .I1(\u0/u5/X [4]),
        .I2(\u0/u5/X [3]),
        .I3(\u0/u5/X [2]),
        .I4(\u0/u5/X [6]),
        .I5(\u0/u5/X [1]),
        .O(\u0/out5 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__47
       (.I0(\u0/u6/X [41]),
        .I1(\u0/u6/X [40]),
        .I2(\u0/u6/X [39]),
        .I3(\u0/u6/X [38]),
        .I4(\u0/u6/X [42]),
        .I5(\u0/u6/X [37]),
        .O(\u0/out6 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__48
       (.I0(\u0/u6/X [17]),
        .I1(\u0/u6/X [16]),
        .I2(\u0/u6/X [15]),
        .I3(\u0/u6/X [14]),
        .I4(\u0/u6/X [18]),
        .I5(\u0/u6/X [13]),
        .O(\u0/out6 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__49
       (.I0(\u0/u6/X [35]),
        .I1(\u0/u6/X [34]),
        .I2(\u0/u6/X [33]),
        .I3(\u0/u6/X [32]),
        .I4(\u0/u6/X [36]),
        .I5(\u0/u6/X [31]),
        .O(\u0/out6 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__5
       (.I0(\u0/u0/X [29]),
        .I1(\u0/u0/X [28]),
        .I2(\u0/u0/X [27]),
        .I3(\u0/u0/X [26]),
        .I4(\u0/u0/X [30]),
        .I5(\u0/u0/X [25]),
        .O(\u0/out0 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__50
       (.I0(\u0/u6/X [11]),
        .I1(\u0/u6/X [10]),
        .I2(\u0/u6/X [9]),
        .I3(\u0/u6/X [8]),
        .I4(\u0/u6/X [12]),
        .I5(\u0/u6/X [7]),
        .O(\u0/out6 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__51
       (.I0(\u0/u6/X [47]),
        .I1(\u0/u6/X [46]),
        .I2(\u0/u6/X [45]),
        .I3(\u0/u6/X [44]),
        .I4(\u0/u6/X [48]),
        .I5(\u0/u6/X [43]),
        .O(\u0/out6 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__52
       (.I0(\u0/u6/X [23]),
        .I1(\u0/u6/X [22]),
        .I2(\u0/u6/X [21]),
        .I3(\u0/u6/X [20]),
        .I4(\u0/u6/X [24]),
        .I5(\u0/u6/X [19]),
        .O(\u0/out6 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__53
       (.I0(\u0/u6/X [29]),
        .I1(\u0/u6/X [28]),
        .I2(\u0/u6/X [27]),
        .I3(\u0/u6/X [26]),
        .I4(\u0/u6/X [30]),
        .I5(\u0/u6/X [25]),
        .O(\u0/out6 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__54
       (.I0(\u0/u6/X [5]),
        .I1(\u0/u6/X [4]),
        .I2(\u0/u6/X [3]),
        .I3(\u0/u6/X [2]),
        .I4(\u0/u6/X [6]),
        .I5(\u0/u6/X [1]),
        .O(\u0/out6 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__55
       (.I0(\u0/u7/X [41]),
        .I1(\u0/u7/X [40]),
        .I2(\u0/u7/X [39]),
        .I3(\u0/u7/X [38]),
        .I4(\u0/u7/X [42]),
        .I5(\u0/u7/X [37]),
        .O(\u0/out7 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__56
       (.I0(\u0/u7/X [17]),
        .I1(\u0/u7/X [16]),
        .I2(\u0/u7/X [15]),
        .I3(\u0/u7/X [14]),
        .I4(\u0/u7/X [18]),
        .I5(\u0/u7/X [13]),
        .O(\u0/out7 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__57
       (.I0(\u0/u7/X [35]),
        .I1(\u0/u7/X [34]),
        .I2(\u0/u7/X [33]),
        .I3(\u0/u7/X [32]),
        .I4(\u0/u7/X [36]),
        .I5(\u0/u7/X [31]),
        .O(\u0/out7 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__58
       (.I0(\u0/u7/X [11]),
        .I1(\u0/u7/X [10]),
        .I2(\u0/u7/X [9]),
        .I3(\u0/u7/X [8]),
        .I4(\u0/u7/X [12]),
        .I5(\u0/u7/X [7]),
        .O(\u0/out7 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__59
       (.I0(\u0/u7/X [47]),
        .I1(\u0/u7/X [46]),
        .I2(\u0/u7/X [45]),
        .I3(\u0/u7/X [44]),
        .I4(\u0/u7/X [48]),
        .I5(\u0/u7/X [43]),
        .O(\u0/out7 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__6
       (.I0(\u0/u0/X [5]),
        .I1(\u0/u0/X [4]),
        .I2(\u0/u0/X [3]),
        .I3(\u0/u0/X [2]),
        .I4(\u0/u0/X [6]),
        .I5(\u0/u0/X [1]),
        .O(\u0/out0 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__60
       (.I0(\u0/u7/X [23]),
        .I1(\u0/u7/X [22]),
        .I2(\u0/u7/X [21]),
        .I3(\u0/u7/X [20]),
        .I4(\u0/u7/X [24]),
        .I5(\u0/u7/X [19]),
        .O(\u0/out7 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__61
       (.I0(\u0/u7/X [29]),
        .I1(\u0/u7/X [28]),
        .I2(\u0/u7/X [27]),
        .I3(\u0/u7/X [26]),
        .I4(\u0/u7/X [30]),
        .I5(\u0/u7/X [25]),
        .O(\u0/out7 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__62
       (.I0(\u0/u7/X [5]),
        .I1(\u0/u7/X [4]),
        .I2(\u0/u7/X [3]),
        .I3(\u0/u7/X [2]),
        .I4(\u0/u7/X [6]),
        .I5(\u0/u7/X [1]),
        .O(\u0/out7 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__63
       (.I0(\u0/u8/X [41]),
        .I1(\u0/u8/X [40]),
        .I2(\u0/u8/X [39]),
        .I3(\u0/u8/X [38]),
        .I4(\u0/u8/X [42]),
        .I5(\u0/u8/X [37]),
        .O(\u0/out8 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__64
       (.I0(\u0/u8/X [17]),
        .I1(\u0/u8/X [16]),
        .I2(\u0/u8/X [15]),
        .I3(\u0/u8/X [14]),
        .I4(\u0/u8/X [18]),
        .I5(\u0/u8/X [13]),
        .O(\u0/out8 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__65
       (.I0(\u0/u8/X [35]),
        .I1(\u0/u8/X [34]),
        .I2(\u0/u8/X [33]),
        .I3(\u0/u8/X [32]),
        .I4(\u0/u8/X [36]),
        .I5(\u0/u8/X [31]),
        .O(\u0/out8 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__66
       (.I0(\u0/u8/X [11]),
        .I1(\u0/u8/X [10]),
        .I2(\u0/u8/X [9]),
        .I3(\u0/u8/X [8]),
        .I4(\u0/u8/X [12]),
        .I5(\u0/u8/X [7]),
        .O(\u0/out8 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__67
       (.I0(\u0/u8/X [47]),
        .I1(\u0/u8/X [46]),
        .I2(\u0/u8/X [45]),
        .I3(\u0/u8/X [44]),
        .I4(\u0/u8/X [48]),
        .I5(\u0/u8/X [43]),
        .O(\u0/out8 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__68
       (.I0(\u0/u8/X [23]),
        .I1(\u0/u8/X [22]),
        .I2(\u0/u8/X [21]),
        .I3(\u0/u8/X [20]),
        .I4(\u0/u8/X [24]),
        .I5(\u0/u8/X [19]),
        .O(\u0/out8 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__69
       (.I0(\u0/u8/X [29]),
        .I1(\u0/u8/X [28]),
        .I2(\u0/u8/X [27]),
        .I3(\u0/u8/X [26]),
        .I4(\u0/u8/X [30]),
        .I5(\u0/u8/X [25]),
        .O(\u0/out8 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__7
       (.I0(\u0/u1/X [41]),
        .I1(\u0/u1/X [40]),
        .I2(\u0/u1/X [39]),
        .I3(\u0/u1/X [38]),
        .I4(\u0/u1/X [42]),
        .I5(\u0/u1/X [37]),
        .O(\u0/out1 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__70
       (.I0(\u0/u8/X [5]),
        .I1(\u0/u8/X [4]),
        .I2(\u0/u8/X [3]),
        .I3(\u0/u8/X [2]),
        .I4(\u0/u8/X [6]),
        .I5(\u0/u8/X [1]),
        .O(\u0/out8 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__71
       (.I0(\u0/u9/X [41]),
        .I1(\u0/u9/X [40]),
        .I2(\u0/u9/X [39]),
        .I3(\u0/u9/X [38]),
        .I4(\u0/u9/X [42]),
        .I5(\u0/u9/X [37]),
        .O(\u0/out9 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__72
       (.I0(\u0/u9/X [17]),
        .I1(\u0/u9/X [16]),
        .I2(\u0/u9/X [15]),
        .I3(\u0/u9/X [14]),
        .I4(\u0/u9/X [18]),
        .I5(\u0/u9/X [13]),
        .O(\u0/out9 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__73
       (.I0(\u0/u9/X [35]),
        .I1(\u0/u9/X [34]),
        .I2(\u0/u9/X [33]),
        .I3(\u0/u9/X [32]),
        .I4(\u0/u9/X [36]),
        .I5(\u0/u9/X [31]),
        .O(\u0/out9 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__74
       (.I0(\u0/u9/X [11]),
        .I1(\u0/u9/X [10]),
        .I2(\u0/u9/X [9]),
        .I3(\u0/u9/X [8]),
        .I4(\u0/u9/X [12]),
        .I5(\u0/u9/X [7]),
        .O(\u0/out9 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__75
       (.I0(\u0/u9/X [47]),
        .I1(\u0/u9/X [46]),
        .I2(\u0/u9/X [45]),
        .I3(\u0/u9/X [44]),
        .I4(\u0/u9/X [48]),
        .I5(\u0/u9/X [43]),
        .O(\u0/out9 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__76
       (.I0(\u0/u9/X [23]),
        .I1(\u0/u9/X [22]),
        .I2(\u0/u9/X [21]),
        .I3(\u0/u9/X [20]),
        .I4(\u0/u9/X [24]),
        .I5(\u0/u9/X [19]),
        .O(\u0/out9 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__77
       (.I0(\u0/u9/X [29]),
        .I1(\u0/u9/X [28]),
        .I2(\u0/u9/X [27]),
        .I3(\u0/u9/X [26]),
        .I4(\u0/u9/X [30]),
        .I5(\u0/u9/X [25]),
        .O(\u0/out9 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__78
       (.I0(\u0/u9/X [5]),
        .I1(\u0/u9/X [4]),
        .I2(\u0/u9/X [3]),
        .I3(\u0/u9/X [2]),
        .I4(\u0/u9/X [6]),
        .I5(\u0/u9/X [1]),
        .O(\u0/out9 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__79
       (.I0(\u0/u10/X [41]),
        .I1(\u0/u10/X [40]),
        .I2(\u0/u10/X [39]),
        .I3(\u0/u10/X [38]),
        .I4(\u0/u10/X [42]),
        .I5(\u0/u10/X [37]),
        .O(\u0/out10 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__8
       (.I0(\u0/u1/X [17]),
        .I1(\u0/u1/X [16]),
        .I2(\u0/u1/X [15]),
        .I3(\u0/u1/X [14]),
        .I4(\u0/u1/X [18]),
        .I5(\u0/u1/X [13]),
        .O(\u0/out1 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__80
       (.I0(\u0/u10/X [17]),
        .I1(\u0/u10/X [16]),
        .I2(\u0/u10/X [15]),
        .I3(\u0/u10/X [14]),
        .I4(\u0/u10/X [18]),
        .I5(\u0/u10/X [13]),
        .O(\u0/out10 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__81
       (.I0(\u0/u10/X [35]),
        .I1(\u0/u10/X [34]),
        .I2(\u0/u10/X [33]),
        .I3(\u0/u10/X [32]),
        .I4(\u0/u10/X [36]),
        .I5(\u0/u10/X [31]),
        .O(\u0/out10 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__82
       (.I0(\u0/u10/X [11]),
        .I1(\u0/u10/X [10]),
        .I2(\u0/u10/X [9]),
        .I3(\u0/u10/X [8]),
        .I4(\u0/u10/X [12]),
        .I5(\u0/u10/X [7]),
        .O(\u0/out10 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__83
       (.I0(\u0/u10/X [47]),
        .I1(\u0/u10/X [46]),
        .I2(\u0/u10/X [45]),
        .I3(\u0/u10/X [44]),
        .I4(\u0/u10/X [48]),
        .I5(\u0/u10/X [43]),
        .O(\u0/out10 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__84
       (.I0(\u0/u10/X [23]),
        .I1(\u0/u10/X [22]),
        .I2(\u0/u10/X [21]),
        .I3(\u0/u10/X [20]),
        .I4(\u0/u10/X [24]),
        .I5(\u0/u10/X [19]),
        .O(\u0/out10 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__85
       (.I0(\u0/u10/X [29]),
        .I1(\u0/u10/X [28]),
        .I2(\u0/u10/X [27]),
        .I3(\u0/u10/X [26]),
        .I4(\u0/u10/X [30]),
        .I5(\u0/u10/X [25]),
        .O(\u0/out10 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__86
       (.I0(\u0/u10/X [5]),
        .I1(\u0/u10/X [4]),
        .I2(\u0/u10/X [3]),
        .I3(\u0/u10/X [2]),
        .I4(\u0/u10/X [6]),
        .I5(\u0/u10/X [1]),
        .O(\u0/out10 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__87
       (.I0(\u0/u11/X [41]),
        .I1(\u0/u11/X [40]),
        .I2(\u0/u11/X [39]),
        .I3(\u0/u11/X [38]),
        .I4(\u0/u11/X [42]),
        .I5(\u0/u11/X [37]),
        .O(\u0/out11 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__88
       (.I0(\u0/u11/X [17]),
        .I1(\u0/u11/X [16]),
        .I2(\u0/u11/X [15]),
        .I3(\u0/u11/X [14]),
        .I4(\u0/u11/X [18]),
        .I5(\u0/u11/X [13]),
        .O(\u0/out11 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__89
       (.I0(\u0/u11/X [35]),
        .I1(\u0/u11/X [34]),
        .I2(\u0/u11/X [33]),
        .I3(\u0/u11/X [32]),
        .I4(\u0/u11/X [36]),
        .I5(\u0/u11/X [31]),
        .O(\u0/out11 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__9
       (.I0(\u0/u1/X [35]),
        .I1(\u0/u1/X [34]),
        .I2(\u0/u1/X [33]),
        .I3(\u0/u1/X [32]),
        .I4(\u0/u1/X [36]),
        .I5(\u0/u1/X [31]),
        .O(\u0/out1 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__90
       (.I0(\u0/u11/X [11]),
        .I1(\u0/u11/X [10]),
        .I2(\u0/u11/X [9]),
        .I3(\u0/u11/X [8]),
        .I4(\u0/u11/X [12]),
        .I5(\u0/u11/X [7]),
        .O(\u0/out11 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__91
       (.I0(\u0/u11/X [47]),
        .I1(\u0/u11/X [46]),
        .I2(\u0/u11/X [45]),
        .I3(\u0/u11/X [44]),
        .I4(\u0/u11/X [48]),
        .I5(\u0/u11/X [43]),
        .O(\u0/out11 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h99D249B5E827B4C6)) 
    g0_b3__92
       (.I0(\u0/u11/X [23]),
        .I1(\u0/u11/X [22]),
        .I2(\u0/u11/X [21]),
        .I3(\u0/u11/X [20]),
        .I4(\u0/u11/X [24]),
        .I5(\u0/u11/X [19]),
        .O(\u0/out11 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1AA787B86C4BD962)) 
    g0_b3__93
       (.I0(\u0/u11/X [29]),
        .I1(\u0/u11/X [28]),
        .I2(\u0/u11/X [27]),
        .I3(\u0/u11/X [26]),
        .I4(\u0/u11/X [30]),
        .I5(\u0/u11/X [25]),
        .O(\u0/out11 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9A27279C9D522AE5)) 
    g0_b3__94
       (.I0(\u0/u11/X [5]),
        .I1(\u0/u11/X [4]),
        .I2(\u0/u11/X [3]),
        .I3(\u0/u11/X [2]),
        .I4(\u0/u11/X [6]),
        .I5(\u0/u11/X [1]),
        .O(\u0/out11 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h994E4B9C69A526DA)) 
    g0_b3__95
       (.I0(\u0/u12/X [41]),
        .I1(\u0/u12/X [40]),
        .I2(\u0/u12/X [39]),
        .I3(\u0/u12/X [38]),
        .I4(\u0/u12/X [42]),
        .I5(\u0/u12/X [37]),
        .O(\u0/out12 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h966669397A89964D)) 
    g0_b3__96
       (.I0(\u0/u12/X [17]),
        .I1(\u0/u12/X [16]),
        .I2(\u0/u12/X [15]),
        .I3(\u0/u12/X [14]),
        .I4(\u0/u12/X [18]),
        .I5(\u0/u12/X [13]),
        .O(\u0/out12 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC3D86867AC63929D)) 
    g0_b3__97
       (.I0(\u0/u12/X [35]),
        .I1(\u0/u12/X [34]),
        .I2(\u0/u12/X [33]),
        .I3(\u0/u12/X [32]),
        .I4(\u0/u12/X [36]),
        .I5(\u0/u12/X [31]),
        .O(\u0/out12 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC927965A69D2992D)) 
    g0_b3__98
       (.I0(\u0/u12/X [11]),
        .I1(\u0/u12/X [10]),
        .I2(\u0/u12/X [9]),
        .I3(\u0/u12/X [8]),
        .I4(\u0/u12/X [12]),
        .I5(\u0/u12/X [7]),
        .O(\u0/out12 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87E49C72691E4B65)) 
    g0_b3__99
       (.I0(\u0/u12/X [47]),
        .I1(\u0/u12/X [46]),
        .I2(\u0/u12/X [45]),
        .I3(\u0/u12/X [44]),
        .I4(\u0/u12/X [48]),
        .I5(\u0/u12/X [43]),
        .O(\u0/out12 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[0]),
        .Q(key_b_r_reg_n_0_),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[10]),
        .Q(\key_b_r_reg_n_0_[0][10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[11]),
        .Q(\key_b_r_reg_n_0_[0][11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[12]),
        .Q(\key_b_r_reg_n_0_[0][12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[13]),
        .Q(\key_b_r_reg_n_0_[0][13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[14]),
        .Q(\key_b_r_reg_n_0_[0][14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[15]),
        .Q(\key_b_r_reg_n_0_[0][15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[16]),
        .Q(\key_b_r_reg_n_0_[0][16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[17]),
        .Q(\key_b_r_reg_n_0_[0][17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[18]),
        .Q(\key_b_r_reg_n_0_[0][18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[19]),
        .Q(\key_b_r_reg_n_0_[0][19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[1]),
        .Q(\key_b_r_reg_n_0_[0][1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[20]),
        .Q(\key_b_r_reg_n_0_[0][20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[21]),
        .Q(\key_b_r_reg_n_0_[0][21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[22]),
        .Q(\key_b_r_reg_n_0_[0][22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[23]),
        .Q(\key_b_r_reg_n_0_[0][23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[24]),
        .Q(\key_b_r_reg_n_0_[0][24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[25]),
        .Q(\key_b_r_reg_n_0_[0][25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[26]),
        .Q(\key_b_r_reg_n_0_[0][26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[27]),
        .Q(\key_b_r_reg_n_0_[0][27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[28]),
        .Q(\key_b_r_reg_n_0_[0][28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[29]),
        .Q(\key_b_r_reg_n_0_[0][29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[2]),
        .Q(\key_b_r_reg_n_0_[0][2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[30]),
        .Q(\key_b_r_reg_n_0_[0][30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[31]),
        .Q(\key_b_r_reg_n_0_[0][31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[32]),
        .Q(\key_b_r_reg_n_0_[0][32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[33]),
        .Q(\key_b_r_reg_n_0_[0][33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[34]),
        .Q(\key_b_r_reg_n_0_[0][34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[35]),
        .Q(\key_b_r_reg_n_0_[0][35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[36]),
        .Q(\key_b_r_reg_n_0_[0][36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[37]),
        .Q(\key_b_r_reg_n_0_[0][37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[38]),
        .Q(\key_b_r_reg_n_0_[0][38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[39]),
        .Q(\key_b_r_reg_n_0_[0][39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[3]),
        .Q(\key_b_r_reg_n_0_[0][3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[40]),
        .Q(\key_b_r_reg_n_0_[0][40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[41]),
        .Q(\key_b_r_reg_n_0_[0][41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[42]),
        .Q(\key_b_r_reg_n_0_[0][42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[43]),
        .Q(\key_b_r_reg_n_0_[0][43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[44]),
        .Q(\key_b_r_reg_n_0_[0][44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[45]),
        .Q(\key_b_r_reg_n_0_[0][45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[46]),
        .Q(\key_b_r_reg_n_0_[0][46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[47]),
        .Q(\key_b_r_reg_n_0_[0][47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[48]),
        .Q(\key_b_r_reg_n_0_[0][48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[49]),
        .Q(\key_b_r_reg_n_0_[0][49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[4]),
        .Q(\key_b_r_reg_n_0_[0][4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[50]),
        .Q(\key_b_r_reg_n_0_[0][50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[51]),
        .Q(\key_b_r_reg_n_0_[0][51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[52]),
        .Q(\key_b_r_reg_n_0_[0][52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[53]),
        .Q(\key_b_r_reg_n_0_[0][53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[54]),
        .Q(\key_b_r_reg_n_0_[0][54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[55]),
        .Q(\key_b_r_reg_n_0_[0][55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[5]),
        .Q(\key_b_r_reg_n_0_[0][5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[6]),
        .Q(\key_b_r_reg_n_0_[0][6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[7]),
        .Q(\key_b_r_reg_n_0_[0][7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[8]),
        .Q(\key_b_r_reg_n_0_[0][8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \key_b_r_reg[0][9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key2[9]),
        .Q(\key_b_r_reg_n_0_[0][9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][0]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][0]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_b_r_reg_n_0_),
        .Q(key_b_r_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][10]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][10]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][10] ),
        .Q(\key_b_r_reg[16][10]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][11]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][11]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][11] ),
        .Q(\key_b_r_reg[16][11]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][12]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][12]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][12] ),
        .Q(\key_b_r_reg[16][12]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][13]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][13]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][13] ),
        .Q(\key_b_r_reg[16][13]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][14]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][14]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][14] ),
        .Q(\key_b_r_reg[16][14]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][15]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][15]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][15] ),
        .Q(\key_b_r_reg[16][15]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][16]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][16]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][16] ),
        .Q(\key_b_r_reg[16][16]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][17]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][17]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][17] ),
        .Q(\key_b_r_reg[16][17]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][18]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][18]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][18] ),
        .Q(\key_b_r_reg[16][18]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][19]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][19]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][19] ),
        .Q(\key_b_r_reg[16][19]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][1]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][1]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][1] ),
        .Q(\key_b_r_reg[16][1]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][20]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][20]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][20] ),
        .Q(\key_b_r_reg[16][20]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][21]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][21]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][21] ),
        .Q(\key_b_r_reg[16][21]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][22]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][22]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][22] ),
        .Q(\key_b_r_reg[16][22]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][23]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][23]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][23] ),
        .Q(\key_b_r_reg[16][23]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][24]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][24]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][24] ),
        .Q(\key_b_r_reg[16][24]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][25]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][25]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][25] ),
        .Q(\key_b_r_reg[16][25]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][26]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][26]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][26] ),
        .Q(\key_b_r_reg[16][26]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][27]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][27]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][27] ),
        .Q(\key_b_r_reg[16][27]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][28]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][28]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][28] ),
        .Q(\key_b_r_reg[16][28]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][29]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][29]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][29] ),
        .Q(\key_b_r_reg[16][29]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][2]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][2]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][2] ),
        .Q(\key_b_r_reg[16][2]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][30]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][30]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][30] ),
        .Q(\key_b_r_reg[16][30]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][31]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][31]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][31] ),
        .Q(\key_b_r_reg[16][31]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][32]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][32]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][32] ),
        .Q(\key_b_r_reg[16][32]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][33]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][33]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][33] ),
        .Q(\key_b_r_reg[16][33]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][34]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][34]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][34] ),
        .Q(\key_b_r_reg[16][34]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][35]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][35]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][35] ),
        .Q(\key_b_r_reg[16][35]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][36]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][36]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][36] ),
        .Q(\key_b_r_reg[16][36]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][37]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][37]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][37] ),
        .Q(\key_b_r_reg[16][37]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][38]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][38]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][38] ),
        .Q(\key_b_r_reg[16][38]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][39]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][39]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][39] ),
        .Q(\key_b_r_reg[16][39]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][3]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][3]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][3] ),
        .Q(\key_b_r_reg[16][3]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][40]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][40]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][40] ),
        .Q(\key_b_r_reg[16][40]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][41]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][41]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][41] ),
        .Q(\key_b_r_reg[16][41]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][42]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][42]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][42] ),
        .Q(\key_b_r_reg[16][42]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][43]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][43]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][43] ),
        .Q(\key_b_r_reg[16][43]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][44]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][44]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][44] ),
        .Q(\key_b_r_reg[16][44]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][45]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][45]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][45] ),
        .Q(\key_b_r_reg[16][45]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][46]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][46]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][46] ),
        .Q(\key_b_r_reg[16][46]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][47]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][47]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][47] ),
        .Q(\key_b_r_reg[16][47]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][48]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][48]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][48] ),
        .Q(\key_b_r_reg[16][48]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][49]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][49]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][49] ),
        .Q(\key_b_r_reg[16][49]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][4]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][4]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][4] ),
        .Q(\key_b_r_reg[16][4]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][50]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][50]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][50] ),
        .Q(\key_b_r_reg[16][50]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][51]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][51]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][51] ),
        .Q(\key_b_r_reg[16][51]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][52]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][52]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][52] ),
        .Q(\key_b_r_reg[16][52]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][53]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][53]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][53] ),
        .Q(\key_b_r_reg[16][53]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][54]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][54]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][54] ),
        .Q(\key_b_r_reg[16][54]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][55]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][55]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][55] ),
        .Q(\key_b_r_reg[16][55]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][5]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][5]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][5] ),
        .Q(\key_b_r_reg[16][5]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][6]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][6]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][6] ),
        .Q(\key_b_r_reg[16][6]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][7]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][7]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][7] ),
        .Q(\key_b_r_reg[16][7]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][8]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][8]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][8] ),
        .Q(\key_b_r_reg[16][8]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_b_r_reg[16] " *) 
  (* srl_name = "des3_perf_0/\key_b_r_reg[16][9]_srl16 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_b_r_reg[16][9]_srl16 
       (.A0(\<const1>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const1>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_b_r_reg_n_0_[0][9] ),
        .Q(\key_b_r_reg[16][9]_srl16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][0]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][0]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[0]),
        .Q31(key_c_r_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][0]_srl32_i_1 
       (.I0(key1[0]),
        .I1(key3[0]),
        .I2(decrypt),
        .O(key_c[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][10]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][10]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[10]),
        .Q31(\key_c_r_reg[31][10]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][10]_srl32_i_1 
       (.I0(key1[10]),
        .I1(key3[10]),
        .I2(decrypt),
        .O(key_c[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][11]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][11]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[11]),
        .Q31(\key_c_r_reg[31][11]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][11]_srl32_i_1 
       (.I0(key1[11]),
        .I1(key3[11]),
        .I2(decrypt),
        .O(key_c[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][12]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][12]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[12]),
        .Q31(\key_c_r_reg[31][12]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][12]_srl32_i_1 
       (.I0(key1[12]),
        .I1(key3[12]),
        .I2(decrypt),
        .O(key_c[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][13]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][13]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[13]),
        .Q31(\key_c_r_reg[31][13]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][13]_srl32_i_1 
       (.I0(key1[13]),
        .I1(key3[13]),
        .I2(decrypt),
        .O(key_c[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][14]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][14]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[14]),
        .Q31(\key_c_r_reg[31][14]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][14]_srl32_i_1 
       (.I0(key1[14]),
        .I1(key3[14]),
        .I2(decrypt),
        .O(key_c[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][15]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][15]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[15]),
        .Q31(\key_c_r_reg[31][15]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][15]_srl32_i_1 
       (.I0(key1[15]),
        .I1(key3[15]),
        .I2(decrypt),
        .O(key_c[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][16]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][16]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[16]),
        .Q31(\key_c_r_reg[31][16]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][16]_srl32_i_1 
       (.I0(key1[16]),
        .I1(key3[16]),
        .I2(decrypt),
        .O(key_c[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][17]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][17]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[17]),
        .Q31(\key_c_r_reg[31][17]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][17]_srl32_i_1 
       (.I0(key1[17]),
        .I1(key3[17]),
        .I2(decrypt),
        .O(key_c[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][18]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][18]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[18]),
        .Q31(\key_c_r_reg[31][18]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][18]_srl32_i_1 
       (.I0(key1[18]),
        .I1(key3[18]),
        .I2(decrypt),
        .O(key_c[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][19]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][19]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[19]),
        .Q31(\key_c_r_reg[31][19]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][19]_srl32_i_1 
       (.I0(key1[19]),
        .I1(key3[19]),
        .I2(decrypt),
        .O(key_c[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][1]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][1]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[1]),
        .Q31(\key_c_r_reg[31][1]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][1]_srl32_i_1 
       (.I0(key1[1]),
        .I1(key3[1]),
        .I2(decrypt),
        .O(key_c[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][20]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][20]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[20]),
        .Q31(\key_c_r_reg[31][20]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][20]_srl32_i_1 
       (.I0(key1[20]),
        .I1(key3[20]),
        .I2(decrypt),
        .O(key_c[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][21]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][21]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[21]),
        .Q31(\key_c_r_reg[31][21]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][21]_srl32_i_1 
       (.I0(key1[21]),
        .I1(key3[21]),
        .I2(decrypt),
        .O(key_c[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][22]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][22]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[22]),
        .Q31(\key_c_r_reg[31][22]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][22]_srl32_i_1 
       (.I0(key1[22]),
        .I1(key3[22]),
        .I2(decrypt),
        .O(key_c[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][23]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][23]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[23]),
        .Q31(\key_c_r_reg[31][23]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][23]_srl32_i_1 
       (.I0(key1[23]),
        .I1(key3[23]),
        .I2(decrypt),
        .O(key_c[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][24]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][24]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[24]),
        .Q31(\key_c_r_reg[31][24]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][24]_srl32_i_1 
       (.I0(key1[24]),
        .I1(key3[24]),
        .I2(decrypt),
        .O(key_c[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][25]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][25]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[25]),
        .Q31(\key_c_r_reg[31][25]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][25]_srl32_i_1 
       (.I0(key1[25]),
        .I1(key3[25]),
        .I2(decrypt),
        .O(key_c[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][26]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][26]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[26]),
        .Q31(\key_c_r_reg[31][26]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][26]_srl32_i_1 
       (.I0(key1[26]),
        .I1(key3[26]),
        .I2(decrypt),
        .O(key_c[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][27]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][27]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[27]),
        .Q31(\key_c_r_reg[31][27]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][27]_srl32_i_1 
       (.I0(key1[27]),
        .I1(key3[27]),
        .I2(decrypt),
        .O(key_c[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][28]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][28]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[28]),
        .Q31(\key_c_r_reg[31][28]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][28]_srl32_i_1 
       (.I0(key1[28]),
        .I1(key3[28]),
        .I2(decrypt),
        .O(key_c[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][29]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][29]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[29]),
        .Q31(\key_c_r_reg[31][29]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][29]_srl32_i_1 
       (.I0(key1[29]),
        .I1(key3[29]),
        .I2(decrypt),
        .O(key_c[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][2]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][2]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[2]),
        .Q31(\key_c_r_reg[31][2]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][2]_srl32_i_1 
       (.I0(key1[2]),
        .I1(key3[2]),
        .I2(decrypt),
        .O(key_c[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][30]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][30]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[30]),
        .Q31(\key_c_r_reg[31][30]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][30]_srl32_i_1 
       (.I0(key1[30]),
        .I1(key3[30]),
        .I2(decrypt),
        .O(key_c[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][31]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][31]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[31]),
        .Q31(\key_c_r_reg[31][31]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][31]_srl32_i_1 
       (.I0(key1[31]),
        .I1(key3[31]),
        .I2(decrypt),
        .O(key_c[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][32]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][32]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[32]),
        .Q31(\key_c_r_reg[31][32]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][32]_srl32_i_1 
       (.I0(key1[32]),
        .I1(key3[32]),
        .I2(decrypt),
        .O(key_c[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][33]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][33]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[33]),
        .Q31(\key_c_r_reg[31][33]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][33]_srl32_i_1 
       (.I0(key1[33]),
        .I1(key3[33]),
        .I2(decrypt),
        .O(key_c[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][34]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][34]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[34]),
        .Q31(\key_c_r_reg[31][34]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][34]_srl32_i_1 
       (.I0(key1[34]),
        .I1(key3[34]),
        .I2(decrypt),
        .O(key_c[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][35]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][35]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[35]),
        .Q31(\key_c_r_reg[31][35]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][35]_srl32_i_1 
       (.I0(key1[35]),
        .I1(key3[35]),
        .I2(decrypt),
        .O(key_c[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][36]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][36]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[36]),
        .Q31(\key_c_r_reg[31][36]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][36]_srl32_i_1 
       (.I0(key1[36]),
        .I1(key3[36]),
        .I2(decrypt),
        .O(key_c[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][37]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][37]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[37]),
        .Q31(\key_c_r_reg[31][37]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][37]_srl32_i_1 
       (.I0(key1[37]),
        .I1(key3[37]),
        .I2(decrypt),
        .O(key_c[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][38]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][38]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[38]),
        .Q31(\key_c_r_reg[31][38]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][38]_srl32_i_1 
       (.I0(key1[38]),
        .I1(key3[38]),
        .I2(decrypt),
        .O(key_c[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][39]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][39]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[39]),
        .Q31(\key_c_r_reg[31][39]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][39]_srl32_i_1 
       (.I0(key1[39]),
        .I1(key3[39]),
        .I2(decrypt),
        .O(key_c[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][3]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][3]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[3]),
        .Q31(\key_c_r_reg[31][3]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][3]_srl32_i_1 
       (.I0(key1[3]),
        .I1(key3[3]),
        .I2(decrypt),
        .O(key_c[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][40]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][40]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[40]),
        .Q31(\key_c_r_reg[31][40]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][40]_srl32_i_1 
       (.I0(key1[40]),
        .I1(key3[40]),
        .I2(decrypt),
        .O(key_c[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][41]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][41]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[41]),
        .Q31(\key_c_r_reg[31][41]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][41]_srl32_i_1 
       (.I0(key1[41]),
        .I1(key3[41]),
        .I2(decrypt),
        .O(key_c[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][42]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][42]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[42]),
        .Q31(\key_c_r_reg[31][42]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][42]_srl32_i_1 
       (.I0(key1[42]),
        .I1(key3[42]),
        .I2(decrypt),
        .O(key_c[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][43]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][43]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[43]),
        .Q31(\key_c_r_reg[31][43]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][43]_srl32_i_1 
       (.I0(key1[43]),
        .I1(key3[43]),
        .I2(decrypt),
        .O(key_c[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][44]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][44]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[44]),
        .Q31(\key_c_r_reg[31][44]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][44]_srl32_i_1 
       (.I0(key1[44]),
        .I1(key3[44]),
        .I2(decrypt),
        .O(key_c[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][45]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][45]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[45]),
        .Q31(\key_c_r_reg[31][45]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][45]_srl32_i_1 
       (.I0(key1[45]),
        .I1(key3[45]),
        .I2(decrypt),
        .O(key_c[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][46]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][46]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[46]),
        .Q31(\key_c_r_reg[31][46]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][46]_srl32_i_1 
       (.I0(key1[46]),
        .I1(key3[46]),
        .I2(decrypt),
        .O(key_c[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][47]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][47]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[47]),
        .Q31(\key_c_r_reg[31][47]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][47]_srl32_i_1 
       (.I0(key1[47]),
        .I1(key3[47]),
        .I2(decrypt),
        .O(key_c[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][48]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][48]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[48]),
        .Q31(\key_c_r_reg[31][48]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][48]_srl32_i_1 
       (.I0(key1[48]),
        .I1(key3[48]),
        .I2(decrypt),
        .O(key_c[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][49]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][49]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[49]),
        .Q31(\key_c_r_reg[31][49]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][49]_srl32_i_1 
       (.I0(key1[49]),
        .I1(key3[49]),
        .I2(decrypt),
        .O(key_c[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][4]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][4]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[4]),
        .Q31(\key_c_r_reg[31][4]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][4]_srl32_i_1 
       (.I0(key1[4]),
        .I1(key3[4]),
        .I2(decrypt),
        .O(key_c[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][50]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][50]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[50]),
        .Q31(\key_c_r_reg[31][50]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][50]_srl32_i_1 
       (.I0(key1[50]),
        .I1(key3[50]),
        .I2(decrypt),
        .O(key_c[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][51]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][51]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[51]),
        .Q31(\key_c_r_reg[31][51]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][51]_srl32_i_1 
       (.I0(key1[51]),
        .I1(key3[51]),
        .I2(decrypt),
        .O(key_c[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][52]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][52]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[52]),
        .Q31(\key_c_r_reg[31][52]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][52]_srl32_i_1 
       (.I0(key1[52]),
        .I1(key3[52]),
        .I2(decrypt),
        .O(key_c[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][53]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][53]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[53]),
        .Q31(\key_c_r_reg[31][53]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][53]_srl32_i_1 
       (.I0(key1[53]),
        .I1(key3[53]),
        .I2(decrypt),
        .O(key_c[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][54]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][54]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[54]),
        .Q31(\key_c_r_reg[31][54]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][54]_srl32_i_1 
       (.I0(key1[54]),
        .I1(key3[54]),
        .I2(decrypt),
        .O(key_c[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][55]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][55]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[55]),
        .Q31(\key_c_r_reg[31][55]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][55]_srl32_i_1 
       (.I0(key1[55]),
        .I1(key3[55]),
        .I2(decrypt),
        .O(key_c[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][5]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][5]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[5]),
        .Q31(\key_c_r_reg[31][5]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][5]_srl32_i_1 
       (.I0(key1[5]),
        .I1(key3[5]),
        .I2(decrypt),
        .O(key_c[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][6]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][6]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[6]),
        .Q31(\key_c_r_reg[31][6]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][6]_srl32_i_1 
       (.I0(key1[6]),
        .I1(key3[6]),
        .I2(decrypt),
        .O(key_c[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][7]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][7]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[7]),
        .Q31(\key_c_r_reg[31][7]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][7]_srl32_i_1 
       (.I0(key1[7]),
        .I1(key3[7]),
        .I2(decrypt),
        .O(key_c[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][8]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][8]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[8]),
        .Q31(\key_c_r_reg[31][8]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][8]_srl32_i_1 
       (.I0(key1[8]),
        .I1(key3[8]),
        .I2(decrypt),
        .O(key_c[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[31] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[31][9]_srl32 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[31][9]_srl32 
       (.A({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c[9]),
        .Q31(\key_c_r_reg[31][9]_srl32_n_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_c_r_reg[31][9]_srl32_i_1 
       (.I0(key1[9]),
        .I1(key3[9]),
        .I2(decrypt),
        .O(key_c[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][0]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][0]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(key_c_r_reg),
        .Q(\key_c_r_reg[33][0]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][10]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][10]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][10]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][10]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][11]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][11]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][11]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][11]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][12]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][12]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][12]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][12]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][13]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][13]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][13]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][13]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][14]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][14]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][14]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][14]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][15]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][15]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][15]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][15]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][16]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][16]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][16]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][16]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][17]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][17]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][17]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][17]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][18]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][18]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][18]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][18]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][19]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][19]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][19]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][19]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][1]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][1]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][1]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][1]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][20]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][20]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][20]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][20]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][21]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][21]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][21]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][21]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][22]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][22]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][22]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][22]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][23]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][23]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][23]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][23]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][24]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][24]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][24]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][24]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][25]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][25]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][25]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][25]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][26]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][26]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][26]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][26]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][27]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][27]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][27]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][27]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][28]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][28]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][28]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][28]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][29]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][29]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][29]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][29]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][2]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][2]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][2]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][2]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][30]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][30]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][30]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][30]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][31]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][31]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][31]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][31]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][32]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][32]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][32]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][32]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][33]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][33]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][33]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][33]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][34]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][34]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][34]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][34]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][35]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][35]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][35]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][35]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][36]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][36]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][36]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][36]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][37]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][37]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][37]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][37]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][38]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][38]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][38]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][38]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][39]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][39]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][39]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][39]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][3]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][3]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][3]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][3]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][40]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][40]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][40]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][40]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][41]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][41]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][41]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][41]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][42]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][42]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][42]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][42]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][43]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][43]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][43]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][43]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][44]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][44]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][44]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][44]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][45]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][45]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][45]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][45]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][46]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][46]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][46]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][46]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][47]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][47]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][47]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][47]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][48]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][48]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][48]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][48]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][49]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][49]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][49]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][49]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][4]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][4]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][4]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][4]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][50]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][50]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][50]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][50]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][51]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][51]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][51]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][51]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][52]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][52]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][52]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][52]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][53]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][53]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][53]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][53]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][54]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][54]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][54]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][54]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][55]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][55]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][55]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][55]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][5]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][5]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][5]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][5]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][6]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][6]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][6]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][6]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][7]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][7]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][7]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][7]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][8]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][8]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][8]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][8]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "SRLC32E" *) 
  (* srl_bus_name = "des3_perf_0/\key_c_r_reg[33] " *) 
  (* srl_name = "des3_perf_0/\key_c_r_reg[33][9]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \key_c_r_reg[33][9]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(\key_c_r_reg[31][9]_srl32_n_1 ),
        .Q(\key_c_r_reg[33][9]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[0]_i_1 
       (.I0(key3[0]),
        .I1(key1[0]),
        .I2(decrypt),
        .O(key_a[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[10]_i_1 
       (.I0(key3[10]),
        .I1(key1[10]),
        .I2(decrypt),
        .O(key_a[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[11]_i_1 
       (.I0(key3[11]),
        .I1(key1[11]),
        .I2(decrypt),
        .O(key_a[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[12]_i_1 
       (.I0(key3[12]),
        .I1(key1[12]),
        .I2(decrypt),
        .O(key_a[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[13]_i_1 
       (.I0(key3[13]),
        .I1(key1[13]),
        .I2(decrypt),
        .O(key_a[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[14]_i_1 
       (.I0(key3[14]),
        .I1(key1[14]),
        .I2(decrypt),
        .O(key_a[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[15]_i_1 
       (.I0(key3[15]),
        .I1(key1[15]),
        .I2(decrypt),
        .O(key_a[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[16]_i_1 
       (.I0(key3[16]),
        .I1(key1[16]),
        .I2(decrypt),
        .O(key_a[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[17]_i_1 
       (.I0(key3[17]),
        .I1(key1[17]),
        .I2(decrypt),
        .O(key_a[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[18]_i_1 
       (.I0(key3[18]),
        .I1(key1[18]),
        .I2(decrypt),
        .O(key_a[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[19]_i_1 
       (.I0(key3[19]),
        .I1(key1[19]),
        .I2(decrypt),
        .O(key_a[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[1]_i_1 
       (.I0(key3[1]),
        .I1(key1[1]),
        .I2(decrypt),
        .O(key_a[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[20]_i_1 
       (.I0(key3[20]),
        .I1(key1[20]),
        .I2(decrypt),
        .O(key_a[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[21]_i_1 
       (.I0(key3[21]),
        .I1(key1[21]),
        .I2(decrypt),
        .O(key_a[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[22]_i_1 
       (.I0(key3[22]),
        .I1(key1[22]),
        .I2(decrypt),
        .O(key_a[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[23]_i_1 
       (.I0(key3[23]),
        .I1(key1[23]),
        .I2(decrypt),
        .O(key_a[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[24]_i_1 
       (.I0(key3[24]),
        .I1(key1[24]),
        .I2(decrypt),
        .O(key_a[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[25]_i_1 
       (.I0(key3[25]),
        .I1(key1[25]),
        .I2(decrypt),
        .O(key_a[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[26]_i_1 
       (.I0(key3[26]),
        .I1(key1[26]),
        .I2(decrypt),
        .O(key_a[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[27]_i_1 
       (.I0(key3[27]),
        .I1(key1[27]),
        .I2(decrypt),
        .O(key_a[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[28]_i_1 
       (.I0(key3[28]),
        .I1(key1[28]),
        .I2(decrypt),
        .O(key_a[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[29]_i_1 
       (.I0(key3[29]),
        .I1(key1[29]),
        .I2(decrypt),
        .O(key_a[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[2]_i_1 
       (.I0(key3[2]),
        .I1(key1[2]),
        .I2(decrypt),
        .O(key_a[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[30]_i_1 
       (.I0(key3[30]),
        .I1(key1[30]),
        .I2(decrypt),
        .O(key_a[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[31]_i_1 
       (.I0(key3[31]),
        .I1(key1[31]),
        .I2(decrypt),
        .O(key_a[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[32]_i_1 
       (.I0(key3[32]),
        .I1(key1[32]),
        .I2(decrypt),
        .O(key_a[32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[33]_i_1 
       (.I0(key3[33]),
        .I1(key1[33]),
        .I2(decrypt),
        .O(key_a[33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[34]_i_1 
       (.I0(key3[34]),
        .I1(key1[34]),
        .I2(decrypt),
        .O(key_a[34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[35]_i_1 
       (.I0(key3[35]),
        .I1(key1[35]),
        .I2(decrypt),
        .O(key_a[35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[36]_i_1 
       (.I0(key3[36]),
        .I1(key1[36]),
        .I2(decrypt),
        .O(key_a[36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[37]_i_1 
       (.I0(key3[37]),
        .I1(key1[37]),
        .I2(decrypt),
        .O(key_a[37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[38]_i_1 
       (.I0(key3[38]),
        .I1(key1[38]),
        .I2(decrypt),
        .O(key_a[38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[39]_i_1 
       (.I0(key3[39]),
        .I1(key1[39]),
        .I2(decrypt),
        .O(key_a[39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[3]_i_1 
       (.I0(key3[3]),
        .I1(key1[3]),
        .I2(decrypt),
        .O(key_a[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[40]_i_1 
       (.I0(key3[40]),
        .I1(key1[40]),
        .I2(decrypt),
        .O(key_a[40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[41]_i_1 
       (.I0(key3[41]),
        .I1(key1[41]),
        .I2(decrypt),
        .O(key_a[41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[42]_i_1 
       (.I0(key3[42]),
        .I1(key1[42]),
        .I2(decrypt),
        .O(key_a[42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[43]_i_1 
       (.I0(key3[43]),
        .I1(key1[43]),
        .I2(decrypt),
        .O(key_a[43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[44]_i_1 
       (.I0(key3[44]),
        .I1(key1[44]),
        .I2(decrypt),
        .O(key_a[44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[45]_i_1 
       (.I0(key3[45]),
        .I1(key1[45]),
        .I2(decrypt),
        .O(key_a[45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[46]_i_1 
       (.I0(key3[46]),
        .I1(key1[46]),
        .I2(decrypt),
        .O(key_a[46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[47]_i_1 
       (.I0(key3[47]),
        .I1(key1[47]),
        .I2(decrypt),
        .O(key_a[47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[48]_i_1 
       (.I0(key3[48]),
        .I1(key1[48]),
        .I2(decrypt),
        .O(key_a[48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[49]_i_1 
       (.I0(key3[49]),
        .I1(key1[49]),
        .I2(decrypt),
        .O(key_a[49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[4]_i_1 
       (.I0(key3[4]),
        .I1(key1[4]),
        .I2(decrypt),
        .O(key_a[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[50]_i_1 
       (.I0(key3[50]),
        .I1(key1[50]),
        .I2(decrypt),
        .O(key_a[50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[51]_i_1 
       (.I0(key3[51]),
        .I1(key1[51]),
        .I2(decrypt),
        .O(key_a[51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[52]_i_1 
       (.I0(key3[52]),
        .I1(key1[52]),
        .I2(decrypt),
        .O(key_a[52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[53]_i_1 
       (.I0(key3[53]),
        .I1(key1[53]),
        .I2(decrypt),
        .O(key_a[53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[54]_i_1 
       (.I0(key3[54]),
        .I1(key1[54]),
        .I2(decrypt),
        .O(key_a[54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[55]_i_1 
       (.I0(key3[55]),
        .I1(key1[55]),
        .I2(decrypt),
        .O(key_a[55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[5]_i_1 
       (.I0(key3[5]),
        .I1(key1[5]),
        .I2(decrypt),
        .O(key_a[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[6]_i_1 
       (.I0(key3[6]),
        .I1(key1[6]),
        .I2(decrypt),
        .O(key_a[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[7]_i_1 
       (.I0(key3[7]),
        .I1(key1[7]),
        .I2(decrypt),
        .O(key_a[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[8]_i_1 
       (.I0(key3[8]),
        .I1(key1[8]),
        .I2(decrypt),
        .O(key_a[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \key_r[9]_i_1 
       (.I0(key3[9]),
        .I1(key1[9]),
        .I2(decrypt),
        .O(key_a[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [42]),
        .Q(\u0/L0 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [43]),
        .Q(\u0/L0 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [44]),
        .Q(\u0/L0 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [45]),
        .Q(\u0/L0 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [46]),
        .Q(\u0/L0 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [47]),
        .Q(\u0/L0 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [48]),
        .Q(\u0/L0 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [49]),
        .Q(\u0/L0 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [50]),
        .Q(\u0/L0 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [51]),
        .Q(\u0/L0 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [33]),
        .Q(\u0/L0 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [52]),
        .Q(\u0/L0 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [53]),
        .Q(\u0/L0 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [54]),
        .Q(\u0/L0 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [55]),
        .Q(\u0/L0 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [56]),
        .Q(\u0/L0 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [57]),
        .Q(\u0/L0 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [58]),
        .Q(\u0/L0 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [59]),
        .Q(\u0/L0 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [60]),
        .Q(\u0/L0 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [61]),
        .Q(\u0/L0 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [34]),
        .Q(\u0/L0 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [62]),
        .Q(\u0/L0 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [63]),
        .Q(\u0/L0 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [64]),
        .Q(\u0/L0 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [35]),
        .Q(\u0/L0 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [36]),
        .Q(\u0/L0 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [37]),
        .Q(\u0/L0 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [38]),
        .Q(\u0/L0 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [39]),
        .Q(\u0/L0 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [40]),
        .Q(\u0/L0 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L0_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/IP [41]),
        .Q(\u0/L0 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [10]),
        .Q(\u0/L10 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [11]),
        .Q(\u0/L10 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [12]),
        .Q(\u0/L10 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [13]),
        .Q(\u0/L10 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [14]),
        .Q(\u0/L10 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [15]),
        .Q(\u0/L10 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [16]),
        .Q(\u0/L10 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [17]),
        .Q(\u0/L10 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [18]),
        .Q(\u0/L10 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [19]),
        .Q(\u0/L10 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [1]),
        .Q(\u0/L10 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [20]),
        .Q(\u0/L10 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [21]),
        .Q(\u0/L10 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [22]),
        .Q(\u0/L10 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [23]),
        .Q(\u0/L10 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [24]),
        .Q(\u0/L10 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [25]),
        .Q(\u0/L10 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [26]),
        .Q(\u0/L10 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [27]),
        .Q(\u0/L10 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [28]),
        .Q(\u0/L10 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [29]),
        .Q(\u0/L10 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [2]),
        .Q(\u0/L10 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [30]),
        .Q(\u0/L10 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [31]),
        .Q(\u0/L10 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [32]),
        .Q(\u0/L10 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [3]),
        .Q(\u0/L10 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [4]),
        .Q(\u0/L10 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [5]),
        .Q(\u0/L10 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [6]),
        .Q(\u0/L10 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [7]),
        .Q(\u0/L10 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [8]),
        .Q(\u0/L10 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L10_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R9 [9]),
        .Q(\u0/L10 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_ ),
        .Q(\u0/L11 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[11] ),
        .Q(\u0/L11 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[12] ),
        .Q(\u0/L11 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[13] ),
        .Q(\u0/L11 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[14] ),
        .Q(\u0/L11 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[15] ),
        .Q(\u0/L11 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[16] ),
        .Q(\u0/L11 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[17] ),
        .Q(\u0/L11 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[18] ),
        .Q(\u0/L11 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[19] ),
        .Q(\u0/L11 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[1] ),
        .Q(\u0/L11 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[20] ),
        .Q(\u0/L11 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[21] ),
        .Q(\u0/L11 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[22] ),
        .Q(\u0/L11 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[23] ),
        .Q(\u0/L11 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[24] ),
        .Q(\u0/L11 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[25] ),
        .Q(\u0/L11 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[26] ),
        .Q(\u0/L11 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[27] ),
        .Q(\u0/L11 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[28] ),
        .Q(\u0/L11 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[29] ),
        .Q(\u0/L11 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[2] ),
        .Q(\u0/L11 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[30] ),
        .Q(\u0/L11 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[31] ),
        .Q(\u0/L11 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[32] ),
        .Q(\u0/L11 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[3] ),
        .Q(\u0/L11 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[4] ),
        .Q(\u0/L11 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[5] ),
        .Q(\u0/L11 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[6] ),
        .Q(\u0/L11 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[7] ),
        .Q(\u0/L11 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[8] ),
        .Q(\u0/L11 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L11_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10_reg_n_0_[9] ),
        .Q(\u0/L11 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [10]),
        .Q(\u0/L12 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [11]),
        .Q(\u0/L12 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [12]),
        .Q(\u0/L12 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [13]),
        .Q(\u0/L12 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [14]),
        .Q(\u0/L12 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [15]),
        .Q(\u0/L12 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [16]),
        .Q(\u0/L12 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [17]),
        .Q(\u0/L12 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [18]),
        .Q(\u0/L12 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [19]),
        .Q(\u0/L12 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [1]),
        .Q(\u0/L12 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [20]),
        .Q(\u0/L12 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [21]),
        .Q(\u0/L12 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [22]),
        .Q(\u0/L12 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [23]),
        .Q(\u0/L12 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [24]),
        .Q(\u0/L12 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [25]),
        .Q(\u0/L12 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [26]),
        .Q(\u0/L12 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [27]),
        .Q(\u0/L12 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [28]),
        .Q(\u0/L12 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [29]),
        .Q(\u0/L12 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [2]),
        .Q(\u0/L12 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [30]),
        .Q(\u0/L12 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [31]),
        .Q(\u0/L12 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [32]),
        .Q(\u0/L12 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [3]),
        .Q(\u0/L12 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [4]),
        .Q(\u0/L12 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [5]),
        .Q(\u0/L12 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [6]),
        .Q(\u0/L12 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [7]),
        .Q(\u0/L12 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [8]),
        .Q(\u0/L12 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L12_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R11 [9]),
        .Q(\u0/L12 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [10]),
        .Q(\u0/L13 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [11]),
        .Q(\u0/L13 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [12]),
        .Q(\u0/L13 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [13]),
        .Q(\u0/L13 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [14]),
        .Q(\u0/L13 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [15]),
        .Q(\u0/L13 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [16]),
        .Q(\u0/L13 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [17]),
        .Q(\u0/L13 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [18]),
        .Q(\u0/L13 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [19]),
        .Q(\u0/L13 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [1]),
        .Q(\u0/L13 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [20]),
        .Q(\u0/L13 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [21]),
        .Q(\u0/L13 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [22]),
        .Q(\u0/L13 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [23]),
        .Q(\u0/L13 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [24]),
        .Q(\u0/L13 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [25]),
        .Q(\u0/L13 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [26]),
        .Q(\u0/L13 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [27]),
        .Q(\u0/L13 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [28]),
        .Q(\u0/L13 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [29]),
        .Q(\u0/L13 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [2]),
        .Q(\u0/L13 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [30]),
        .Q(\u0/L13 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [31]),
        .Q(\u0/L13 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [32]),
        .Q(\u0/L13 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [3]),
        .Q(\u0/L13 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [4]),
        .Q(\u0/L13 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [5]),
        .Q(\u0/L13 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [6]),
        .Q(\u0/L13 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [7]),
        .Q(\u0/L13 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [8]),
        .Q(\u0/L13 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L13_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R12 [9]),
        .Q(\u0/L13 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [10]),
        .Q(\u0/L14 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [11]),
        .Q(\u0/L14 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [12]),
        .Q(\u0/L14 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [13]),
        .Q(\u0/L14 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [14]),
        .Q(\u0/L14 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [15]),
        .Q(\u0/L14 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [16]),
        .Q(\u0/L14 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [17]),
        .Q(\u0/L14 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [18]),
        .Q(\u0/L14 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [19]),
        .Q(\u0/L14 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [1]),
        .Q(\u0/L14 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [20]),
        .Q(\u0/L14 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [21]),
        .Q(\u0/L14 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [22]),
        .Q(\u0/L14 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [23]),
        .Q(\u0/L14 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [24]),
        .Q(\u0/L14 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [25]),
        .Q(\u0/L14 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [26]),
        .Q(\u0/L14 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [27]),
        .Q(\u0/L14 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [28]),
        .Q(\u0/L14 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [29]),
        .Q(\u0/L14 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [2]),
        .Q(\u0/L14 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [30]),
        .Q(\u0/L14 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [31]),
        .Q(\u0/L14 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [32]),
        .Q(\u0/L14 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [3]),
        .Q(\u0/L14 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [4]),
        .Q(\u0/L14 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [5]),
        .Q(\u0/L14 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [6]),
        .Q(\u0/L14 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [7]),
        .Q(\u0/L14 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [8]),
        .Q(\u0/L14 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L14_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R13 [9]),
        .Q(\u0/L14 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [10]),
        .Q(\u0/L1 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [11]),
        .Q(\u0/L1 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [12]),
        .Q(\u0/L1 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [13]),
        .Q(\u0/L1 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [14]),
        .Q(\u0/L1 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [15]),
        .Q(\u0/L1 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [16]),
        .Q(\u0/L1 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [17]),
        .Q(\u0/L1 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [18]),
        .Q(\u0/L1 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [19]),
        .Q(\u0/L1 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [1]),
        .Q(\u0/L1 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [20]),
        .Q(\u0/L1 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [21]),
        .Q(\u0/L1 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [22]),
        .Q(\u0/L1 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [23]),
        .Q(\u0/L1 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [24]),
        .Q(\u0/L1 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [25]),
        .Q(\u0/L1 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [26]),
        .Q(\u0/L1 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [27]),
        .Q(\u0/L1 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [28]),
        .Q(\u0/L1 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [29]),
        .Q(\u0/L1 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [2]),
        .Q(\u0/L1 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [30]),
        .Q(\u0/L1 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [31]),
        .Q(\u0/L1 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [32]),
        .Q(\u0/L1 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [3]),
        .Q(\u0/L1 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [4]),
        .Q(\u0/L1 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [5]),
        .Q(\u0/L1 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [6]),
        .Q(\u0/L1 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [7]),
        .Q(\u0/L1 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [8]),
        .Q(\u0/L1 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R0 [9]),
        .Q(\u0/L1 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [10]),
        .Q(\u0/L2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [11]),
        .Q(\u0/L2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [12]),
        .Q(\u0/L2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [13]),
        .Q(\u0/L2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [14]),
        .Q(\u0/L2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [15]),
        .Q(\u0/L2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [16]),
        .Q(\u0/L2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [17]),
        .Q(\u0/L2 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [18]),
        .Q(\u0/L2 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [19]),
        .Q(\u0/L2 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [1]),
        .Q(\u0/L2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [20]),
        .Q(\u0/L2 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [21]),
        .Q(\u0/L2 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [22]),
        .Q(\u0/L2 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [23]),
        .Q(\u0/L2 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [24]),
        .Q(\u0/L2 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [25]),
        .Q(\u0/L2 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [26]),
        .Q(\u0/L2 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [27]),
        .Q(\u0/L2 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [28]),
        .Q(\u0/L2 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [29]),
        .Q(\u0/L2 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [2]),
        .Q(\u0/L2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [30]),
        .Q(\u0/L2 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [31]),
        .Q(\u0/L2 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [32]),
        .Q(\u0/L2 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [3]),
        .Q(\u0/L2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [4]),
        .Q(\u0/L2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [5]),
        .Q(\u0/L2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [6]),
        .Q(\u0/L2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [7]),
        .Q(\u0/L2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [8]),
        .Q(\u0/L2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L2_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R1 [9]),
        .Q(\u0/L2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [10]),
        .Q(\u0/L3 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [11]),
        .Q(\u0/L3 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [12]),
        .Q(\u0/L3 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [13]),
        .Q(\u0/L3 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [14]),
        .Q(\u0/L3 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [15]),
        .Q(\u0/L3 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [16]),
        .Q(\u0/L3 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [17]),
        .Q(\u0/L3 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [18]),
        .Q(\u0/L3 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [19]),
        .Q(\u0/L3 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [1]),
        .Q(\u0/L3 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [20]),
        .Q(\u0/L3 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [21]),
        .Q(\u0/L3 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [22]),
        .Q(\u0/L3 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [23]),
        .Q(\u0/L3 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [24]),
        .Q(\u0/L3 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [25]),
        .Q(\u0/L3 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [26]),
        .Q(\u0/L3 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [27]),
        .Q(\u0/L3 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [28]),
        .Q(\u0/L3 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [29]),
        .Q(\u0/L3 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [2]),
        .Q(\u0/L3 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [30]),
        .Q(\u0/L3 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [31]),
        .Q(\u0/L3 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [32]),
        .Q(\u0/L3 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [3]),
        .Q(\u0/L3 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [4]),
        .Q(\u0/L3 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [5]),
        .Q(\u0/L3 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [6]),
        .Q(\u0/L3 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [7]),
        .Q(\u0/L3 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [8]),
        .Q(\u0/L3 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L3_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R2 [9]),
        .Q(\u0/L3 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [10]),
        .Q(\u0/L4 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [11]),
        .Q(\u0/L4 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [12]),
        .Q(\u0/L4 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [13]),
        .Q(\u0/L4 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [14]),
        .Q(\u0/L4 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [15]),
        .Q(\u0/L4 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [16]),
        .Q(\u0/L4 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [17]),
        .Q(\u0/L4 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [18]),
        .Q(\u0/L4 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [19]),
        .Q(\u0/L4 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [1]),
        .Q(\u0/L4 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [20]),
        .Q(\u0/L4 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [21]),
        .Q(\u0/L4 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [22]),
        .Q(\u0/L4 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [23]),
        .Q(\u0/L4 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [24]),
        .Q(\u0/L4 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [25]),
        .Q(\u0/L4 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [26]),
        .Q(\u0/L4 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [27]),
        .Q(\u0/L4 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [28]),
        .Q(\u0/L4 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [29]),
        .Q(\u0/L4 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [2]),
        .Q(\u0/L4 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [30]),
        .Q(\u0/L4 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [31]),
        .Q(\u0/L4 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [32]),
        .Q(\u0/L4 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [3]),
        .Q(\u0/L4 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [4]),
        .Q(\u0/L4 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [5]),
        .Q(\u0/L4 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [6]),
        .Q(\u0/L4 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [7]),
        .Q(\u0/L4 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [8]),
        .Q(\u0/L4 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L4_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R3 [9]),
        .Q(\u0/L4 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [10]),
        .Q(\u0/L5 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [11]),
        .Q(\u0/L5 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [12]),
        .Q(\u0/L5 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [13]),
        .Q(\u0/L5 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [14]),
        .Q(\u0/L5 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [15]),
        .Q(\u0/L5 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [16]),
        .Q(\u0/L5 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [17]),
        .Q(\u0/L5 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [18]),
        .Q(\u0/L5 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [19]),
        .Q(\u0/L5 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [1]),
        .Q(\u0/L5 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [20]),
        .Q(\u0/L5 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [21]),
        .Q(\u0/L5 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [22]),
        .Q(\u0/L5 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [23]),
        .Q(\u0/L5 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [24]),
        .Q(\u0/L5 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [25]),
        .Q(\u0/L5 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [26]),
        .Q(\u0/L5 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [27]),
        .Q(\u0/L5 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [28]),
        .Q(\u0/L5 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [29]),
        .Q(\u0/L5 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [2]),
        .Q(\u0/L5 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [30]),
        .Q(\u0/L5 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [31]),
        .Q(\u0/L5 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [32]),
        .Q(\u0/L5 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [3]),
        .Q(\u0/L5 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [4]),
        .Q(\u0/L5 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [5]),
        .Q(\u0/L5 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [6]),
        .Q(\u0/L5 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [7]),
        .Q(\u0/L5 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [8]),
        .Q(\u0/L5 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L5_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R4 [9]),
        .Q(\u0/L5 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [10]),
        .Q(\u0/L6 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [11]),
        .Q(\u0/L6 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [12]),
        .Q(\u0/L6 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [13]),
        .Q(\u0/L6 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [14]),
        .Q(\u0/L6 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [15]),
        .Q(\u0/L6 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [16]),
        .Q(\u0/L6 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [17]),
        .Q(\u0/L6 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [18]),
        .Q(\u0/L6 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [19]),
        .Q(\u0/L6 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [1]),
        .Q(\u0/L6 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [20]),
        .Q(\u0/L6 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [21]),
        .Q(\u0/L6 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [22]),
        .Q(\u0/L6 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [23]),
        .Q(\u0/L6 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [24]),
        .Q(\u0/L6 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [25]),
        .Q(\u0/L6 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [26]),
        .Q(\u0/L6 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [27]),
        .Q(\u0/L6 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [28]),
        .Q(\u0/L6 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [29]),
        .Q(\u0/L6 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [2]),
        .Q(\u0/L6 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [30]),
        .Q(\u0/L6 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [31]),
        .Q(\u0/L6 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [32]),
        .Q(\u0/L6 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [3]),
        .Q(\u0/L6 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [4]),
        .Q(\u0/L6 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [5]),
        .Q(\u0/L6 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [6]),
        .Q(\u0/L6 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [7]),
        .Q(\u0/L6 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [8]),
        .Q(\u0/L6 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L6_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R5 [9]),
        .Q(\u0/L6 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [10]),
        .Q(\u0/L7 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [11]),
        .Q(\u0/L7 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [12]),
        .Q(\u0/L7 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [13]),
        .Q(\u0/L7 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [14]),
        .Q(\u0/L7 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [15]),
        .Q(\u0/L7 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [16]),
        .Q(\u0/L7 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [17]),
        .Q(\u0/L7 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [18]),
        .Q(\u0/L7 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [19]),
        .Q(\u0/L7 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [1]),
        .Q(\u0/L7 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [20]),
        .Q(\u0/L7 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [21]),
        .Q(\u0/L7 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [22]),
        .Q(\u0/L7 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [23]),
        .Q(\u0/L7 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [24]),
        .Q(\u0/L7 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [25]),
        .Q(\u0/L7 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [26]),
        .Q(\u0/L7 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [27]),
        .Q(\u0/L7 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [28]),
        .Q(\u0/L7 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [29]),
        .Q(\u0/L7 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [2]),
        .Q(\u0/L7 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [30]),
        .Q(\u0/L7 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [31]),
        .Q(\u0/L7 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [32]),
        .Q(\u0/L7 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [3]),
        .Q(\u0/L7 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [4]),
        .Q(\u0/L7 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [5]),
        .Q(\u0/L7 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [6]),
        .Q(\u0/L7 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [7]),
        .Q(\u0/L7 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [8]),
        .Q(\u0/L7 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L7_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R6 [9]),
        .Q(\u0/L7 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [10]),
        .Q(\u0/L8 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [11]),
        .Q(\u0/L8 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [12]),
        .Q(\u0/L8 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [13]),
        .Q(\u0/L8 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [14]),
        .Q(\u0/L8 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [15]),
        .Q(\u0/L8 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [16]),
        .Q(\u0/L8 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [17]),
        .Q(\u0/L8 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [18]),
        .Q(\u0/L8 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [19]),
        .Q(\u0/L8 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [1]),
        .Q(\u0/L8 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [20]),
        .Q(\u0/L8 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [21]),
        .Q(\u0/L8 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [22]),
        .Q(\u0/L8 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [23]),
        .Q(\u0/L8 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [24]),
        .Q(\u0/L8 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [25]),
        .Q(\u0/L8 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [26]),
        .Q(\u0/L8 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [27]),
        .Q(\u0/L8 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [28]),
        .Q(\u0/L8 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [29]),
        .Q(\u0/L8 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [2]),
        .Q(\u0/L8 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [30]),
        .Q(\u0/L8 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [31]),
        .Q(\u0/L8 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [32]),
        .Q(\u0/L8 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [3]),
        .Q(\u0/L8 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [4]),
        .Q(\u0/L8 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [5]),
        .Q(\u0/L8 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [6]),
        .Q(\u0/L8 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [7]),
        .Q(\u0/L8 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [8]),
        .Q(\u0/L8 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L8_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R7 [9]),
        .Q(\u0/L8 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [10]),
        .Q(\u0/L9 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [11]),
        .Q(\u0/L9 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [12]),
        .Q(\u0/L9 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [13]),
        .Q(\u0/L9 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [14]),
        .Q(\u0/L9 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [15]),
        .Q(\u0/L9 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [16]),
        .Q(\u0/L9 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [17]),
        .Q(\u0/L9 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [18]),
        .Q(\u0/L9 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [19]),
        .Q(\u0/L9 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [1]),
        .Q(\u0/L9 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [20]),
        .Q(\u0/L9 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [21]),
        .Q(\u0/L9 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [22]),
        .Q(\u0/L9 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [23]),
        .Q(\u0/L9 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [24]),
        .Q(\u0/L9 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [25]),
        .Q(\u0/L9 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [26]),
        .Q(\u0/L9 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [27]),
        .Q(\u0/L9 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [28]),
        .Q(\u0/L9 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [29]),
        .Q(\u0/L9 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [2]),
        .Q(\u0/L9 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [30]),
        .Q(\u0/L9 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [31]),
        .Q(\u0/L9 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [32]),
        .Q(\u0/L9 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [3]),
        .Q(\u0/L9 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [4]),
        .Q(\u0/L9 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [5]),
        .Q(\u0/L9 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [6]),
        .Q(\u0/L9 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [7]),
        .Q(\u0/L9 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [8]),
        .Q(\u0/L9 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/L9_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R8 [9]),
        .Q(\u0/L9 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[10]_i_1 
       (.I0(\u0/IP [10]),
        .I1(\u0/out0 [10]),
        .O(\u0/R00 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[11]_i_1 
       (.I0(\u0/IP [11]),
        .I1(\u0/out0 [11]),
        .O(\u0/R00 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[12]_i_1 
       (.I0(\u0/IP [12]),
        .I1(\u0/out0 [12]),
        .O(\u0/R00 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[13]_i_1 
       (.I0(\u0/IP [13]),
        .I1(\u0/out0 [13]),
        .O(\u0/R00 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[14]_i_1 
       (.I0(\u0/IP [14]),
        .I1(\u0/out0 [14]),
        .O(\u0/R00 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[15]_i_1 
       (.I0(\u0/IP [15]),
        .I1(\u0/out0 [15]),
        .O(\u0/R00 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[16]_i_1 
       (.I0(\u0/IP [16]),
        .I1(\u0/out0 [16]),
        .O(\u0/R00 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[17]_i_1 
       (.I0(\u0/IP [17]),
        .I1(\u0/out0 [17]),
        .O(\u0/R00 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[18]_i_1 
       (.I0(\u0/IP [18]),
        .I1(\u0/out0 [18]),
        .O(\u0/R00 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[19]_i_1 
       (.I0(\u0/IP [19]),
        .I1(\u0/out0 [19]),
        .O(\u0/R00 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[1]_i_1 
       (.I0(\u0/IP [1]),
        .I1(\u0/out0 [1]),
        .O(\u0/R00 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[20]_i_1 
       (.I0(\u0/IP [20]),
        .I1(\u0/out0 [20]),
        .O(\u0/R00 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[21]_i_1 
       (.I0(\u0/IP [21]),
        .I1(\u0/out0 [21]),
        .O(\u0/R00 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[22]_i_1 
       (.I0(\u0/IP [22]),
        .I1(\u0/out0 [22]),
        .O(\u0/R00 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[23]_i_1 
       (.I0(\u0/IP [23]),
        .I1(\u0/out0 [23]),
        .O(\u0/R00 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[24]_i_1 
       (.I0(\u0/IP [24]),
        .I1(\u0/out0 [24]),
        .O(\u0/R00 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[25]_i_1 
       (.I0(\u0/IP [25]),
        .I1(\u0/out0 [25]),
        .O(\u0/R00 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[26]_i_1 
       (.I0(\u0/IP [26]),
        .I1(\u0/out0 [26]),
        .O(\u0/R00 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[27]_i_1 
       (.I0(\u0/IP [27]),
        .I1(\u0/out0 [27]),
        .O(\u0/R00 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[28]_i_1 
       (.I0(\u0/IP [28]),
        .I1(\u0/out0 [28]),
        .O(\u0/R00 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[29]_i_1 
       (.I0(\u0/IP [29]),
        .I1(\u0/out0 [29]),
        .O(\u0/R00 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[2]_i_1 
       (.I0(\u0/IP [2]),
        .I1(\u0/out0 [2]),
        .O(\u0/R00 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[30]_i_1 
       (.I0(\u0/IP [30]),
        .I1(\u0/out0 [30]),
        .O(\u0/R00 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[31]_i_1 
       (.I0(\u0/IP [31]),
        .I1(\u0/out0 [31]),
        .O(\u0/R00 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[32]_i_1 
       (.I0(\u0/IP [32]),
        .I1(\u0/out0 [32]),
        .O(\u0/R00 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[3]_i_1 
       (.I0(\u0/IP [3]),
        .I1(\u0/out0 [3]),
        .O(\u0/R00 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[4]_i_1 
       (.I0(\u0/IP [4]),
        .I1(\u0/out0 [4]),
        .O(\u0/R00 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[5]_i_1 
       (.I0(\u0/IP [5]),
        .I1(\u0/out0 [5]),
        .O(\u0/R00 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[6]_i_1 
       (.I0(\u0/IP [6]),
        .I1(\u0/out0 [6]),
        .O(\u0/R00 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[7]_i_1 
       (.I0(\u0/IP [7]),
        .I1(\u0/out0 [7]),
        .O(\u0/R00 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[8]_i_1 
       (.I0(\u0/IP [8]),
        .I1(\u0/out0 [8]),
        .O(\u0/R00 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R0[9]_i_1 
       (.I0(\u0/IP [9]),
        .I1(\u0/out0 [9]),
        .O(\u0/R00 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [22]),
        .Q(\u0/R0 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [21]),
        .Q(\u0/R0 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [20]),
        .Q(\u0/R0 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [19]),
        .Q(\u0/R0 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [18]),
        .Q(\u0/R0 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [17]),
        .Q(\u0/R0 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [16]),
        .Q(\u0/R0 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [15]),
        .Q(\u0/R0 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [14]),
        .Q(\u0/R0 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [13]),
        .Q(\u0/R0 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [31]),
        .Q(\u0/R0 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [12]),
        .Q(\u0/R0 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [11]),
        .Q(\u0/R0 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [10]),
        .Q(\u0/R0 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [9]),
        .Q(\u0/R0 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [8]),
        .Q(\u0/R0 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [7]),
        .Q(\u0/R0 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [6]),
        .Q(\u0/R0 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [5]),
        .Q(\u0/R0 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [4]),
        .Q(\u0/R0 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [3]),
        .Q(\u0/R0 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [30]),
        .Q(\u0/R0 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [2]),
        .Q(\u0/R0 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [1]),
        .Q(\u0/R0 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [0]),
        .Q(\u0/R0 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [29]),
        .Q(\u0/R0 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [28]),
        .Q(\u0/R0 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [27]),
        .Q(\u0/R0 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [26]),
        .Q(\u0/R0 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [25]),
        .Q(\u0/R0 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [24]),
        .Q(\u0/R0 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R0_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R00 [23]),
        .Q(\u0/R0 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[10]_i_1 
       (.I0(\u0/L9 [10]),
        .I1(\u0/out10 [10]),
        .O(\u0/R100 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[11]_i_1 
       (.I0(\u0/L9 [11]),
        .I1(\u0/out10 [11]),
        .O(\u0/R100 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[12]_i_1 
       (.I0(\u0/L9 [12]),
        .I1(\u0/out10 [12]),
        .O(\u0/R100 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[13]_i_1 
       (.I0(\u0/L9 [13]),
        .I1(\u0/out10 [13]),
        .O(\u0/R100 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[14]_i_1 
       (.I0(\u0/L9 [14]),
        .I1(\u0/out10 [14]),
        .O(\u0/R100 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[15]_i_1 
       (.I0(\u0/L9 [15]),
        .I1(\u0/out10 [15]),
        .O(\u0/R100 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[16]_i_1 
       (.I0(\u0/L9 [16]),
        .I1(\u0/out10 [16]),
        .O(\u0/R100 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[17]_i_1 
       (.I0(\u0/L9 [17]),
        .I1(\u0/out10 [17]),
        .O(\u0/R100 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[18]_i_1 
       (.I0(\u0/L9 [18]),
        .I1(\u0/out10 [18]),
        .O(\u0/R100 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[19]_i_1 
       (.I0(\u0/L9 [19]),
        .I1(\u0/out10 [19]),
        .O(\u0/R100 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[1]_i_1 
       (.I0(\u0/L9 [1]),
        .I1(\u0/out10 [1]),
        .O(\u0/R100 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[20]_i_1 
       (.I0(\u0/L9 [20]),
        .I1(\u0/out10 [20]),
        .O(\u0/R100 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[21]_i_1 
       (.I0(\u0/L9 [21]),
        .I1(\u0/out10 [21]),
        .O(\u0/R100 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[22]_i_1 
       (.I0(\u0/L9 [22]),
        .I1(\u0/out10 [22]),
        .O(\u0/R100 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[23]_i_1 
       (.I0(\u0/L9 [23]),
        .I1(\u0/out10 [23]),
        .O(\u0/R100 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[24]_i_1 
       (.I0(\u0/L9 [24]),
        .I1(\u0/out10 [24]),
        .O(\u0/R100 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[25]_i_1 
       (.I0(\u0/L9 [25]),
        .I1(\u0/out10 [25]),
        .O(\u0/R100 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[26]_i_1 
       (.I0(\u0/L9 [26]),
        .I1(\u0/out10 [26]),
        .O(\u0/R100 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[27]_i_1 
       (.I0(\u0/L9 [27]),
        .I1(\u0/out10 [27]),
        .O(\u0/R100 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[28]_i_1 
       (.I0(\u0/L9 [28]),
        .I1(\u0/out10 [28]),
        .O(\u0/R100 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[29]_i_1 
       (.I0(\u0/L9 [29]),
        .I1(\u0/out10 [29]),
        .O(\u0/R100 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[2]_i_1 
       (.I0(\u0/L9 [2]),
        .I1(\u0/out10 [2]),
        .O(\u0/R100 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[30]_i_1 
       (.I0(\u0/L9 [30]),
        .I1(\u0/out10 [30]),
        .O(\u0/R100 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[31]_i_1 
       (.I0(\u0/L9 [31]),
        .I1(\u0/out10 [31]),
        .O(\u0/R100 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[32]_i_1 
       (.I0(\u0/L9 [32]),
        .I1(\u0/out10 [32]),
        .O(\u0/R100 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[3]_i_1 
       (.I0(\u0/L9 [3]),
        .I1(\u0/out10 [3]),
        .O(\u0/R100 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[4]_i_1 
       (.I0(\u0/L9 [4]),
        .I1(\u0/out10 [4]),
        .O(\u0/R100 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[5]_i_1 
       (.I0(\u0/L9 [5]),
        .I1(\u0/out10 [5]),
        .O(\u0/R100 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[6]_i_1 
       (.I0(\u0/L9 [6]),
        .I1(\u0/out10 [6]),
        .O(\u0/R100 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[7]_i_1 
       (.I0(\u0/L9 [7]),
        .I1(\u0/out10 [7]),
        .O(\u0/R100 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[8]_i_1 
       (.I0(\u0/L9 [8]),
        .I1(\u0/out10 [8]),
        .O(\u0/R100 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R10[9]_i_1 
       (.I0(\u0/L9 [9]),
        .I1(\u0/out10 [9]),
        .O(\u0/R100 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [22]),
        .Q(\u0/R10_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [21]),
        .Q(\u0/R10_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [20]),
        .Q(\u0/R10_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [19]),
        .Q(\u0/R10_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [18]),
        .Q(\u0/R10_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [17]),
        .Q(\u0/R10_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [16]),
        .Q(\u0/R10_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [15]),
        .Q(\u0/R10_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [14]),
        .Q(\u0/R10_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [13]),
        .Q(\u0/R10_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [31]),
        .Q(\u0/R10_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [12]),
        .Q(\u0/R10_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [11]),
        .Q(\u0/R10_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [10]),
        .Q(\u0/R10_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [9]),
        .Q(\u0/R10_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [8]),
        .Q(\u0/R10_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [7]),
        .Q(\u0/R10_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [6]),
        .Q(\u0/R10_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [5]),
        .Q(\u0/R10_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [4]),
        .Q(\u0/R10_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [3]),
        .Q(\u0/R10_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [30]),
        .Q(\u0/R10_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [2]),
        .Q(\u0/R10_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [1]),
        .Q(\u0/R10_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [0]),
        .Q(\u0/R10_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [29]),
        .Q(\u0/R10_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [28]),
        .Q(\u0/R10_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [27]),
        .Q(\u0/R10_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [26]),
        .Q(\u0/R10_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [25]),
        .Q(\u0/R10_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [24]),
        .Q(\u0/R10_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R10_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R100 [23]),
        .Q(\u0/R10_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[10]_i_1 
       (.I0(\u0/L10 [10]),
        .I1(\u0/out11 [10]),
        .O(\u0/R110 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[11]_i_1 
       (.I0(\u0/L10 [11]),
        .I1(\u0/out11 [11]),
        .O(\u0/R110 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[12]_i_1 
       (.I0(\u0/L10 [12]),
        .I1(\u0/out11 [12]),
        .O(\u0/R110 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[13]_i_1 
       (.I0(\u0/L10 [13]),
        .I1(\u0/out11 [13]),
        .O(\u0/R110 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[14]_i_1 
       (.I0(\u0/L10 [14]),
        .I1(\u0/out11 [14]),
        .O(\u0/R110 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[15]_i_1 
       (.I0(\u0/L10 [15]),
        .I1(\u0/out11 [15]),
        .O(\u0/R110 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[16]_i_1 
       (.I0(\u0/L10 [16]),
        .I1(\u0/out11 [16]),
        .O(\u0/R110 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[17]_i_1 
       (.I0(\u0/L10 [17]),
        .I1(\u0/out11 [17]),
        .O(\u0/R110 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[18]_i_1 
       (.I0(\u0/L10 [18]),
        .I1(\u0/out11 [18]),
        .O(\u0/R110 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[19]_i_1 
       (.I0(\u0/L10 [19]),
        .I1(\u0/out11 [19]),
        .O(\u0/R110 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[1]_i_1 
       (.I0(\u0/L10 [1]),
        .I1(\u0/out11 [1]),
        .O(\u0/R110 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[20]_i_1 
       (.I0(\u0/L10 [20]),
        .I1(\u0/out11 [20]),
        .O(\u0/R110 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[21]_i_1 
       (.I0(\u0/L10 [21]),
        .I1(\u0/out11 [21]),
        .O(\u0/R110 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[22]_i_1 
       (.I0(\u0/L10 [22]),
        .I1(\u0/out11 [22]),
        .O(\u0/R110 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[23]_i_1 
       (.I0(\u0/L10 [23]),
        .I1(\u0/out11 [23]),
        .O(\u0/R110 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[24]_i_1 
       (.I0(\u0/L10 [24]),
        .I1(\u0/out11 [24]),
        .O(\u0/R110 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[25]_i_1 
       (.I0(\u0/L10 [25]),
        .I1(\u0/out11 [25]),
        .O(\u0/R110 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[26]_i_1 
       (.I0(\u0/L10 [26]),
        .I1(\u0/out11 [26]),
        .O(\u0/R110 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[27]_i_1 
       (.I0(\u0/L10 [27]),
        .I1(\u0/out11 [27]),
        .O(\u0/R110 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[28]_i_1 
       (.I0(\u0/L10 [28]),
        .I1(\u0/out11 [28]),
        .O(\u0/R110 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[29]_i_1 
       (.I0(\u0/L10 [29]),
        .I1(\u0/out11 [29]),
        .O(\u0/R110 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[2]_i_1 
       (.I0(\u0/L10 [2]),
        .I1(\u0/out11 [2]),
        .O(\u0/R110 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[30]_i_1 
       (.I0(\u0/L10 [30]),
        .I1(\u0/out11 [30]),
        .O(\u0/R110 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[31]_i_1 
       (.I0(\u0/L10 [31]),
        .I1(\u0/out11 [31]),
        .O(\u0/R110 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[32]_i_1 
       (.I0(\u0/L10 [32]),
        .I1(\u0/out11 [32]),
        .O(\u0/R110 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[3]_i_1 
       (.I0(\u0/L10 [3]),
        .I1(\u0/out11 [3]),
        .O(\u0/R110 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[4]_i_1 
       (.I0(\u0/L10 [4]),
        .I1(\u0/out11 [4]),
        .O(\u0/R110 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[5]_i_1 
       (.I0(\u0/L10 [5]),
        .I1(\u0/out11 [5]),
        .O(\u0/R110 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[6]_i_1 
       (.I0(\u0/L10 [6]),
        .I1(\u0/out11 [6]),
        .O(\u0/R110 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[7]_i_1 
       (.I0(\u0/L10 [7]),
        .I1(\u0/out11 [7]),
        .O(\u0/R110 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[8]_i_1 
       (.I0(\u0/L10 [8]),
        .I1(\u0/out11 [8]),
        .O(\u0/R110 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R11[9]_i_1 
       (.I0(\u0/L10 [9]),
        .I1(\u0/out11 [9]),
        .O(\u0/R110 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [22]),
        .Q(\u0/R11 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [21]),
        .Q(\u0/R11 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [20]),
        .Q(\u0/R11 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [19]),
        .Q(\u0/R11 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [18]),
        .Q(\u0/R11 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [17]),
        .Q(\u0/R11 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [16]),
        .Q(\u0/R11 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [15]),
        .Q(\u0/R11 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [14]),
        .Q(\u0/R11 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [13]),
        .Q(\u0/R11 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [31]),
        .Q(\u0/R11 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [12]),
        .Q(\u0/R11 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [11]),
        .Q(\u0/R11 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [10]),
        .Q(\u0/R11 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [9]),
        .Q(\u0/R11 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [8]),
        .Q(\u0/R11 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [7]),
        .Q(\u0/R11 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [6]),
        .Q(\u0/R11 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [5]),
        .Q(\u0/R11 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [4]),
        .Q(\u0/R11 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [3]),
        .Q(\u0/R11 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [30]),
        .Q(\u0/R11 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [2]),
        .Q(\u0/R11 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [1]),
        .Q(\u0/R11 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [0]),
        .Q(\u0/R11 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [29]),
        .Q(\u0/R11 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [28]),
        .Q(\u0/R11 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [27]),
        .Q(\u0/R11 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [26]),
        .Q(\u0/R11 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [25]),
        .Q(\u0/R11 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [24]),
        .Q(\u0/R11 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R11_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R110 [23]),
        .Q(\u0/R11 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[10]_i_1 
       (.I0(\u0/L11 [10]),
        .I1(\u0/out12 [10]),
        .O(\u0/R120 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[11]_i_1 
       (.I0(\u0/L11 [11]),
        .I1(\u0/out12 [11]),
        .O(\u0/R120 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[12]_i_1 
       (.I0(\u0/L11 [12]),
        .I1(\u0/out12 [12]),
        .O(\u0/R120 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[13]_i_1 
       (.I0(\u0/L11 [13]),
        .I1(\u0/out12 [13]),
        .O(\u0/R120 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[14]_i_1 
       (.I0(\u0/L11 [14]),
        .I1(\u0/out12 [14]),
        .O(\u0/R120 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[15]_i_1 
       (.I0(\u0/L11 [15]),
        .I1(\u0/out12 [15]),
        .O(\u0/R120 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[16]_i_1 
       (.I0(\u0/L11 [16]),
        .I1(\u0/out12 [16]),
        .O(\u0/R120 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[17]_i_1 
       (.I0(\u0/L11 [17]),
        .I1(\u0/out12 [17]),
        .O(\u0/R120 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[18]_i_1 
       (.I0(\u0/L11 [18]),
        .I1(\u0/out12 [18]),
        .O(\u0/R120 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[19]_i_1 
       (.I0(\u0/L11 [19]),
        .I1(\u0/out12 [19]),
        .O(\u0/R120 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[1]_i_1 
       (.I0(\u0/L11 [1]),
        .I1(\u0/out12 [1]),
        .O(\u0/R120 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[20]_i_1 
       (.I0(\u0/L11 [20]),
        .I1(\u0/out12 [20]),
        .O(\u0/R120 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[21]_i_1 
       (.I0(\u0/L11 [21]),
        .I1(\u0/out12 [21]),
        .O(\u0/R120 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[22]_i_1 
       (.I0(\u0/L11 [22]),
        .I1(\u0/out12 [22]),
        .O(\u0/R120 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[23]_i_1 
       (.I0(\u0/L11 [23]),
        .I1(\u0/out12 [23]),
        .O(\u0/R120 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[24]_i_1 
       (.I0(\u0/L11 [24]),
        .I1(\u0/out12 [24]),
        .O(\u0/R120 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[25]_i_1 
       (.I0(\u0/L11 [25]),
        .I1(\u0/out12 [25]),
        .O(\u0/R120 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[26]_i_1 
       (.I0(\u0/L11 [26]),
        .I1(\u0/out12 [26]),
        .O(\u0/R120 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[27]_i_1 
       (.I0(\u0/L11 [27]),
        .I1(\u0/out12 [27]),
        .O(\u0/R120 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[28]_i_1 
       (.I0(\u0/L11 [28]),
        .I1(\u0/out12 [28]),
        .O(\u0/R120 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[29]_i_1 
       (.I0(\u0/L11 [29]),
        .I1(\u0/out12 [29]),
        .O(\u0/R120 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[2]_i_1 
       (.I0(\u0/L11 [2]),
        .I1(\u0/out12 [2]),
        .O(\u0/R120 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[30]_i_1 
       (.I0(\u0/L11 [30]),
        .I1(\u0/out12 [30]),
        .O(\u0/R120 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[31]_i_1 
       (.I0(\u0/L11 [31]),
        .I1(\u0/out12 [31]),
        .O(\u0/R120 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[32]_i_1 
       (.I0(\u0/L11 [32]),
        .I1(\u0/out12 [32]),
        .O(\u0/R120 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[3]_i_1 
       (.I0(\u0/L11 [3]),
        .I1(\u0/out12 [3]),
        .O(\u0/R120 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[4]_i_1 
       (.I0(\u0/L11 [4]),
        .I1(\u0/out12 [4]),
        .O(\u0/R120 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[5]_i_1 
       (.I0(\u0/L11 [5]),
        .I1(\u0/out12 [5]),
        .O(\u0/R120 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[6]_i_1 
       (.I0(\u0/L11 [6]),
        .I1(\u0/out12 [6]),
        .O(\u0/R120 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[7]_i_1 
       (.I0(\u0/L11 [7]),
        .I1(\u0/out12 [7]),
        .O(\u0/R120 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[8]_i_1 
       (.I0(\u0/L11 [8]),
        .I1(\u0/out12 [8]),
        .O(\u0/R120 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R12[9]_i_1 
       (.I0(\u0/L11 [9]),
        .I1(\u0/out12 [9]),
        .O(\u0/R120 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [22]),
        .Q(\u0/R12 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [21]),
        .Q(\u0/R12 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [20]),
        .Q(\u0/R12 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [19]),
        .Q(\u0/R12 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [18]),
        .Q(\u0/R12 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [17]),
        .Q(\u0/R12 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [16]),
        .Q(\u0/R12 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [15]),
        .Q(\u0/R12 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [14]),
        .Q(\u0/R12 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [13]),
        .Q(\u0/R12 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [31]),
        .Q(\u0/R12 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [12]),
        .Q(\u0/R12 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [11]),
        .Q(\u0/R12 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [10]),
        .Q(\u0/R12 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [9]),
        .Q(\u0/R12 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [8]),
        .Q(\u0/R12 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [7]),
        .Q(\u0/R12 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [6]),
        .Q(\u0/R12 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [5]),
        .Q(\u0/R12 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [4]),
        .Q(\u0/R12 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [3]),
        .Q(\u0/R12 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [30]),
        .Q(\u0/R12 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [2]),
        .Q(\u0/R12 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [1]),
        .Q(\u0/R12 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [0]),
        .Q(\u0/R12 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [29]),
        .Q(\u0/R12 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [28]),
        .Q(\u0/R12 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [27]),
        .Q(\u0/R12 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [26]),
        .Q(\u0/R12 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [25]),
        .Q(\u0/R12 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [24]),
        .Q(\u0/R12 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R12_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R120 [23]),
        .Q(\u0/R12 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[10]_i_1 
       (.I0(\u0/L12 [10]),
        .I1(\u0/out13 [10]),
        .O(\u0/R130 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[11]_i_1 
       (.I0(\u0/L12 [11]),
        .I1(\u0/out13 [11]),
        .O(\u0/R130 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[12]_i_1 
       (.I0(\u0/L12 [12]),
        .I1(\u0/out13 [12]),
        .O(\u0/R130 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[13]_i_1 
       (.I0(\u0/L12 [13]),
        .I1(\u0/out13 [13]),
        .O(\u0/R130 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[14]_i_1 
       (.I0(\u0/L12 [14]),
        .I1(\u0/out13 [14]),
        .O(\u0/R130 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[15]_i_1 
       (.I0(\u0/L12 [15]),
        .I1(\u0/out13 [15]),
        .O(\u0/R130 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[16]_i_1 
       (.I0(\u0/L12 [16]),
        .I1(\u0/out13 [16]),
        .O(\u0/R130 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[17]_i_1 
       (.I0(\u0/L12 [17]),
        .I1(\u0/out13 [17]),
        .O(\u0/R130 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[18]_i_1 
       (.I0(\u0/L12 [18]),
        .I1(\u0/out13 [18]),
        .O(\u0/R130 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[19]_i_1 
       (.I0(\u0/L12 [19]),
        .I1(\u0/out13 [19]),
        .O(\u0/R130 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[1]_i_1 
       (.I0(\u0/L12 [1]),
        .I1(\u0/out13 [1]),
        .O(\u0/R130 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[20]_i_1 
       (.I0(\u0/L12 [20]),
        .I1(\u0/out13 [20]),
        .O(\u0/R130 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[21]_i_1 
       (.I0(\u0/L12 [21]),
        .I1(\u0/out13 [21]),
        .O(\u0/R130 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[22]_i_1 
       (.I0(\u0/L12 [22]),
        .I1(\u0/out13 [22]),
        .O(\u0/R130 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[23]_i_1 
       (.I0(\u0/L12 [23]),
        .I1(\u0/out13 [23]),
        .O(\u0/R130 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[24]_i_1 
       (.I0(\u0/L12 [24]),
        .I1(\u0/out13 [24]),
        .O(\u0/R130 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[25]_i_1 
       (.I0(\u0/L12 [25]),
        .I1(\u0/out13 [25]),
        .O(\u0/R130 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[26]_i_1 
       (.I0(\u0/L12 [26]),
        .I1(\u0/out13 [26]),
        .O(\u0/R130 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[27]_i_1 
       (.I0(\u0/L12 [27]),
        .I1(\u0/out13 [27]),
        .O(\u0/R130 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[28]_i_1 
       (.I0(\u0/L12 [28]),
        .I1(\u0/out13 [28]),
        .O(\u0/R130 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[29]_i_1 
       (.I0(\u0/L12 [29]),
        .I1(\u0/out13 [29]),
        .O(\u0/R130 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[2]_i_1 
       (.I0(\u0/L12 [2]),
        .I1(\u0/out13 [2]),
        .O(\u0/R130 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[30]_i_1 
       (.I0(\u0/L12 [30]),
        .I1(\u0/out13 [30]),
        .O(\u0/R130 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[31]_i_1 
       (.I0(\u0/L12 [31]),
        .I1(\u0/out13 [31]),
        .O(\u0/R130 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[32]_i_1 
       (.I0(\u0/L12 [32]),
        .I1(\u0/out13 [32]),
        .O(\u0/R130 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[3]_i_1 
       (.I0(\u0/L12 [3]),
        .I1(\u0/out13 [3]),
        .O(\u0/R130 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[4]_i_1 
       (.I0(\u0/L12 [4]),
        .I1(\u0/out13 [4]),
        .O(\u0/R130 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[5]_i_1 
       (.I0(\u0/L12 [5]),
        .I1(\u0/out13 [5]),
        .O(\u0/R130 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[6]_i_1 
       (.I0(\u0/L12 [6]),
        .I1(\u0/out13 [6]),
        .O(\u0/R130 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[7]_i_1 
       (.I0(\u0/L12 [7]),
        .I1(\u0/out13 [7]),
        .O(\u0/R130 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[8]_i_1 
       (.I0(\u0/L12 [8]),
        .I1(\u0/out13 [8]),
        .O(\u0/R130 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R13[9]_i_1 
       (.I0(\u0/L12 [9]),
        .I1(\u0/out13 [9]),
        .O(\u0/R130 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [22]),
        .Q(\u0/R13 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [21]),
        .Q(\u0/R13 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [20]),
        .Q(\u0/R13 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [19]),
        .Q(\u0/R13 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [18]),
        .Q(\u0/R13 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [17]),
        .Q(\u0/R13 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [16]),
        .Q(\u0/R13 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [15]),
        .Q(\u0/R13 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [14]),
        .Q(\u0/R13 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [13]),
        .Q(\u0/R13 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [31]),
        .Q(\u0/R13 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [12]),
        .Q(\u0/R13 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [11]),
        .Q(\u0/R13 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [10]),
        .Q(\u0/R13 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [9]),
        .Q(\u0/R13 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [8]),
        .Q(\u0/R13 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [7]),
        .Q(\u0/R13 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [6]),
        .Q(\u0/R13 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [5]),
        .Q(\u0/R13 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [4]),
        .Q(\u0/R13 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [3]),
        .Q(\u0/R13 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [30]),
        .Q(\u0/R13 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [2]),
        .Q(\u0/R13 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [1]),
        .Q(\u0/R13 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [0]),
        .Q(\u0/R13 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [29]),
        .Q(\u0/R13 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [28]),
        .Q(\u0/R13 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [27]),
        .Q(\u0/R13 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [26]),
        .Q(\u0/R13 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [25]),
        .Q(\u0/R13 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [24]),
        .Q(\u0/R13 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R13_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R130 [23]),
        .Q(\u0/R13 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[10]_i_1 
       (.I0(\u0/L13 [10]),
        .I1(\u0/out14 [10]),
        .O(\u0/R140 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[11]_i_1 
       (.I0(\u0/L13 [11]),
        .I1(\u0/out14 [11]),
        .O(\u0/R140 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[12]_i_1 
       (.I0(\u0/L13 [12]),
        .I1(\u0/out14 [12]),
        .O(\u0/R140 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[13]_i_1 
       (.I0(\u0/L13 [13]),
        .I1(\u0/out14 [13]),
        .O(\u0/R140 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[14]_i_1 
       (.I0(\u0/L13 [14]),
        .I1(\u0/out14 [14]),
        .O(\u0/R140 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[15]_i_1 
       (.I0(\u0/L13 [15]),
        .I1(\u0/out14 [15]),
        .O(\u0/R140 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[16]_i_1 
       (.I0(\u0/L13 [16]),
        .I1(\u0/out14 [16]),
        .O(\u0/R140 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[17]_i_1 
       (.I0(\u0/L13 [17]),
        .I1(\u0/out14 [17]),
        .O(\u0/R140 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[18]_i_1 
       (.I0(\u0/L13 [18]),
        .I1(\u0/out14 [18]),
        .O(\u0/R140 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[19]_i_1 
       (.I0(\u0/L13 [19]),
        .I1(\u0/out14 [19]),
        .O(\u0/R140 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[1]_i_1 
       (.I0(\u0/L13 [1]),
        .I1(\u0/out14 [1]),
        .O(\u0/R140 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[20]_i_1 
       (.I0(\u0/L13 [20]),
        .I1(\u0/out14 [20]),
        .O(\u0/R140 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[21]_i_1 
       (.I0(\u0/L13 [21]),
        .I1(\u0/out14 [21]),
        .O(\u0/R140 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[22]_i_1 
       (.I0(\u0/L13 [22]),
        .I1(\u0/out14 [22]),
        .O(\u0/R140 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[23]_i_1 
       (.I0(\u0/L13 [23]),
        .I1(\u0/out14 [23]),
        .O(\u0/R140 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[24]_i_1 
       (.I0(\u0/L13 [24]),
        .I1(\u0/out14 [24]),
        .O(\u0/R140 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[25]_i_1 
       (.I0(\u0/L13 [25]),
        .I1(\u0/out14 [25]),
        .O(\u0/R140 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[26]_i_1 
       (.I0(\u0/L13 [26]),
        .I1(\u0/out14 [26]),
        .O(\u0/R140 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[27]_i_1 
       (.I0(\u0/L13 [27]),
        .I1(\u0/out14 [27]),
        .O(\u0/R140 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[28]_i_1 
       (.I0(\u0/L13 [28]),
        .I1(\u0/out14 [28]),
        .O(\u0/R140 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[29]_i_1 
       (.I0(\u0/L13 [29]),
        .I1(\u0/out14 [29]),
        .O(\u0/R140 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[2]_i_1 
       (.I0(\u0/L13 [2]),
        .I1(\u0/out14 [2]),
        .O(\u0/R140 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[30]_i_1 
       (.I0(\u0/L13 [30]),
        .I1(\u0/out14 [30]),
        .O(\u0/R140 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[31]_i_1 
       (.I0(\u0/L13 [31]),
        .I1(\u0/out14 [31]),
        .O(\u0/R140 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[32]_i_1 
       (.I0(\u0/L13 [32]),
        .I1(\u0/out14 [32]),
        .O(\u0/R140 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[3]_i_1 
       (.I0(\u0/L13 [3]),
        .I1(\u0/out14 [3]),
        .O(\u0/R140 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[4]_i_1 
       (.I0(\u0/L13 [4]),
        .I1(\u0/out14 [4]),
        .O(\u0/R140 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[5]_i_1 
       (.I0(\u0/L13 [5]),
        .I1(\u0/out14 [5]),
        .O(\u0/R140 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[6]_i_1 
       (.I0(\u0/L13 [6]),
        .I1(\u0/out14 [6]),
        .O(\u0/R140 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[7]_i_1 
       (.I0(\u0/L13 [7]),
        .I1(\u0/out14 [7]),
        .O(\u0/R140 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[8]_i_1 
       (.I0(\u0/L13 [8]),
        .I1(\u0/out14 [8]),
        .O(\u0/R140 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R14[9]_i_1 
       (.I0(\u0/L13 [9]),
        .I1(\u0/out14 [9]),
        .O(\u0/R140 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [22]),
        .Q(\u0/FP [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [21]),
        .Q(\u0/FP [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [20]),
        .Q(\u0/FP [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [19]),
        .Q(\u0/FP [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [18]),
        .Q(\u0/FP [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [17]),
        .Q(\u0/FP [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [16]),
        .Q(\u0/FP [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [15]),
        .Q(\u0/FP [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [14]),
        .Q(\u0/FP [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [13]),
        .Q(\u0/FP [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [31]),
        .Q(\u0/FP [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [12]),
        .Q(\u0/FP [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [11]),
        .Q(\u0/FP [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [10]),
        .Q(\u0/FP [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [9]),
        .Q(\u0/FP [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [8]),
        .Q(\u0/FP [56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [7]),
        .Q(\u0/FP [57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [6]),
        .Q(\u0/FP [58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [5]),
        .Q(\u0/FP [59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [4]),
        .Q(\u0/FP [60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [3]),
        .Q(\u0/FP [61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [30]),
        .Q(\u0/FP [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [2]),
        .Q(\u0/FP [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [1]),
        .Q(\u0/FP [63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [0]),
        .Q(\u0/FP [64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [29]),
        .Q(\u0/FP [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [28]),
        .Q(\u0/FP [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [27]),
        .Q(\u0/FP [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [26]),
        .Q(\u0/FP [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [25]),
        .Q(\u0/FP [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [24]),
        .Q(\u0/FP [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R14_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R140 [23]),
        .Q(\u0/FP [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[10]_i_1 
       (.I0(\u0/L0 [10]),
        .I1(\u0/out1 [10]),
        .O(\u0/R10 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[11]_i_1 
       (.I0(\u0/L0 [11]),
        .I1(\u0/out1 [11]),
        .O(\u0/R10 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[12]_i_1 
       (.I0(\u0/L0 [12]),
        .I1(\u0/out1 [12]),
        .O(\u0/R10 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[13]_i_1 
       (.I0(\u0/L0 [13]),
        .I1(\u0/out1 [13]),
        .O(\u0/R10 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[14]_i_1 
       (.I0(\u0/L0 [14]),
        .I1(\u0/out1 [14]),
        .O(\u0/R10 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[15]_i_1 
       (.I0(\u0/L0 [15]),
        .I1(\u0/out1 [15]),
        .O(\u0/R10 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[16]_i_1 
       (.I0(\u0/L0 [16]),
        .I1(\u0/out1 [16]),
        .O(\u0/R10 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[17]_i_1 
       (.I0(\u0/L0 [17]),
        .I1(\u0/out1 [17]),
        .O(\u0/R10 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[18]_i_1 
       (.I0(\u0/L0 [18]),
        .I1(\u0/out1 [18]),
        .O(\u0/R10 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[19]_i_1 
       (.I0(\u0/L0 [19]),
        .I1(\u0/out1 [19]),
        .O(\u0/R10 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[1]_i_1 
       (.I0(\u0/L0 [1]),
        .I1(\u0/out1 [1]),
        .O(\u0/R10 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[20]_i_1 
       (.I0(\u0/L0 [20]),
        .I1(\u0/out1 [20]),
        .O(\u0/R10 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[21]_i_1 
       (.I0(\u0/L0 [21]),
        .I1(\u0/out1 [21]),
        .O(\u0/R10 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[22]_i_1 
       (.I0(\u0/L0 [22]),
        .I1(\u0/out1 [22]),
        .O(\u0/R10 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[23]_i_1 
       (.I0(\u0/L0 [23]),
        .I1(\u0/out1 [23]),
        .O(\u0/R10 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[24]_i_1 
       (.I0(\u0/L0 [24]),
        .I1(\u0/out1 [24]),
        .O(\u0/R10 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[25]_i_1 
       (.I0(\u0/L0 [25]),
        .I1(\u0/out1 [25]),
        .O(\u0/R10 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[26]_i_1 
       (.I0(\u0/L0 [26]),
        .I1(\u0/out1 [26]),
        .O(\u0/R10 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[27]_i_1 
       (.I0(\u0/L0 [27]),
        .I1(\u0/out1 [27]),
        .O(\u0/R10 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[28]_i_1 
       (.I0(\u0/L0 [28]),
        .I1(\u0/out1 [28]),
        .O(\u0/R10 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[29]_i_1 
       (.I0(\u0/L0 [29]),
        .I1(\u0/out1 [29]),
        .O(\u0/R10 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[2]_i_1 
       (.I0(\u0/L0 [2]),
        .I1(\u0/out1 [2]),
        .O(\u0/R10 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[30]_i_1 
       (.I0(\u0/L0 [30]),
        .I1(\u0/out1 [30]),
        .O(\u0/R10 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[31]_i_1 
       (.I0(\u0/L0 [31]),
        .I1(\u0/out1 [31]),
        .O(\u0/R10 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[32]_i_1 
       (.I0(\u0/L0 [32]),
        .I1(\u0/out1 [32]),
        .O(\u0/R10 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[3]_i_1 
       (.I0(\u0/L0 [3]),
        .I1(\u0/out1 [3]),
        .O(\u0/R10 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[4]_i_1 
       (.I0(\u0/L0 [4]),
        .I1(\u0/out1 [4]),
        .O(\u0/R10 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[5]_i_1 
       (.I0(\u0/L0 [5]),
        .I1(\u0/out1 [5]),
        .O(\u0/R10 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[6]_i_1 
       (.I0(\u0/L0 [6]),
        .I1(\u0/out1 [6]),
        .O(\u0/R10 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[7]_i_1 
       (.I0(\u0/L0 [7]),
        .I1(\u0/out1 [7]),
        .O(\u0/R10 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[8]_i_1 
       (.I0(\u0/L0 [8]),
        .I1(\u0/out1 [8]),
        .O(\u0/R10 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R1[9]_i_1 
       (.I0(\u0/L0 [9]),
        .I1(\u0/out1 [9]),
        .O(\u0/R10 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [22]),
        .Q(\u0/R1 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [21]),
        .Q(\u0/R1 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [20]),
        .Q(\u0/R1 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [19]),
        .Q(\u0/R1 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [18]),
        .Q(\u0/R1 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [17]),
        .Q(\u0/R1 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [16]),
        .Q(\u0/R1 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [15]),
        .Q(\u0/R1 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [14]),
        .Q(\u0/R1 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [13]),
        .Q(\u0/R1 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [31]),
        .Q(\u0/R1 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [12]),
        .Q(\u0/R1 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [11]),
        .Q(\u0/R1 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [10]),
        .Q(\u0/R1 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [9]),
        .Q(\u0/R1 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [8]),
        .Q(\u0/R1 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [7]),
        .Q(\u0/R1 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [6]),
        .Q(\u0/R1 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [5]),
        .Q(\u0/R1 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [4]),
        .Q(\u0/R1 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [3]),
        .Q(\u0/R1 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [30]),
        .Q(\u0/R1 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [2]),
        .Q(\u0/R1 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [1]),
        .Q(\u0/R1 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [0]),
        .Q(\u0/R1 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [29]),
        .Q(\u0/R1 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [28]),
        .Q(\u0/R1 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [27]),
        .Q(\u0/R1 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [26]),
        .Q(\u0/R1 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [25]),
        .Q(\u0/R1 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [24]),
        .Q(\u0/R1 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R10 [23]),
        .Q(\u0/R1 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[10]_i_1 
       (.I0(\u0/L1 [10]),
        .I1(\u0/out2 [10]),
        .O(\u0/R20 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[11]_i_1 
       (.I0(\u0/L1 [11]),
        .I1(\u0/out2 [11]),
        .O(\u0/R20 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[12]_i_1 
       (.I0(\u0/L1 [12]),
        .I1(\u0/out2 [12]),
        .O(\u0/R20 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[13]_i_1 
       (.I0(\u0/L1 [13]),
        .I1(\u0/out2 [13]),
        .O(\u0/R20 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[14]_i_1 
       (.I0(\u0/L1 [14]),
        .I1(\u0/out2 [14]),
        .O(\u0/R20 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[15]_i_1 
       (.I0(\u0/L1 [15]),
        .I1(\u0/out2 [15]),
        .O(\u0/R20 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[16]_i_1 
       (.I0(\u0/L1 [16]),
        .I1(\u0/out2 [16]),
        .O(\u0/R20 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[17]_i_1 
       (.I0(\u0/L1 [17]),
        .I1(\u0/out2 [17]),
        .O(\u0/R20 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[18]_i_1 
       (.I0(\u0/L1 [18]),
        .I1(\u0/out2 [18]),
        .O(\u0/R20 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[19]_i_1 
       (.I0(\u0/L1 [19]),
        .I1(\u0/out2 [19]),
        .O(\u0/R20 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[1]_i_1 
       (.I0(\u0/L1 [1]),
        .I1(\u0/out2 [1]),
        .O(\u0/R20 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[20]_i_1 
       (.I0(\u0/L1 [20]),
        .I1(\u0/out2 [20]),
        .O(\u0/R20 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[21]_i_1 
       (.I0(\u0/L1 [21]),
        .I1(\u0/out2 [21]),
        .O(\u0/R20 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[22]_i_1 
       (.I0(\u0/L1 [22]),
        .I1(\u0/out2 [22]),
        .O(\u0/R20 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[23]_i_1 
       (.I0(\u0/L1 [23]),
        .I1(\u0/out2 [23]),
        .O(\u0/R20 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[24]_i_1 
       (.I0(\u0/L1 [24]),
        .I1(\u0/out2 [24]),
        .O(\u0/R20 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[25]_i_1 
       (.I0(\u0/L1 [25]),
        .I1(\u0/out2 [25]),
        .O(\u0/R20 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[26]_i_1 
       (.I0(\u0/L1 [26]),
        .I1(\u0/out2 [26]),
        .O(\u0/R20 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[27]_i_1 
       (.I0(\u0/L1 [27]),
        .I1(\u0/out2 [27]),
        .O(\u0/R20 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[28]_i_1 
       (.I0(\u0/L1 [28]),
        .I1(\u0/out2 [28]),
        .O(\u0/R20 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[29]_i_1 
       (.I0(\u0/L1 [29]),
        .I1(\u0/out2 [29]),
        .O(\u0/R20 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[2]_i_1 
       (.I0(\u0/L1 [2]),
        .I1(\u0/out2 [2]),
        .O(\u0/R20 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[30]_i_1 
       (.I0(\u0/L1 [30]),
        .I1(\u0/out2 [30]),
        .O(\u0/R20 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[31]_i_1 
       (.I0(\u0/L1 [31]),
        .I1(\u0/out2 [31]),
        .O(\u0/R20 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[32]_i_1 
       (.I0(\u0/L1 [32]),
        .I1(\u0/out2 [32]),
        .O(\u0/R20 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[3]_i_1 
       (.I0(\u0/L1 [3]),
        .I1(\u0/out2 [3]),
        .O(\u0/R20 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[4]_i_1 
       (.I0(\u0/L1 [4]),
        .I1(\u0/out2 [4]),
        .O(\u0/R20 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[5]_i_1 
       (.I0(\u0/L1 [5]),
        .I1(\u0/out2 [5]),
        .O(\u0/R20 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[6]_i_1 
       (.I0(\u0/L1 [6]),
        .I1(\u0/out2 [6]),
        .O(\u0/R20 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[7]_i_1 
       (.I0(\u0/L1 [7]),
        .I1(\u0/out2 [7]),
        .O(\u0/R20 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[8]_i_1 
       (.I0(\u0/L1 [8]),
        .I1(\u0/out2 [8]),
        .O(\u0/R20 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R2[9]_i_1 
       (.I0(\u0/L1 [9]),
        .I1(\u0/out2 [9]),
        .O(\u0/R20 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [22]),
        .Q(\u0/R2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [21]),
        .Q(\u0/R2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [20]),
        .Q(\u0/R2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [19]),
        .Q(\u0/R2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [18]),
        .Q(\u0/R2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [17]),
        .Q(\u0/R2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [16]),
        .Q(\u0/R2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [15]),
        .Q(\u0/R2 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [14]),
        .Q(\u0/R2 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [13]),
        .Q(\u0/R2 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [31]),
        .Q(\u0/R2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [12]),
        .Q(\u0/R2 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [11]),
        .Q(\u0/R2 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [10]),
        .Q(\u0/R2 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [9]),
        .Q(\u0/R2 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [8]),
        .Q(\u0/R2 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [7]),
        .Q(\u0/R2 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [6]),
        .Q(\u0/R2 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [5]),
        .Q(\u0/R2 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [4]),
        .Q(\u0/R2 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [3]),
        .Q(\u0/R2 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [30]),
        .Q(\u0/R2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [2]),
        .Q(\u0/R2 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [1]),
        .Q(\u0/R2 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [0]),
        .Q(\u0/R2 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [29]),
        .Q(\u0/R2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [28]),
        .Q(\u0/R2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [27]),
        .Q(\u0/R2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [26]),
        .Q(\u0/R2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [25]),
        .Q(\u0/R2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [24]),
        .Q(\u0/R2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R2_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R20 [23]),
        .Q(\u0/R2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[10]_i_1 
       (.I0(\u0/L2 [10]),
        .I1(\u0/out3 [10]),
        .O(\u0/R30 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[11]_i_1 
       (.I0(\u0/L2 [11]),
        .I1(\u0/out3 [11]),
        .O(\u0/R30 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[12]_i_1 
       (.I0(\u0/L2 [12]),
        .I1(\u0/out3 [12]),
        .O(\u0/R30 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[13]_i_1 
       (.I0(\u0/L2 [13]),
        .I1(\u0/out3 [13]),
        .O(\u0/R30 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[14]_i_1 
       (.I0(\u0/L2 [14]),
        .I1(\u0/out3 [14]),
        .O(\u0/R30 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[15]_i_1 
       (.I0(\u0/L2 [15]),
        .I1(\u0/out3 [15]),
        .O(\u0/R30 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[16]_i_1 
       (.I0(\u0/L2 [16]),
        .I1(\u0/out3 [16]),
        .O(\u0/R30 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[17]_i_1 
       (.I0(\u0/L2 [17]),
        .I1(\u0/out3 [17]),
        .O(\u0/R30 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[18]_i_1 
       (.I0(\u0/L2 [18]),
        .I1(\u0/out3 [18]),
        .O(\u0/R30 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[19]_i_1 
       (.I0(\u0/L2 [19]),
        .I1(\u0/out3 [19]),
        .O(\u0/R30 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[1]_i_1 
       (.I0(\u0/L2 [1]),
        .I1(\u0/out3 [1]),
        .O(\u0/R30 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[20]_i_1 
       (.I0(\u0/L2 [20]),
        .I1(\u0/out3 [20]),
        .O(\u0/R30 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[21]_i_1 
       (.I0(\u0/L2 [21]),
        .I1(\u0/out3 [21]),
        .O(\u0/R30 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[22]_i_1 
       (.I0(\u0/L2 [22]),
        .I1(\u0/out3 [22]),
        .O(\u0/R30 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[23]_i_1 
       (.I0(\u0/L2 [23]),
        .I1(\u0/out3 [23]),
        .O(\u0/R30 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[24]_i_1 
       (.I0(\u0/L2 [24]),
        .I1(\u0/out3 [24]),
        .O(\u0/R30 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[25]_i_1 
       (.I0(\u0/L2 [25]),
        .I1(\u0/out3 [25]),
        .O(\u0/R30 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[26]_i_1 
       (.I0(\u0/L2 [26]),
        .I1(\u0/out3 [26]),
        .O(\u0/R30 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[27]_i_1 
       (.I0(\u0/L2 [27]),
        .I1(\u0/out3 [27]),
        .O(\u0/R30 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[28]_i_1 
       (.I0(\u0/L2 [28]),
        .I1(\u0/out3 [28]),
        .O(\u0/R30 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[29]_i_1 
       (.I0(\u0/L2 [29]),
        .I1(\u0/out3 [29]),
        .O(\u0/R30 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[2]_i_1 
       (.I0(\u0/L2 [2]),
        .I1(\u0/out3 [2]),
        .O(\u0/R30 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[30]_i_1 
       (.I0(\u0/L2 [30]),
        .I1(\u0/out3 [30]),
        .O(\u0/R30 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[31]_i_1 
       (.I0(\u0/L2 [31]),
        .I1(\u0/out3 [31]),
        .O(\u0/R30 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[32]_i_1 
       (.I0(\u0/L2 [32]),
        .I1(\u0/out3 [32]),
        .O(\u0/R30 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[3]_i_1 
       (.I0(\u0/L2 [3]),
        .I1(\u0/out3 [3]),
        .O(\u0/R30 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[4]_i_1 
       (.I0(\u0/L2 [4]),
        .I1(\u0/out3 [4]),
        .O(\u0/R30 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[5]_i_1 
       (.I0(\u0/L2 [5]),
        .I1(\u0/out3 [5]),
        .O(\u0/R30 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[6]_i_1 
       (.I0(\u0/L2 [6]),
        .I1(\u0/out3 [6]),
        .O(\u0/R30 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[7]_i_1 
       (.I0(\u0/L2 [7]),
        .I1(\u0/out3 [7]),
        .O(\u0/R30 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[8]_i_1 
       (.I0(\u0/L2 [8]),
        .I1(\u0/out3 [8]),
        .O(\u0/R30 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R3[9]_i_1 
       (.I0(\u0/L2 [9]),
        .I1(\u0/out3 [9]),
        .O(\u0/R30 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [22]),
        .Q(\u0/R3 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [21]),
        .Q(\u0/R3 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [20]),
        .Q(\u0/R3 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [19]),
        .Q(\u0/R3 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [18]),
        .Q(\u0/R3 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [17]),
        .Q(\u0/R3 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [16]),
        .Q(\u0/R3 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [15]),
        .Q(\u0/R3 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [14]),
        .Q(\u0/R3 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [13]),
        .Q(\u0/R3 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [31]),
        .Q(\u0/R3 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [12]),
        .Q(\u0/R3 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [11]),
        .Q(\u0/R3 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [10]),
        .Q(\u0/R3 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [9]),
        .Q(\u0/R3 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [8]),
        .Q(\u0/R3 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [7]),
        .Q(\u0/R3 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [6]),
        .Q(\u0/R3 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [5]),
        .Q(\u0/R3 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [4]),
        .Q(\u0/R3 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [3]),
        .Q(\u0/R3 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [30]),
        .Q(\u0/R3 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [2]),
        .Q(\u0/R3 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [1]),
        .Q(\u0/R3 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [0]),
        .Q(\u0/R3 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [29]),
        .Q(\u0/R3 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [28]),
        .Q(\u0/R3 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [27]),
        .Q(\u0/R3 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [26]),
        .Q(\u0/R3 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [25]),
        .Q(\u0/R3 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [24]),
        .Q(\u0/R3 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R3_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R30 [23]),
        .Q(\u0/R3 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[10]_i_1 
       (.I0(\u0/L3 [10]),
        .I1(\u0/out4 [10]),
        .O(\u0/R40 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[11]_i_1 
       (.I0(\u0/L3 [11]),
        .I1(\u0/out4 [11]),
        .O(\u0/R40 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[12]_i_1 
       (.I0(\u0/L3 [12]),
        .I1(\u0/out4 [12]),
        .O(\u0/R40 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[13]_i_1 
       (.I0(\u0/L3 [13]),
        .I1(\u0/out4 [13]),
        .O(\u0/R40 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[14]_i_1 
       (.I0(\u0/L3 [14]),
        .I1(\u0/out4 [14]),
        .O(\u0/R40 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[15]_i_1 
       (.I0(\u0/L3 [15]),
        .I1(\u0/out4 [15]),
        .O(\u0/R40 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[16]_i_1 
       (.I0(\u0/L3 [16]),
        .I1(\u0/out4 [16]),
        .O(\u0/R40 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[17]_i_1 
       (.I0(\u0/L3 [17]),
        .I1(\u0/out4 [17]),
        .O(\u0/R40 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[18]_i_1 
       (.I0(\u0/L3 [18]),
        .I1(\u0/out4 [18]),
        .O(\u0/R40 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[19]_i_1 
       (.I0(\u0/L3 [19]),
        .I1(\u0/out4 [19]),
        .O(\u0/R40 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[1]_i_1 
       (.I0(\u0/L3 [1]),
        .I1(\u0/out4 [1]),
        .O(\u0/R40 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[20]_i_1 
       (.I0(\u0/L3 [20]),
        .I1(\u0/out4 [20]),
        .O(\u0/R40 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[21]_i_1 
       (.I0(\u0/L3 [21]),
        .I1(\u0/out4 [21]),
        .O(\u0/R40 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[22]_i_1 
       (.I0(\u0/L3 [22]),
        .I1(\u0/out4 [22]),
        .O(\u0/R40 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[23]_i_1 
       (.I0(\u0/L3 [23]),
        .I1(\u0/out4 [23]),
        .O(\u0/R40 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[24]_i_1 
       (.I0(\u0/L3 [24]),
        .I1(\u0/out4 [24]),
        .O(\u0/R40 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[25]_i_1 
       (.I0(\u0/L3 [25]),
        .I1(\u0/out4 [25]),
        .O(\u0/R40 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[26]_i_1 
       (.I0(\u0/L3 [26]),
        .I1(\u0/out4 [26]),
        .O(\u0/R40 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[27]_i_1 
       (.I0(\u0/L3 [27]),
        .I1(\u0/out4 [27]),
        .O(\u0/R40 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[28]_i_1 
       (.I0(\u0/L3 [28]),
        .I1(\u0/out4 [28]),
        .O(\u0/R40 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[29]_i_1 
       (.I0(\u0/L3 [29]),
        .I1(\u0/out4 [29]),
        .O(\u0/R40 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[2]_i_1 
       (.I0(\u0/L3 [2]),
        .I1(\u0/out4 [2]),
        .O(\u0/R40 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[30]_i_1 
       (.I0(\u0/L3 [30]),
        .I1(\u0/out4 [30]),
        .O(\u0/R40 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[31]_i_1 
       (.I0(\u0/L3 [31]),
        .I1(\u0/out4 [31]),
        .O(\u0/R40 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[32]_i_1 
       (.I0(\u0/L3 [32]),
        .I1(\u0/out4 [32]),
        .O(\u0/R40 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[3]_i_1 
       (.I0(\u0/L3 [3]),
        .I1(\u0/out4 [3]),
        .O(\u0/R40 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[4]_i_1 
       (.I0(\u0/L3 [4]),
        .I1(\u0/out4 [4]),
        .O(\u0/R40 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[5]_i_1 
       (.I0(\u0/L3 [5]),
        .I1(\u0/out4 [5]),
        .O(\u0/R40 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[6]_i_1 
       (.I0(\u0/L3 [6]),
        .I1(\u0/out4 [6]),
        .O(\u0/R40 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[7]_i_1 
       (.I0(\u0/L3 [7]),
        .I1(\u0/out4 [7]),
        .O(\u0/R40 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[8]_i_1 
       (.I0(\u0/L3 [8]),
        .I1(\u0/out4 [8]),
        .O(\u0/R40 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R4[9]_i_1 
       (.I0(\u0/L3 [9]),
        .I1(\u0/out4 [9]),
        .O(\u0/R40 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [22]),
        .Q(\u0/R4 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [21]),
        .Q(\u0/R4 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [20]),
        .Q(\u0/R4 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [19]),
        .Q(\u0/R4 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [18]),
        .Q(\u0/R4 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [17]),
        .Q(\u0/R4 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [16]),
        .Q(\u0/R4 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [15]),
        .Q(\u0/R4 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [14]),
        .Q(\u0/R4 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [13]),
        .Q(\u0/R4 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [31]),
        .Q(\u0/R4 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [12]),
        .Q(\u0/R4 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [11]),
        .Q(\u0/R4 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [10]),
        .Q(\u0/R4 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [9]),
        .Q(\u0/R4 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [8]),
        .Q(\u0/R4 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [7]),
        .Q(\u0/R4 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [6]),
        .Q(\u0/R4 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [5]),
        .Q(\u0/R4 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [4]),
        .Q(\u0/R4 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [3]),
        .Q(\u0/R4 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [30]),
        .Q(\u0/R4 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [2]),
        .Q(\u0/R4 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [1]),
        .Q(\u0/R4 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [0]),
        .Q(\u0/R4 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [29]),
        .Q(\u0/R4 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [28]),
        .Q(\u0/R4 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [27]),
        .Q(\u0/R4 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [26]),
        .Q(\u0/R4 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [25]),
        .Q(\u0/R4 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [24]),
        .Q(\u0/R4 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R4_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R40 [23]),
        .Q(\u0/R4 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[10]_i_1 
       (.I0(\u0/L4 [10]),
        .I1(\u0/out5 [10]),
        .O(\u0/R50 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[11]_i_1 
       (.I0(\u0/L4 [11]),
        .I1(\u0/out5 [11]),
        .O(\u0/R50 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[12]_i_1 
       (.I0(\u0/L4 [12]),
        .I1(\u0/out5 [12]),
        .O(\u0/R50 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[13]_i_1 
       (.I0(\u0/L4 [13]),
        .I1(\u0/out5 [13]),
        .O(\u0/R50 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[14]_i_1 
       (.I0(\u0/L4 [14]),
        .I1(\u0/out5 [14]),
        .O(\u0/R50 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[15]_i_1 
       (.I0(\u0/L4 [15]),
        .I1(\u0/out5 [15]),
        .O(\u0/R50 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[16]_i_1 
       (.I0(\u0/L4 [16]),
        .I1(\u0/out5 [16]),
        .O(\u0/R50 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[17]_i_1 
       (.I0(\u0/L4 [17]),
        .I1(\u0/out5 [17]),
        .O(\u0/R50 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[18]_i_1 
       (.I0(\u0/L4 [18]),
        .I1(\u0/out5 [18]),
        .O(\u0/R50 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[19]_i_1 
       (.I0(\u0/L4 [19]),
        .I1(\u0/out5 [19]),
        .O(\u0/R50 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[1]_i_1 
       (.I0(\u0/L4 [1]),
        .I1(\u0/out5 [1]),
        .O(\u0/R50 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[20]_i_1 
       (.I0(\u0/L4 [20]),
        .I1(\u0/out5 [20]),
        .O(\u0/R50 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[21]_i_1 
       (.I0(\u0/L4 [21]),
        .I1(\u0/out5 [21]),
        .O(\u0/R50 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[22]_i_1 
       (.I0(\u0/L4 [22]),
        .I1(\u0/out5 [22]),
        .O(\u0/R50 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[23]_i_1 
       (.I0(\u0/L4 [23]),
        .I1(\u0/out5 [23]),
        .O(\u0/R50 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[24]_i_1 
       (.I0(\u0/L4 [24]),
        .I1(\u0/out5 [24]),
        .O(\u0/R50 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[25]_i_1 
       (.I0(\u0/L4 [25]),
        .I1(\u0/out5 [25]),
        .O(\u0/R50 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[26]_i_1 
       (.I0(\u0/L4 [26]),
        .I1(\u0/out5 [26]),
        .O(\u0/R50 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[27]_i_1 
       (.I0(\u0/L4 [27]),
        .I1(\u0/out5 [27]),
        .O(\u0/R50 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[28]_i_1 
       (.I0(\u0/L4 [28]),
        .I1(\u0/out5 [28]),
        .O(\u0/R50 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[29]_i_1 
       (.I0(\u0/L4 [29]),
        .I1(\u0/out5 [29]),
        .O(\u0/R50 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[2]_i_1 
       (.I0(\u0/L4 [2]),
        .I1(\u0/out5 [2]),
        .O(\u0/R50 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[30]_i_1 
       (.I0(\u0/L4 [30]),
        .I1(\u0/out5 [30]),
        .O(\u0/R50 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[31]_i_1 
       (.I0(\u0/L4 [31]),
        .I1(\u0/out5 [31]),
        .O(\u0/R50 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[32]_i_1 
       (.I0(\u0/L4 [32]),
        .I1(\u0/out5 [32]),
        .O(\u0/R50 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[3]_i_1 
       (.I0(\u0/L4 [3]),
        .I1(\u0/out5 [3]),
        .O(\u0/R50 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[4]_i_1 
       (.I0(\u0/L4 [4]),
        .I1(\u0/out5 [4]),
        .O(\u0/R50 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[5]_i_1 
       (.I0(\u0/L4 [5]),
        .I1(\u0/out5 [5]),
        .O(\u0/R50 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[6]_i_1 
       (.I0(\u0/L4 [6]),
        .I1(\u0/out5 [6]),
        .O(\u0/R50 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[7]_i_1 
       (.I0(\u0/L4 [7]),
        .I1(\u0/out5 [7]),
        .O(\u0/R50 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[8]_i_1 
       (.I0(\u0/L4 [8]),
        .I1(\u0/out5 [8]),
        .O(\u0/R50 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R5[9]_i_1 
       (.I0(\u0/L4 [9]),
        .I1(\u0/out5 [9]),
        .O(\u0/R50 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [22]),
        .Q(\u0/R5 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [21]),
        .Q(\u0/R5 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [20]),
        .Q(\u0/R5 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [19]),
        .Q(\u0/R5 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [18]),
        .Q(\u0/R5 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [17]),
        .Q(\u0/R5 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [16]),
        .Q(\u0/R5 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [15]),
        .Q(\u0/R5 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [14]),
        .Q(\u0/R5 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [13]),
        .Q(\u0/R5 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [31]),
        .Q(\u0/R5 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [12]),
        .Q(\u0/R5 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [11]),
        .Q(\u0/R5 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [10]),
        .Q(\u0/R5 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [9]),
        .Q(\u0/R5 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [8]),
        .Q(\u0/R5 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [7]),
        .Q(\u0/R5 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [6]),
        .Q(\u0/R5 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [5]),
        .Q(\u0/R5 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [4]),
        .Q(\u0/R5 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [3]),
        .Q(\u0/R5 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [30]),
        .Q(\u0/R5 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [2]),
        .Q(\u0/R5 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [1]),
        .Q(\u0/R5 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [0]),
        .Q(\u0/R5 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [29]),
        .Q(\u0/R5 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [28]),
        .Q(\u0/R5 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [27]),
        .Q(\u0/R5 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [26]),
        .Q(\u0/R5 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [25]),
        .Q(\u0/R5 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [24]),
        .Q(\u0/R5 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R5_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R50 [23]),
        .Q(\u0/R5 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[10]_i_1 
       (.I0(\u0/L5 [10]),
        .I1(\u0/out6 [10]),
        .O(\u0/R60 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[11]_i_1 
       (.I0(\u0/L5 [11]),
        .I1(\u0/out6 [11]),
        .O(\u0/R60 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[12]_i_1 
       (.I0(\u0/L5 [12]),
        .I1(\u0/out6 [12]),
        .O(\u0/R60 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[13]_i_1 
       (.I0(\u0/L5 [13]),
        .I1(\u0/out6 [13]),
        .O(\u0/R60 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[14]_i_1 
       (.I0(\u0/L5 [14]),
        .I1(\u0/out6 [14]),
        .O(\u0/R60 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[15]_i_1 
       (.I0(\u0/L5 [15]),
        .I1(\u0/out6 [15]),
        .O(\u0/R60 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[16]_i_1 
       (.I0(\u0/L5 [16]),
        .I1(\u0/out6 [16]),
        .O(\u0/R60 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[17]_i_1 
       (.I0(\u0/L5 [17]),
        .I1(\u0/out6 [17]),
        .O(\u0/R60 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[18]_i_1 
       (.I0(\u0/L5 [18]),
        .I1(\u0/out6 [18]),
        .O(\u0/R60 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[19]_i_1 
       (.I0(\u0/L5 [19]),
        .I1(\u0/out6 [19]),
        .O(\u0/R60 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[1]_i_1 
       (.I0(\u0/L5 [1]),
        .I1(\u0/out6 [1]),
        .O(\u0/R60 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[20]_i_1 
       (.I0(\u0/L5 [20]),
        .I1(\u0/out6 [20]),
        .O(\u0/R60 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[21]_i_1 
       (.I0(\u0/L5 [21]),
        .I1(\u0/out6 [21]),
        .O(\u0/R60 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[22]_i_1 
       (.I0(\u0/L5 [22]),
        .I1(\u0/out6 [22]),
        .O(\u0/R60 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[23]_i_1 
       (.I0(\u0/L5 [23]),
        .I1(\u0/out6 [23]),
        .O(\u0/R60 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[24]_i_1 
       (.I0(\u0/L5 [24]),
        .I1(\u0/out6 [24]),
        .O(\u0/R60 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[25]_i_1 
       (.I0(\u0/L5 [25]),
        .I1(\u0/out6 [25]),
        .O(\u0/R60 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[26]_i_1 
       (.I0(\u0/L5 [26]),
        .I1(\u0/out6 [26]),
        .O(\u0/R60 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[27]_i_1 
       (.I0(\u0/L5 [27]),
        .I1(\u0/out6 [27]),
        .O(\u0/R60 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[28]_i_1 
       (.I0(\u0/L5 [28]),
        .I1(\u0/out6 [28]),
        .O(\u0/R60 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[29]_i_1 
       (.I0(\u0/L5 [29]),
        .I1(\u0/out6 [29]),
        .O(\u0/R60 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[2]_i_1 
       (.I0(\u0/L5 [2]),
        .I1(\u0/out6 [2]),
        .O(\u0/R60 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[30]_i_1 
       (.I0(\u0/L5 [30]),
        .I1(\u0/out6 [30]),
        .O(\u0/R60 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[31]_i_1 
       (.I0(\u0/L5 [31]),
        .I1(\u0/out6 [31]),
        .O(\u0/R60 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[32]_i_1 
       (.I0(\u0/L5 [32]),
        .I1(\u0/out6 [32]),
        .O(\u0/R60 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[3]_i_1 
       (.I0(\u0/L5 [3]),
        .I1(\u0/out6 [3]),
        .O(\u0/R60 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[4]_i_1 
       (.I0(\u0/L5 [4]),
        .I1(\u0/out6 [4]),
        .O(\u0/R60 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[5]_i_1 
       (.I0(\u0/L5 [5]),
        .I1(\u0/out6 [5]),
        .O(\u0/R60 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[6]_i_1 
       (.I0(\u0/L5 [6]),
        .I1(\u0/out6 [6]),
        .O(\u0/R60 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[7]_i_1 
       (.I0(\u0/L5 [7]),
        .I1(\u0/out6 [7]),
        .O(\u0/R60 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[8]_i_1 
       (.I0(\u0/L5 [8]),
        .I1(\u0/out6 [8]),
        .O(\u0/R60 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R6[9]_i_1 
       (.I0(\u0/L5 [9]),
        .I1(\u0/out6 [9]),
        .O(\u0/R60 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [22]),
        .Q(\u0/R6 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [21]),
        .Q(\u0/R6 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [20]),
        .Q(\u0/R6 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [19]),
        .Q(\u0/R6 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [18]),
        .Q(\u0/R6 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [17]),
        .Q(\u0/R6 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [16]),
        .Q(\u0/R6 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [15]),
        .Q(\u0/R6 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [14]),
        .Q(\u0/R6 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [13]),
        .Q(\u0/R6 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [31]),
        .Q(\u0/R6 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [12]),
        .Q(\u0/R6 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [11]),
        .Q(\u0/R6 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [10]),
        .Q(\u0/R6 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [9]),
        .Q(\u0/R6 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [8]),
        .Q(\u0/R6 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [7]),
        .Q(\u0/R6 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [6]),
        .Q(\u0/R6 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [5]),
        .Q(\u0/R6 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [4]),
        .Q(\u0/R6 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [3]),
        .Q(\u0/R6 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [30]),
        .Q(\u0/R6 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [2]),
        .Q(\u0/R6 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [1]),
        .Q(\u0/R6 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [0]),
        .Q(\u0/R6 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [29]),
        .Q(\u0/R6 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [28]),
        .Q(\u0/R6 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [27]),
        .Q(\u0/R6 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [26]),
        .Q(\u0/R6 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [25]),
        .Q(\u0/R6 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [24]),
        .Q(\u0/R6 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R6_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R60 [23]),
        .Q(\u0/R6 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[10]_i_1 
       (.I0(\u0/L6 [10]),
        .I1(\u0/out7 [10]),
        .O(\u0/R70 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[11]_i_1 
       (.I0(\u0/L6 [11]),
        .I1(\u0/out7 [11]),
        .O(\u0/R70 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[12]_i_1 
       (.I0(\u0/L6 [12]),
        .I1(\u0/out7 [12]),
        .O(\u0/R70 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[13]_i_1 
       (.I0(\u0/L6 [13]),
        .I1(\u0/out7 [13]),
        .O(\u0/R70 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[14]_i_1 
       (.I0(\u0/L6 [14]),
        .I1(\u0/out7 [14]),
        .O(\u0/R70 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[15]_i_1 
       (.I0(\u0/L6 [15]),
        .I1(\u0/out7 [15]),
        .O(\u0/R70 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[16]_i_1 
       (.I0(\u0/L6 [16]),
        .I1(\u0/out7 [16]),
        .O(\u0/R70 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[17]_i_1 
       (.I0(\u0/L6 [17]),
        .I1(\u0/out7 [17]),
        .O(\u0/R70 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[18]_i_1 
       (.I0(\u0/L6 [18]),
        .I1(\u0/out7 [18]),
        .O(\u0/R70 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[19]_i_1 
       (.I0(\u0/L6 [19]),
        .I1(\u0/out7 [19]),
        .O(\u0/R70 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[1]_i_1 
       (.I0(\u0/L6 [1]),
        .I1(\u0/out7 [1]),
        .O(\u0/R70 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[20]_i_1 
       (.I0(\u0/L6 [20]),
        .I1(\u0/out7 [20]),
        .O(\u0/R70 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[21]_i_1 
       (.I0(\u0/L6 [21]),
        .I1(\u0/out7 [21]),
        .O(\u0/R70 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[22]_i_1 
       (.I0(\u0/L6 [22]),
        .I1(\u0/out7 [22]),
        .O(\u0/R70 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[23]_i_1 
       (.I0(\u0/L6 [23]),
        .I1(\u0/out7 [23]),
        .O(\u0/R70 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[24]_i_1 
       (.I0(\u0/L6 [24]),
        .I1(\u0/out7 [24]),
        .O(\u0/R70 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[25]_i_1 
       (.I0(\u0/L6 [25]),
        .I1(\u0/out7 [25]),
        .O(\u0/R70 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[26]_i_1 
       (.I0(\u0/L6 [26]),
        .I1(\u0/out7 [26]),
        .O(\u0/R70 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[27]_i_1 
       (.I0(\u0/L6 [27]),
        .I1(\u0/out7 [27]),
        .O(\u0/R70 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[28]_i_1 
       (.I0(\u0/L6 [28]),
        .I1(\u0/out7 [28]),
        .O(\u0/R70 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[29]_i_1 
       (.I0(\u0/L6 [29]),
        .I1(\u0/out7 [29]),
        .O(\u0/R70 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[2]_i_1 
       (.I0(\u0/L6 [2]),
        .I1(\u0/out7 [2]),
        .O(\u0/R70 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[30]_i_1 
       (.I0(\u0/L6 [30]),
        .I1(\u0/out7 [30]),
        .O(\u0/R70 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[31]_i_1 
       (.I0(\u0/L6 [31]),
        .I1(\u0/out7 [31]),
        .O(\u0/R70 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[32]_i_1 
       (.I0(\u0/L6 [32]),
        .I1(\u0/out7 [32]),
        .O(\u0/R70 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[3]_i_1 
       (.I0(\u0/L6 [3]),
        .I1(\u0/out7 [3]),
        .O(\u0/R70 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[4]_i_1 
       (.I0(\u0/L6 [4]),
        .I1(\u0/out7 [4]),
        .O(\u0/R70 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[5]_i_1 
       (.I0(\u0/L6 [5]),
        .I1(\u0/out7 [5]),
        .O(\u0/R70 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[6]_i_1 
       (.I0(\u0/L6 [6]),
        .I1(\u0/out7 [6]),
        .O(\u0/R70 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[7]_i_1 
       (.I0(\u0/L6 [7]),
        .I1(\u0/out7 [7]),
        .O(\u0/R70 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[8]_i_1 
       (.I0(\u0/L6 [8]),
        .I1(\u0/out7 [8]),
        .O(\u0/R70 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R7[9]_i_1 
       (.I0(\u0/L6 [9]),
        .I1(\u0/out7 [9]),
        .O(\u0/R70 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [22]),
        .Q(\u0/R7 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [21]),
        .Q(\u0/R7 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [20]),
        .Q(\u0/R7 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [19]),
        .Q(\u0/R7 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [18]),
        .Q(\u0/R7 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [17]),
        .Q(\u0/R7 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [16]),
        .Q(\u0/R7 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [15]),
        .Q(\u0/R7 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [14]),
        .Q(\u0/R7 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [13]),
        .Q(\u0/R7 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [31]),
        .Q(\u0/R7 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [12]),
        .Q(\u0/R7 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [11]),
        .Q(\u0/R7 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [10]),
        .Q(\u0/R7 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [9]),
        .Q(\u0/R7 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [8]),
        .Q(\u0/R7 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [7]),
        .Q(\u0/R7 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [6]),
        .Q(\u0/R7 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [5]),
        .Q(\u0/R7 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [4]),
        .Q(\u0/R7 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [3]),
        .Q(\u0/R7 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [30]),
        .Q(\u0/R7 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [2]),
        .Q(\u0/R7 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [1]),
        .Q(\u0/R7 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [0]),
        .Q(\u0/R7 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [29]),
        .Q(\u0/R7 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [28]),
        .Q(\u0/R7 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [27]),
        .Q(\u0/R7 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [26]),
        .Q(\u0/R7 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [25]),
        .Q(\u0/R7 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [24]),
        .Q(\u0/R7 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R7_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R70 [23]),
        .Q(\u0/R7 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[10]_i_1 
       (.I0(\u0/L7 [10]),
        .I1(\u0/out8 [10]),
        .O(\u0/R80 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[11]_i_1 
       (.I0(\u0/L7 [11]),
        .I1(\u0/out8 [11]),
        .O(\u0/R80 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[12]_i_1 
       (.I0(\u0/L7 [12]),
        .I1(\u0/out8 [12]),
        .O(\u0/R80 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[13]_i_1 
       (.I0(\u0/L7 [13]),
        .I1(\u0/out8 [13]),
        .O(\u0/R80 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[14]_i_1 
       (.I0(\u0/L7 [14]),
        .I1(\u0/out8 [14]),
        .O(\u0/R80 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[15]_i_1 
       (.I0(\u0/L7 [15]),
        .I1(\u0/out8 [15]),
        .O(\u0/R80 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[16]_i_1 
       (.I0(\u0/L7 [16]),
        .I1(\u0/out8 [16]),
        .O(\u0/R80 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[17]_i_1 
       (.I0(\u0/L7 [17]),
        .I1(\u0/out8 [17]),
        .O(\u0/R80 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[18]_i_1 
       (.I0(\u0/L7 [18]),
        .I1(\u0/out8 [18]),
        .O(\u0/R80 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[19]_i_1 
       (.I0(\u0/L7 [19]),
        .I1(\u0/out8 [19]),
        .O(\u0/R80 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[1]_i_1 
       (.I0(\u0/L7 [1]),
        .I1(\u0/out8 [1]),
        .O(\u0/R80 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[20]_i_1 
       (.I0(\u0/L7 [20]),
        .I1(\u0/out8 [20]),
        .O(\u0/R80 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[21]_i_1 
       (.I0(\u0/L7 [21]),
        .I1(\u0/out8 [21]),
        .O(\u0/R80 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[22]_i_1 
       (.I0(\u0/L7 [22]),
        .I1(\u0/out8 [22]),
        .O(\u0/R80 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[23]_i_1 
       (.I0(\u0/L7 [23]),
        .I1(\u0/out8 [23]),
        .O(\u0/R80 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[24]_i_1 
       (.I0(\u0/L7 [24]),
        .I1(\u0/out8 [24]),
        .O(\u0/R80 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[25]_i_1 
       (.I0(\u0/L7 [25]),
        .I1(\u0/out8 [25]),
        .O(\u0/R80 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[26]_i_1 
       (.I0(\u0/L7 [26]),
        .I1(\u0/out8 [26]),
        .O(\u0/R80 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[27]_i_1 
       (.I0(\u0/L7 [27]),
        .I1(\u0/out8 [27]),
        .O(\u0/R80 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[28]_i_1 
       (.I0(\u0/L7 [28]),
        .I1(\u0/out8 [28]),
        .O(\u0/R80 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[29]_i_1 
       (.I0(\u0/L7 [29]),
        .I1(\u0/out8 [29]),
        .O(\u0/R80 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[2]_i_1 
       (.I0(\u0/L7 [2]),
        .I1(\u0/out8 [2]),
        .O(\u0/R80 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[30]_i_1 
       (.I0(\u0/L7 [30]),
        .I1(\u0/out8 [30]),
        .O(\u0/R80 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[31]_i_1 
       (.I0(\u0/L7 [31]),
        .I1(\u0/out8 [31]),
        .O(\u0/R80 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[32]_i_1 
       (.I0(\u0/L7 [32]),
        .I1(\u0/out8 [32]),
        .O(\u0/R80 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[3]_i_1 
       (.I0(\u0/L7 [3]),
        .I1(\u0/out8 [3]),
        .O(\u0/R80 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[4]_i_1 
       (.I0(\u0/L7 [4]),
        .I1(\u0/out8 [4]),
        .O(\u0/R80 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[5]_i_1 
       (.I0(\u0/L7 [5]),
        .I1(\u0/out8 [5]),
        .O(\u0/R80 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[6]_i_1 
       (.I0(\u0/L7 [6]),
        .I1(\u0/out8 [6]),
        .O(\u0/R80 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[7]_i_1 
       (.I0(\u0/L7 [7]),
        .I1(\u0/out8 [7]),
        .O(\u0/R80 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[8]_i_1 
       (.I0(\u0/L7 [8]),
        .I1(\u0/out8 [8]),
        .O(\u0/R80 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R8[9]_i_1 
       (.I0(\u0/L7 [9]),
        .I1(\u0/out8 [9]),
        .O(\u0/R80 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [22]),
        .Q(\u0/R8 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [21]),
        .Q(\u0/R8 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [20]),
        .Q(\u0/R8 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [19]),
        .Q(\u0/R8 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [18]),
        .Q(\u0/R8 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [17]),
        .Q(\u0/R8 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [16]),
        .Q(\u0/R8 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [15]),
        .Q(\u0/R8 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [14]),
        .Q(\u0/R8 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [13]),
        .Q(\u0/R8 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [31]),
        .Q(\u0/R8 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [12]),
        .Q(\u0/R8 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [11]),
        .Q(\u0/R8 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [10]),
        .Q(\u0/R8 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [9]),
        .Q(\u0/R8 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [8]),
        .Q(\u0/R8 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [7]),
        .Q(\u0/R8 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [6]),
        .Q(\u0/R8 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [5]),
        .Q(\u0/R8 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [4]),
        .Q(\u0/R8 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [3]),
        .Q(\u0/R8 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [30]),
        .Q(\u0/R8 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [2]),
        .Q(\u0/R8 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [1]),
        .Q(\u0/R8 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [0]),
        .Q(\u0/R8 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [29]),
        .Q(\u0/R8 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [28]),
        .Q(\u0/R8 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [27]),
        .Q(\u0/R8 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [26]),
        .Q(\u0/R8 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [25]),
        .Q(\u0/R8 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [24]),
        .Q(\u0/R8 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R8_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R80 [23]),
        .Q(\u0/R8 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[10]_i_1 
       (.I0(\u0/L8 [10]),
        .I1(\u0/out9 [10]),
        .O(\u0/R90 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[11]_i_1 
       (.I0(\u0/L8 [11]),
        .I1(\u0/out9 [11]),
        .O(\u0/R90 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[12]_i_1 
       (.I0(\u0/L8 [12]),
        .I1(\u0/out9 [12]),
        .O(\u0/R90 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[13]_i_1 
       (.I0(\u0/L8 [13]),
        .I1(\u0/out9 [13]),
        .O(\u0/R90 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[14]_i_1 
       (.I0(\u0/L8 [14]),
        .I1(\u0/out9 [14]),
        .O(\u0/R90 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[15]_i_1 
       (.I0(\u0/L8 [15]),
        .I1(\u0/out9 [15]),
        .O(\u0/R90 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[16]_i_1 
       (.I0(\u0/L8 [16]),
        .I1(\u0/out9 [16]),
        .O(\u0/R90 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[17]_i_1 
       (.I0(\u0/L8 [17]),
        .I1(\u0/out9 [17]),
        .O(\u0/R90 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[18]_i_1 
       (.I0(\u0/L8 [18]),
        .I1(\u0/out9 [18]),
        .O(\u0/R90 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[19]_i_1 
       (.I0(\u0/L8 [19]),
        .I1(\u0/out9 [19]),
        .O(\u0/R90 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[1]_i_1 
       (.I0(\u0/L8 [1]),
        .I1(\u0/out9 [1]),
        .O(\u0/R90 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[20]_i_1 
       (.I0(\u0/L8 [20]),
        .I1(\u0/out9 [20]),
        .O(\u0/R90 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[21]_i_1 
       (.I0(\u0/L8 [21]),
        .I1(\u0/out9 [21]),
        .O(\u0/R90 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[22]_i_1 
       (.I0(\u0/L8 [22]),
        .I1(\u0/out9 [22]),
        .O(\u0/R90 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[23]_i_1 
       (.I0(\u0/L8 [23]),
        .I1(\u0/out9 [23]),
        .O(\u0/R90 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[24]_i_1 
       (.I0(\u0/L8 [24]),
        .I1(\u0/out9 [24]),
        .O(\u0/R90 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[25]_i_1 
       (.I0(\u0/L8 [25]),
        .I1(\u0/out9 [25]),
        .O(\u0/R90 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[26]_i_1 
       (.I0(\u0/L8 [26]),
        .I1(\u0/out9 [26]),
        .O(\u0/R90 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[27]_i_1 
       (.I0(\u0/L8 [27]),
        .I1(\u0/out9 [27]),
        .O(\u0/R90 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[28]_i_1 
       (.I0(\u0/L8 [28]),
        .I1(\u0/out9 [28]),
        .O(\u0/R90 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[29]_i_1 
       (.I0(\u0/L8 [29]),
        .I1(\u0/out9 [29]),
        .O(\u0/R90 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[2]_i_1 
       (.I0(\u0/L8 [2]),
        .I1(\u0/out9 [2]),
        .O(\u0/R90 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[30]_i_1 
       (.I0(\u0/L8 [30]),
        .I1(\u0/out9 [30]),
        .O(\u0/R90 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[31]_i_1 
       (.I0(\u0/L8 [31]),
        .I1(\u0/out9 [31]),
        .O(\u0/R90 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[32]_i_1 
       (.I0(\u0/L8 [32]),
        .I1(\u0/out9 [32]),
        .O(\u0/R90 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[3]_i_1 
       (.I0(\u0/L8 [3]),
        .I1(\u0/out9 [3]),
        .O(\u0/R90 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[4]_i_1 
       (.I0(\u0/L8 [4]),
        .I1(\u0/out9 [4]),
        .O(\u0/R90 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[5]_i_1 
       (.I0(\u0/L8 [5]),
        .I1(\u0/out9 [5]),
        .O(\u0/R90 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[6]_i_1 
       (.I0(\u0/L8 [6]),
        .I1(\u0/out9 [6]),
        .O(\u0/R90 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[7]_i_1 
       (.I0(\u0/L8 [7]),
        .I1(\u0/out9 [7]),
        .O(\u0/R90 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[8]_i_1 
       (.I0(\u0/L8 [8]),
        .I1(\u0/out9 [8]),
        .O(\u0/R90 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/R9[9]_i_1 
       (.I0(\u0/L8 [9]),
        .I1(\u0/out9 [9]),
        .O(\u0/R90 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [22]),
        .Q(\u0/R9 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [21]),
        .Q(\u0/R9 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [20]),
        .Q(\u0/R9 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [19]),
        .Q(\u0/R9 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [18]),
        .Q(\u0/R9 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [17]),
        .Q(\u0/R9 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [16]),
        .Q(\u0/R9 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [15]),
        .Q(\u0/R9 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [14]),
        .Q(\u0/R9 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [13]),
        .Q(\u0/R9 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [31]),
        .Q(\u0/R9 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [12]),
        .Q(\u0/R9 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [11]),
        .Q(\u0/R9 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [10]),
        .Q(\u0/R9 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [9]),
        .Q(\u0/R9 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [8]),
        .Q(\u0/R9 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [7]),
        .Q(\u0/R9 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [6]),
        .Q(\u0/R9 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [5]),
        .Q(\u0/R9 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [4]),
        .Q(\u0/R9 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [3]),
        .Q(\u0/R9 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [30]),
        .Q(\u0/R9 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [2]),
        .Q(\u0/R9 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [1]),
        .Q(\u0/R9 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [0]),
        .Q(\u0/R9 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [29]),
        .Q(\u0/R9 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [28]),
        .Q(\u0/R9 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [27]),
        .Q(\u0/R9 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [26]),
        .Q(\u0/R9 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [25]),
        .Q(\u0/R9 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [24]),
        .Q(\u0/R9 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/R9_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/R90 [23]),
        .Q(\u0/R9 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[0]),
        .Q(\u0/IP [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[10]),
        .Q(\u0/IP [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[11]),
        .Q(\u0/IP [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[12]),
        .Q(\u0/IP [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[13]),
        .Q(\u0/IP [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[14]),
        .Q(\u0/IP [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[15]),
        .Q(\u0/IP [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[16]),
        .Q(\u0/IP [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[17]),
        .Q(\u0/IP [59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[18]),
        .Q(\u0/IP [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[19]),
        .Q(\u0/IP [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[1]),
        .Q(\u0/IP [57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[20]),
        .Q(\u0/IP [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[21]),
        .Q(\u0/IP [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[22]),
        .Q(\u0/IP [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[23]),
        .Q(\u0/IP [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[24]),
        .Q(\u0/IP [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[25]),
        .Q(\u0/IP [60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[26]),
        .Q(\u0/IP [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[27]),
        .Q(\u0/IP [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[28]),
        .Q(\u0/IP [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[29]),
        .Q(\u0/IP [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[2]),
        .Q(\u0/IP [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[30]),
        .Q(\u0/IP [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[31]),
        .Q(\u0/IP [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[32]),
        .Q(\u0/IP [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[33]),
        .Q(\u0/IP [61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[34]),
        .Q(\u0/IP [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[35]),
        .Q(\u0/IP [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[36]),
        .Q(\u0/IP [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[37]),
        .Q(\u0/IP [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[38]),
        .Q(\u0/IP [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[39]),
        .Q(\u0/IP [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[3]),
        .Q(\u0/IP [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[40]),
        .Q(\u0/IP [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[41]),
        .Q(\u0/IP [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[42]),
        .Q(\u0/IP [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[43]),
        .Q(\u0/IP [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[44]),
        .Q(\u0/IP [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[45]),
        .Q(\u0/IP [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[46]),
        .Q(\u0/IP [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[47]),
        .Q(\u0/IP [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[48]),
        .Q(\u0/IP [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[49]),
        .Q(\u0/IP [63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[4]),
        .Q(\u0/IP [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[50]),
        .Q(\u0/IP [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[51]),
        .Q(\u0/IP [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[52]),
        .Q(\u0/IP [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[53]),
        .Q(\u0/IP [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[54]),
        .Q(\u0/IP [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[55]),
        .Q(\u0/IP [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[56]),
        .Q(\u0/IP [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[57]),
        .Q(\u0/IP [64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[58]),
        .Q(\u0/IP [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[59]),
        .Q(\u0/IP [56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[5]),
        .Q(\u0/IP [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[60]),
        .Q(\u0/IP [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[61]),
        .Q(\u0/IP [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[62]),
        .Q(\u0/IP [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[63]),
        .Q(\u0/IP [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[6]),
        .Q(\u0/IP [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[7]),
        .Q(\u0/IP [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[8]),
        .Q(\u0/IP [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desIn_r_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(desIn[9]),
        .Q(\u0/IP [58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[0]_i_1 
       (.I0(\u0/out15 [25]),
        .I1(\u0/L14 [25]),
        .O(\u0/FP [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[10]_i_1 
       (.I0(\u0/out15 [18]),
        .I1(\u0/L14 [18]),
        .O(\u0/FP [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[12]_i_1 
       (.I0(\u0/out15 [10]),
        .I1(\u0/L14 [10]),
        .O(\u0/FP [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[14]_i_1 
       (.I0(\u0/out15 [2]),
        .I1(\u0/L14 [2]),
        .O(\u0/FP [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[16]_i_1 
       (.I0(\u0/out15 [27]),
        .I1(\u0/L14 [27]),
        .O(\u0/FP [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[18]_i_1 
       (.I0(\u0/out15 [19]),
        .I1(\u0/L14 [19]),
        .O(\u0/FP [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[20]_i_1 
       (.I0(\u0/out15 [11]),
        .I1(\u0/L14 [11]),
        .O(\u0/FP [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[22]_i_1 
       (.I0(\u0/out15 [3]),
        .I1(\u0/L14 [3]),
        .O(\u0/FP [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[24]_i_1 
       (.I0(\u0/out15 [28]),
        .I1(\u0/L14 [28]),
        .O(\u0/FP [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[26]_i_1 
       (.I0(\u0/out15 [20]),
        .I1(\u0/L14 [20]),
        .O(\u0/FP [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[28]_i_1 
       (.I0(\u0/out15 [12]),
        .I1(\u0/L14 [12]),
        .O(\u0/FP [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[2]_i_1 
       (.I0(\u0/out15 [17]),
        .I1(\u0/L14 [17]),
        .O(\u0/FP [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[30]_i_1 
       (.I0(\u0/out15 [4]),
        .I1(\u0/L14 [4]),
        .O(\u0/FP [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[32]_i_1 
       (.I0(\u0/out15 [29]),
        .I1(\u0/L14 [29]),
        .O(\u0/FP [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[34]_i_1 
       (.I0(\u0/out15 [21]),
        .I1(\u0/L14 [21]),
        .O(\u0/FP [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[36]_i_1 
       (.I0(\u0/out15 [13]),
        .I1(\u0/L14 [13]),
        .O(\u0/FP [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[38]_i_1 
       (.I0(\u0/out15 [5]),
        .I1(\u0/L14 [5]),
        .O(\u0/FP [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[40]_i_1 
       (.I0(\u0/out15 [30]),
        .I1(\u0/L14 [30]),
        .O(\u0/FP [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[42]_i_1 
       (.I0(\u0/out15 [22]),
        .I1(\u0/L14 [22]),
        .O(\u0/FP [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[44]_i_1 
       (.I0(\u0/out15 [14]),
        .I1(\u0/L14 [14]),
        .O(\u0/FP [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[46]_i_1 
       (.I0(\u0/out15 [6]),
        .I1(\u0/L14 [6]),
        .O(\u0/FP [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[48]_i_1 
       (.I0(\u0/out15 [31]),
        .I1(\u0/L14 [31]),
        .O(\u0/FP [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[4]_i_1 
       (.I0(\u0/out15 [9]),
        .I1(\u0/L14 [9]),
        .O(\u0/FP [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[50]_i_1 
       (.I0(\u0/out15 [23]),
        .I1(\u0/L14 [23]),
        .O(\u0/FP [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[52]_i_1 
       (.I0(\u0/out15 [15]),
        .I1(\u0/L14 [15]),
        .O(\u0/FP [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[54]_i_1 
       (.I0(\u0/out15 [7]),
        .I1(\u0/L14 [7]),
        .O(\u0/FP [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[56]_i_1 
       (.I0(\u0/out15 [32]),
        .I1(\u0/L14 [32]),
        .O(\u0/FP [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[58]_i_1 
       (.I0(\u0/out15 [24]),
        .I1(\u0/L14 [24]),
        .O(\u0/FP [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[60]_i_1 
       (.I0(\u0/out15 [16]),
        .I1(\u0/L14 [16]),
        .O(\u0/FP [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[62]_i_1 
       (.I0(\u0/out15 [8]),
        .I1(\u0/L14 [8]),
        .O(\u0/FP [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[6]_i_1 
       (.I0(\u0/out15 [1]),
        .I1(\u0/L14 [1]),
        .O(\u0/FP [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u0/desOut[8]_i_1 
       (.I0(\u0/out15 [26]),
        .I1(\u0/L14 [26]),
        .O(\u0/FP [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [25]),
        .Q(stage1_out[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [18]),
        .Q(stage1_out[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [50]),
        .Q(stage1_out[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [10]),
        .Q(stage1_out[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [42]),
        .Q(stage1_out[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [2]),
        .Q(stage1_out[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [34]),
        .Q(stage1_out[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [27]),
        .Q(stage1_out[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [59]),
        .Q(stage1_out[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [19]),
        .Q(stage1_out[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [51]),
        .Q(stage1_out[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [57]),
        .Q(stage1_out[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [11]),
        .Q(stage1_out[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [43]),
        .Q(stage1_out[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [3]),
        .Q(stage1_out[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [35]),
        .Q(stage1_out[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [28]),
        .Q(stage1_out[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [60]),
        .Q(stage1_out[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [20]),
        .Q(stage1_out[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [52]),
        .Q(stage1_out[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [12]),
        .Q(stage1_out[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [44]),
        .Q(stage1_out[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [17]),
        .Q(stage1_out[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [4]),
        .Q(stage1_out[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [36]),
        .Q(stage1_out[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [29]),
        .Q(stage1_out[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [61]),
        .Q(stage1_out[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [21]),
        .Q(stage1_out[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [53]),
        .Q(stage1_out[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [13]),
        .Q(stage1_out[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [45]),
        .Q(stage1_out[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [5]),
        .Q(stage1_out[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [37]),
        .Q(stage1_out[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [49]),
        .Q(stage1_out[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [30]),
        .Q(stage1_out[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [62]),
        .Q(stage1_out[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [22]),
        .Q(stage1_out[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [54]),
        .Q(stage1_out[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [14]),
        .Q(stage1_out[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [46]),
        .Q(stage1_out[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [6]),
        .Q(stage1_out[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [38]),
        .Q(stage1_out[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [31]),
        .Q(stage1_out[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [63]),
        .Q(stage1_out[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [9]),
        .Q(stage1_out[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [23]),
        .Q(stage1_out[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [55]),
        .Q(stage1_out[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [15]),
        .Q(stage1_out[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [47]),
        .Q(stage1_out[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [7]),
        .Q(stage1_out[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [39]),
        .Q(stage1_out[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [32]),
        .Q(stage1_out[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [64]),
        .Q(stage1_out[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [24]),
        .Q(stage1_out[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [56]),
        .Q(stage1_out[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [41]),
        .Q(stage1_out[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [16]),
        .Q(stage1_out[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [48]),
        .Q(stage1_out[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [8]),
        .Q(stage1_out[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [40]),
        .Q(stage1_out[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [1]),
        .Q(stage1_out[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [33]),
        .Q(stage1_out[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [26]),
        .Q(stage1_out[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/desOut_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/FP [58]),
        .Q(stage1_out[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[0]),
        .Q(\u0/key_r [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[10]),
        .Q(\u0/key_r [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[11]),
        .Q(\u0/key_r [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[12]),
        .Q(\u0/key_r [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[13]),
        .Q(\u0/key_r [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[14]),
        .Q(\u0/key_r [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[15]),
        .Q(\u0/key_r [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[16]),
        .Q(\u0/key_r [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[17]),
        .Q(\u0/key_r [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[18]),
        .Q(\u0/key_r [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[19]),
        .Q(\u0/key_r [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[1]),
        .Q(\u0/key_r [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[20]),
        .Q(\u0/key_r [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[21]),
        .Q(\u0/key_r [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[22]),
        .Q(\u0/key_r [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[23]),
        .Q(\u0/key_r [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[24]),
        .Q(\u0/key_r [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[25]),
        .Q(\u0/key_r [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[26]),
        .Q(\u0/key_r [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[27]),
        .Q(\u0/key_r [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[28]),
        .Q(\u0/key_r [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[29]),
        .Q(\u0/key_r [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[2]),
        .Q(\u0/key_r [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[30]),
        .Q(\u0/key_r [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[31]),
        .Q(\u0/key_r [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[32]),
        .Q(\u0/key_r [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[33]),
        .Q(\u0/key_r [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[34]),
        .Q(\u0/key_r [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[35]),
        .Q(\u0/key_r [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[36]),
        .Q(\u0/key_r [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[37]),
        .Q(\u0/key_r [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[38]),
        .Q(\u0/key_r [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[39]),
        .Q(\u0/key_r [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[3]),
        .Q(\u0/key_r [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[40]),
        .Q(\u0/key_r [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[41]),
        .Q(\u0/key_r [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[42]),
        .Q(\u0/key_r [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[43]),
        .Q(\u0/key_r [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[44]),
        .Q(\u0/key_r [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[45]),
        .Q(\u0/key_r [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[46]),
        .Q(\u0/key_r [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[47]),
        .Q(\u0/key_r [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[48]),
        .Q(\u0/key_r [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[49]),
        .Q(\u0/key_r [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[4]),
        .Q(\u0/key_r [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[50]),
        .Q(\u0/key_r [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[51]),
        .Q(\u0/key_r [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[52]),
        .Q(\u0/key_r [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[53]),
        .Q(\u0/key_r [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[54]),
        .Q(\u0/key_r [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[55]),
        .Q(\u0/key_r [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[5]),
        .Q(\u0/key_r [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[6]),
        .Q(\u0/key_r [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[7]),
        .Q(\u0/key_r [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[8]),
        .Q(\u0/key_r [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/key_r_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_a[9]),
        .Q(\u0/key_r [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [0]),
        .Q(\u0/uk/K_r0_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [10]),
        .Q(\u0/uk/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [11]),
        .Q(\u0/uk/p_14_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [12]),
        .Q(\u0/uk/p_38_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [13]),
        .Q(\u0/uk/p_7_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [14]),
        .Q(\u0/uk/p_36_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [15]),
        .Q(\u0/uk/p_25_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [16]),
        .Q(\u0/uk/p_27_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [17]),
        .Q(\u0/uk/K_r0_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [18]),
        .Q(\u0/uk/p_37_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [19]),
        .Q(\u0/uk/K_r0_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [1]),
        .Q(\u0/uk/K_r0_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [20]),
        .Q(\u0/uk/p_2_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [21]),
        .Q(\u0/uk/p_24_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [22]),
        .Q(\u0/uk/K_r0_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [23]),
        .Q(\u0/uk/p_30_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [24]),
        .Q(\u0/uk/p_3_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [25]),
        .Q(\u0/uk/K_r0_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [26]),
        .Q(\u0/uk/p_9_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [27]),
        .Q(\u0/uk/p_5_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [28]),
        .Q(\u0/uk/p_20_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [29]),
        .Q(\u0/uk/p_31_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [2]),
        .Q(\u0/uk/K_r0_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [30]),
        .Q(\u0/uk/p_22_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [31]),
        .Q(\u0/uk/K_r0_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [32]),
        .Q(\u0/uk/K_r0_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [33]),
        .Q(\u0/uk/p_39_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [34]),
        .Q(\u0/uk/p_6_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [35]),
        .Q(\u0/uk/K_r0_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [36]),
        .Q(\u0/uk/K_r0_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [37]),
        .Q(\u0/uk/p_26_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [38]),
        .Q(\u0/uk/p_18_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [39]),
        .Q(\u0/uk/p_12_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [3]),
        .Q(\u0/uk/p_11_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [40]),
        .Q(\u0/uk/p_8_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [41]),
        .Q(\u0/uk/p_13_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [42]),
        .Q(\u0/uk/p_29_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [43]),
        .Q(\u0/uk/p_17_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [44]),
        .Q(\u0/uk/p_19_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [45]),
        .Q(\u0/uk/p_33_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [46]),
        .Q(\u0/uk/p_1_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [47]),
        .Q(\u0/uk/p_15_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [48]),
        .Q(\u0/uk/p_4_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [49]),
        .Q(\u0/uk/p_34_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [4]),
        .Q(\u0/uk/K_r0_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [50]),
        .Q(\u0/uk/p_28_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [51]),
        .Q(\u0/uk/p_35_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [52]),
        .Q(\u0/uk/K_r0_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [53]),
        .Q(\u0/uk/K_r0_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [54]),
        .Q(\u0/uk/p_40_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [55]),
        .Q(\u0/uk/K_r0_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [5]),
        .Q(\u0/uk/p_10_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [6]),
        .Q(\u0/uk/p_16_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [7]),
        .Q(\u0/uk/p_21_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [8]),
        .Q(\u0/uk/p_32_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r0_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/key_r [9]),
        .Q(\u0/uk/p_23_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [0]),
        .Q(\u0/uk/K_r10 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [10]),
        .Q(\u0/uk/K_r10 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [11]),
        .Q(\u0/uk/K_r10 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [12]),
        .Q(\u0/uk/K_r10 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [13]),
        .Q(\u0/uk/K_r10 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [14]),
        .Q(\u0/uk/K_r10 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [15]),
        .Q(\u0/uk/K_r10 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [16]),
        .Q(\u0/uk/K_r10 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [17]),
        .Q(\u0/uk/K_r10 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [18]),
        .Q(\u0/uk/K_r10 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [19]),
        .Q(\u0/uk/K_r10 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [1]),
        .Q(\u0/uk/K_r10 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [20]),
        .Q(\u0/uk/K_r10 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [21]),
        .Q(\u0/uk/K_r10 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [22]),
        .Q(\u0/uk/K_r10 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [23]),
        .Q(\u0/uk/K_r10 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [24]),
        .Q(\u0/uk/K_r10 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [25]),
        .Q(\u0/uk/K_r10 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [26]),
        .Q(\u0/uk/K_r10 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [27]),
        .Q(\u0/uk/K_r10 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [28]),
        .Q(\u0/uk/K_r10 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [29]),
        .Q(\u0/uk/K_r10 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [2]),
        .Q(\u0/uk/K_r10 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [30]),
        .Q(\u0/uk/K_r10 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [31]),
        .Q(\u0/uk/K_r10 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [32]),
        .Q(\u0/uk/K_r10 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [33]),
        .Q(\u0/uk/K_r10 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [34]),
        .Q(\u0/uk/K_r10 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [35]),
        .Q(\u0/uk/K_r10 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [36]),
        .Q(\u0/uk/K_r10 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [37]),
        .Q(\u0/uk/K_r10 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [38]),
        .Q(\u0/uk/K_r10 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [39]),
        .Q(\u0/uk/K_r10 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [3]),
        .Q(\u0/uk/K_r10 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [40]),
        .Q(\u0/uk/K_r10 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [41]),
        .Q(\u0/uk/K_r10 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [42]),
        .Q(\u0/uk/K_r10 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [43]),
        .Q(\u0/uk/K_r10 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [44]),
        .Q(\u0/uk/K_r10 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [45]),
        .Q(\u0/uk/K_r10 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [46]),
        .Q(\u0/uk/K_r10 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [47]),
        .Q(\u0/uk/K_r10 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [48]),
        .Q(\u0/uk/K_r10 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [49]),
        .Q(\u0/uk/K_r10 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [4]),
        .Q(\u0/uk/K_r10 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [50]),
        .Q(\u0/uk/K_r10 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [51]),
        .Q(\u0/uk/K_r10 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [52]),
        .Q(\u0/uk/K_r10 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [53]),
        .Q(\u0/uk/K_r10 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [54]),
        .Q(\u0/uk/K_r10 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [55]),
        .Q(\u0/uk/K_r10 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [5]),
        .Q(\u0/uk/K_r10 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [6]),
        .Q(\u0/uk/K_r10 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [7]),
        .Q(\u0/uk/K_r10 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [8]),
        .Q(\u0/uk/K_r10 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r10_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r9 [9]),
        .Q(\u0/uk/K_r10 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [0]),
        .Q(\u0/uk/K_r11 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [10]),
        .Q(\u0/uk/K_r11 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [11]),
        .Q(\u0/uk/K_r11 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [12]),
        .Q(\u0/uk/K_r11 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [13]),
        .Q(\u0/uk/K_r11 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [14]),
        .Q(\u0/uk/K_r11 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [15]),
        .Q(\u0/uk/K_r11 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [16]),
        .Q(\u0/uk/K_r11 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [17]),
        .Q(\u0/uk/K_r11 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [18]),
        .Q(\u0/uk/K_r11 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [19]),
        .Q(\u0/uk/K_r11 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [1]),
        .Q(\u0/uk/K_r11 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [20]),
        .Q(\u0/uk/K_r11 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [21]),
        .Q(\u0/uk/K_r11 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [22]),
        .Q(\u0/uk/K_r11 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [23]),
        .Q(\u0/uk/K_r11 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [24]),
        .Q(\u0/uk/K_r11 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [25]),
        .Q(\u0/uk/K_r11 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [26]),
        .Q(\u0/uk/K_r11 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [27]),
        .Q(\u0/uk/K_r11 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [28]),
        .Q(\u0/uk/K_r11 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [29]),
        .Q(\u0/uk/K_r11 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [2]),
        .Q(\u0/uk/K_r11 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [30]),
        .Q(\u0/uk/K_r11 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [31]),
        .Q(\u0/uk/K_r11 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [32]),
        .Q(\u0/uk/K_r11 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [33]),
        .Q(\u0/uk/K_r11 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [34]),
        .Q(\u0/uk/K_r11 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [35]),
        .Q(\u0/uk/K_r11 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [36]),
        .Q(\u0/uk/K_r11 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [37]),
        .Q(\u0/uk/K_r11 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [38]),
        .Q(\u0/uk/K_r11 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [39]),
        .Q(\u0/uk/K_r11 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [3]),
        .Q(\u0/uk/K_r11 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [40]),
        .Q(\u0/uk/K_r11 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [41]),
        .Q(\u0/uk/K_r11 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [42]),
        .Q(\u0/uk/K_r11 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [43]),
        .Q(\u0/uk/K_r11 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [44]),
        .Q(\u0/uk/K_r11 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [45]),
        .Q(\u0/uk/K_r11 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [46]),
        .Q(\u0/uk/K_r11 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [47]),
        .Q(\u0/uk/K_r11 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [48]),
        .Q(\u0/uk/K_r11 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [49]),
        .Q(\u0/uk/K_r11 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [4]),
        .Q(\u0/uk/K_r11 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [50]),
        .Q(\u0/uk/K_r11 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [51]),
        .Q(\u0/uk/K_r11 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [52]),
        .Q(\u0/uk/K_r11 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [53]),
        .Q(\u0/uk/K_r11 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [54]),
        .Q(\u0/uk/K_r11 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [55]),
        .Q(\u0/uk/K_r11 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [5]),
        .Q(\u0/uk/K_r11 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [6]),
        .Q(\u0/uk/K_r11 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [7]),
        .Q(\u0/uk/K_r11 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [8]),
        .Q(\u0/uk/K_r11 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r11_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r10 [9]),
        .Q(\u0/uk/K_r11 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [0]),
        .Q(\u0/uk/K_r12 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [10]),
        .Q(\u0/uk/K_r12 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [11]),
        .Q(\u0/uk/K_r12 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [12]),
        .Q(\u0/uk/K_r12 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [13]),
        .Q(\u0/uk/K_r12 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [14]),
        .Q(\u0/uk/K_r12 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [15]),
        .Q(\u0/uk/K_r12 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [16]),
        .Q(\u0/uk/K_r12 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [17]),
        .Q(\u0/uk/K_r12 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [18]),
        .Q(\u0/uk/K_r12 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [19]),
        .Q(\u0/uk/K_r12 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [1]),
        .Q(\u0/uk/K_r12 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [20]),
        .Q(\u0/uk/K_r12 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [21]),
        .Q(\u0/uk/K_r12 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [22]),
        .Q(\u0/uk/K_r12 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [23]),
        .Q(\u0/uk/K_r12 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [24]),
        .Q(\u0/uk/K_r12 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [25]),
        .Q(\u0/uk/K_r12 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [26]),
        .Q(\u0/uk/K_r12 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [27]),
        .Q(\u0/uk/K_r12 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [28]),
        .Q(\u0/uk/K_r12 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [29]),
        .Q(\u0/uk/K_r12 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [2]),
        .Q(\u0/uk/K_r12 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [30]),
        .Q(\u0/uk/K_r12 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [31]),
        .Q(\u0/uk/K_r12 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [32]),
        .Q(\u0/uk/K_r12 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [33]),
        .Q(\u0/uk/K_r12 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [34]),
        .Q(\u0/uk/K_r12 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [35]),
        .Q(\u0/uk/K_r12 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [36]),
        .Q(\u0/uk/K_r12 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [37]),
        .Q(\u0/uk/K_r12 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [38]),
        .Q(\u0/uk/K_r12 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [39]),
        .Q(\u0/uk/K_r12 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [3]),
        .Q(\u0/uk/K_r12 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [40]),
        .Q(\u0/uk/K_r12 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [41]),
        .Q(\u0/uk/K_r12 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [42]),
        .Q(\u0/uk/K_r12 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [43]),
        .Q(\u0/uk/K_r12 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [44]),
        .Q(\u0/uk/K_r12 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [45]),
        .Q(\u0/uk/K_r12 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [46]),
        .Q(\u0/uk/K_r12 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [47]),
        .Q(\u0/uk/K_r12 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [48]),
        .Q(\u0/uk/K_r12 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [49]),
        .Q(\u0/uk/K_r12 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [4]),
        .Q(\u0/uk/K_r12 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [50]),
        .Q(\u0/uk/K_r12 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [51]),
        .Q(\u0/uk/K_r12 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [52]),
        .Q(\u0/uk/K_r12 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [53]),
        .Q(\u0/uk/K_r12 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [54]),
        .Q(\u0/uk/K_r12 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [55]),
        .Q(\u0/uk/K_r12 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [5]),
        .Q(\u0/uk/K_r12 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [6]),
        .Q(\u0/uk/K_r12 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [7]),
        .Q(\u0/uk/K_r12 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [8]),
        .Q(\u0/uk/K_r12 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r12_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r11 [9]),
        .Q(\u0/uk/K_r12 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [0]),
        .Q(\u0/uk/K_r13 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [10]),
        .Q(\u0/uk/K_r13 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [11]),
        .Q(\u0/uk/K_r13 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [12]),
        .Q(\u0/uk/K_r13 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [13]),
        .Q(\u0/uk/K_r13 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [14]),
        .Q(\u0/uk/K_r13 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [15]),
        .Q(\u0/uk/K_r13 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [16]),
        .Q(\u0/uk/K_r13 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [17]),
        .Q(\u0/uk/K_r13 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [18]),
        .Q(\u0/uk/K_r13 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [19]),
        .Q(\u0/uk/K_r13 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [1]),
        .Q(\u0/uk/K_r13 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [20]),
        .Q(\u0/uk/K_r13 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [21]),
        .Q(\u0/uk/K_r13 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [22]),
        .Q(\u0/uk/K_r13 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [23]),
        .Q(\u0/uk/K_r13 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [24]),
        .Q(\u0/uk/K_r13 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [25]),
        .Q(\u0/uk/K_r13 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [26]),
        .Q(\u0/uk/K_r13 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [27]),
        .Q(\u0/uk/K_r13 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [28]),
        .Q(\u0/uk/K_r13 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [29]),
        .Q(\u0/uk/K_r13 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [2]),
        .Q(\u0/uk/K_r13 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [30]),
        .Q(\u0/uk/K_r13 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [31]),
        .Q(\u0/uk/K_r13 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [32]),
        .Q(\u0/uk/K_r13 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [33]),
        .Q(\u0/uk/K_r13 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [34]),
        .Q(\u0/uk/K_r13 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [35]),
        .Q(\u0/uk/K_r13 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [36]),
        .Q(\u0/uk/K_r13 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [37]),
        .Q(\u0/uk/K_r13 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [38]),
        .Q(\u0/uk/K_r13 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [39]),
        .Q(\u0/uk/K_r13 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [3]),
        .Q(\u0/uk/K_r13 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [40]),
        .Q(\u0/uk/K_r13 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [41]),
        .Q(\u0/uk/K_r13 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [42]),
        .Q(\u0/uk/K_r13 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [43]),
        .Q(\u0/uk/K_r13 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [44]),
        .Q(\u0/uk/K_r13 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [45]),
        .Q(\u0/uk/K_r13 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [46]),
        .Q(\u0/uk/K_r13 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [47]),
        .Q(\u0/uk/K_r13 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [48]),
        .Q(\u0/uk/K_r13 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [49]),
        .Q(\u0/uk/K_r13 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [4]),
        .Q(\u0/uk/K_r13 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [50]),
        .Q(\u0/uk/K_r13 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [51]),
        .Q(\u0/uk/K_r13 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [52]),
        .Q(\u0/uk/K_r13 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [53]),
        .Q(\u0/uk/K_r13 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [54]),
        .Q(\u0/uk/K_r13 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [55]),
        .Q(\u0/uk/K_r13 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [5]),
        .Q(\u0/uk/K_r13 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [6]),
        .Q(\u0/uk/K_r13 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [7]),
        .Q(\u0/uk/K_r13 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [8]),
        .Q(\u0/uk/K_r13 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r13_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r12 [9]),
        .Q(\u0/uk/K_r13 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [0]),
        .Q(\u0/uk/K_r14_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [10]),
        .Q(\u0/uk/K_r14_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [11]),
        .Q(\u0/uk/K_r14_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [12]),
        .Q(\u0/uk/K_r14_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [13]),
        .Q(\u0/uk/K_r14_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [14]),
        .Q(\u0/uk/K_r14_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [15]),
        .Q(\u0/uk/K_r14_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [16]),
        .Q(\u0/uk/K_r14_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [17]),
        .Q(\u0/uk/K_r14_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [18]),
        .Q(\u0/uk/K_r14_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [19]),
        .Q(\u0/uk/K_r14_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [1]),
        .Q(\u0/uk/K_r14_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [20]),
        .Q(\u0/uk/K_r14_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [21]),
        .Q(\u0/uk/K_r14_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [22]),
        .Q(\u0/uk/K_r14_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [23]),
        .Q(\u0/uk/K_r14_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [24]),
        .Q(\u0/uk/K_r14_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [25]),
        .Q(\u0/uk/K_r14_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [26]),
        .Q(\u0/uk/K_r14_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [27]),
        .Q(\u0/uk/K_r14_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [28]),
        .Q(\u0/uk/K_r14_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [29]),
        .Q(\u0/uk/K_r14_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [2]),
        .Q(\u0/uk/K_r14_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [30]),
        .Q(\u0/uk/K_r14_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [31]),
        .Q(\u0/uk/K_r14_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [32]),
        .Q(\u0/uk/K_r14_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [33]),
        .Q(\u0/uk/K_r14_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [34]),
        .Q(\u0/uk/K_r14_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [35]),
        .Q(\u0/uk/K_r14_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [36]),
        .Q(\u0/uk/K_r14_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [37]),
        .Q(\u0/uk/K_r14_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [38]),
        .Q(\u0/uk/K_r14_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [39]),
        .Q(\u0/uk/K_r14_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [3]),
        .Q(\u0/uk/K_r14_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [40]),
        .Q(\u0/uk/K_r14_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [41]),
        .Q(\u0/uk/K_r14_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [42]),
        .Q(\u0/uk/K_r14_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [43]),
        .Q(\u0/uk/K_r14_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [44]),
        .Q(\u0/uk/K_r14_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [45]),
        .Q(\u0/uk/K_r14_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [46]),
        .Q(\u0/uk/K_r14_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [47]),
        .Q(\u0/uk/K_r14_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [48]),
        .Q(\u0/uk/K_r14_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [49]),
        .Q(\u0/uk/K_r14_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [4]),
        .Q(\u0/uk/K_r14_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [50]),
        .Q(\u0/uk/K_r14_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [51]),
        .Q(\u0/uk/K_r14_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [52]),
        .Q(\u0/uk/K_r14_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [53]),
        .Q(\u0/uk/K_r14_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [54]),
        .Q(\u0/uk/K_r14_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [55]),
        .Q(\u0/uk/K_r14_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [5]),
        .Q(\u0/uk/K_r14_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [6]),
        .Q(\u0/uk/K_r14_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [7]),
        .Q(\u0/uk/K_r14_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [8]),
        .Q(\u0/uk/K_r14_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r14_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r13 [9]),
        .Q(\u0/uk/K_r14_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_ ),
        .Q(\u0/uk/K_r1 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_0_in ),
        .Q(\u0/uk/K_r1 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_14_in ),
        .Q(\u0/uk/K_r1 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_38_in ),
        .Q(\u0/uk/K_r1 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_7_in ),
        .Q(\u0/uk/K_r1 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_36_in ),
        .Q(\u0/uk/K_r1 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_25_in ),
        .Q(\u0/uk/K_r1 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_27_in ),
        .Q(\u0/uk/K_r1 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[17] ),
        .Q(\u0/uk/K_r1 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_37_in ),
        .Q(\u0/uk/K_r1 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[19] ),
        .Q(\u0/uk/K_r1 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[1] ),
        .Q(\u0/uk/K_r1 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_2_in ),
        .Q(\u0/uk/K_r1 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_24_in ),
        .Q(\u0/uk/K_r1 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[22] ),
        .Q(\u0/uk/K_r1 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_30_in ),
        .Q(\u0/uk/K_r1 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_3_in ),
        .Q(\u0/uk/K_r1 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[25] ),
        .Q(\u0/uk/K_r1 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_9_in ),
        .Q(\u0/uk/K_r1 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_5_in ),
        .Q(\u0/uk/K_r1 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_20_in ),
        .Q(\u0/uk/K_r1 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_31_in ),
        .Q(\u0/uk/K_r1 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[2] ),
        .Q(\u0/uk/K_r1 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_22_in ),
        .Q(\u0/uk/K_r1 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[31] ),
        .Q(\u0/uk/K_r1 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[32] ),
        .Q(\u0/uk/K_r1 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_39_in ),
        .Q(\u0/uk/K_r1 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_6_in ),
        .Q(\u0/uk/K_r1 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[35] ),
        .Q(\u0/uk/K_r1 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[36] ),
        .Q(\u0/uk/K_r1 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_26_in ),
        .Q(\u0/uk/K_r1 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_18_in ),
        .Q(\u0/uk/K_r1 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_12_in ),
        .Q(\u0/uk/K_r1 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_11_in ),
        .Q(\u0/uk/K_r1 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_8_in ),
        .Q(\u0/uk/K_r1 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_13_in ),
        .Q(\u0/uk/K_r1 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_29_in ),
        .Q(\u0/uk/K_r1 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_17_in ),
        .Q(\u0/uk/K_r1 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_19_in ),
        .Q(\u0/uk/K_r1 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_33_in ),
        .Q(\u0/uk/K_r1 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_1_in ),
        .Q(\u0/uk/K_r1 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_15_in ),
        .Q(\u0/uk/K_r1 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_4_in ),
        .Q(\u0/uk/K_r1 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_34_in ),
        .Q(\u0/uk/K_r1 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[4] ),
        .Q(\u0/uk/K_r1 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_28_in ),
        .Q(\u0/uk/K_r1 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_35_in ),
        .Q(\u0/uk/K_r1 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[52] ),
        .Q(\u0/uk/K_r1 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[53] ),
        .Q(\u0/uk/K_r1 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_40_in ),
        .Q(\u0/uk/K_r1 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r0_reg_n_0_[55] ),
        .Q(\u0/uk/K_r1 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_10_in ),
        .Q(\u0/uk/K_r1 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_16_in ),
        .Q(\u0/uk/K_r1 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_21_in ),
        .Q(\u0/uk/K_r1 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_32_in ),
        .Q(\u0/uk/K_r1 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_23_in ),
        .Q(\u0/uk/K_r1 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [0]),
        .Q(\u0/uk/K_r2 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [10]),
        .Q(\u0/uk/K_r2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [11]),
        .Q(\u0/uk/K_r2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [12]),
        .Q(\u0/uk/K_r2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [13]),
        .Q(\u0/uk/K_r2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [14]),
        .Q(\u0/uk/K_r2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [15]),
        .Q(\u0/uk/K_r2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [16]),
        .Q(\u0/uk/K_r2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [17]),
        .Q(\u0/uk/K_r2 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [18]),
        .Q(\u0/uk/K_r2 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [19]),
        .Q(\u0/uk/K_r2 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [1]),
        .Q(\u0/uk/K_r2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [20]),
        .Q(\u0/uk/K_r2 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [21]),
        .Q(\u0/uk/K_r2 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [22]),
        .Q(\u0/uk/K_r2 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [23]),
        .Q(\u0/uk/K_r2 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [24]),
        .Q(\u0/uk/K_r2 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [25]),
        .Q(\u0/uk/K_r2 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [26]),
        .Q(\u0/uk/K_r2 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [27]),
        .Q(\u0/uk/K_r2 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [28]),
        .Q(\u0/uk/K_r2 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [29]),
        .Q(\u0/uk/K_r2 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [2]),
        .Q(\u0/uk/K_r2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [30]),
        .Q(\u0/uk/K_r2 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [31]),
        .Q(\u0/uk/K_r2 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [32]),
        .Q(\u0/uk/K_r2 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [33]),
        .Q(\u0/uk/K_r2 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [34]),
        .Q(\u0/uk/K_r2 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [35]),
        .Q(\u0/uk/K_r2 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [36]),
        .Q(\u0/uk/K_r2 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [37]),
        .Q(\u0/uk/K_r2 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [38]),
        .Q(\u0/uk/K_r2 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [39]),
        .Q(\u0/uk/K_r2 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [3]),
        .Q(\u0/uk/K_r2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [40]),
        .Q(\u0/uk/K_r2 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [41]),
        .Q(\u0/uk/K_r2 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [42]),
        .Q(\u0/uk/K_r2 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [43]),
        .Q(\u0/uk/K_r2 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [44]),
        .Q(\u0/uk/K_r2 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [45]),
        .Q(\u0/uk/K_r2 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [46]),
        .Q(\u0/uk/K_r2 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [47]),
        .Q(\u0/uk/K_r2 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [48]),
        .Q(\u0/uk/K_r2 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [49]),
        .Q(\u0/uk/K_r2 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [4]),
        .Q(\u0/uk/K_r2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [50]),
        .Q(\u0/uk/K_r2 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [51]),
        .Q(\u0/uk/K_r2 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [52]),
        .Q(\u0/uk/K_r2 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [53]),
        .Q(\u0/uk/K_r2 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [54]),
        .Q(\u0/uk/K_r2 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [55]),
        .Q(\u0/uk/K_r2 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [5]),
        .Q(\u0/uk/K_r2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [6]),
        .Q(\u0/uk/K_r2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [7]),
        .Q(\u0/uk/K_r2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [8]),
        .Q(\u0/uk/K_r2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r2_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r1 [9]),
        .Q(\u0/uk/K_r2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [0]),
        .Q(\u0/uk/K_r3 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [10]),
        .Q(\u0/uk/K_r3 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [11]),
        .Q(\u0/uk/K_r3 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [12]),
        .Q(\u0/uk/K_r3 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [13]),
        .Q(\u0/uk/K_r3 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [14]),
        .Q(\u0/uk/K_r3 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [15]),
        .Q(\u0/uk/K_r3 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [16]),
        .Q(\u0/uk/K_r3 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [17]),
        .Q(\u0/uk/K_r3 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [18]),
        .Q(\u0/uk/K_r3 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [19]),
        .Q(\u0/uk/K_r3 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [1]),
        .Q(\u0/uk/K_r3 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [20]),
        .Q(\u0/uk/K_r3 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [21]),
        .Q(\u0/uk/K_r3 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [22]),
        .Q(\u0/uk/K_r3 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [23]),
        .Q(\u0/uk/K_r3 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [24]),
        .Q(\u0/uk/K_r3 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [25]),
        .Q(\u0/uk/K_r3 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [26]),
        .Q(\u0/uk/K_r3 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [27]),
        .Q(\u0/uk/K_r3 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [28]),
        .Q(\u0/uk/K_r3 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [29]),
        .Q(\u0/uk/K_r3 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [2]),
        .Q(\u0/uk/K_r3 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [30]),
        .Q(\u0/uk/K_r3 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [31]),
        .Q(\u0/uk/K_r3 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [32]),
        .Q(\u0/uk/K_r3 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [33]),
        .Q(\u0/uk/K_r3 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [34]),
        .Q(\u0/uk/K_r3 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [35]),
        .Q(\u0/uk/K_r3 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [36]),
        .Q(\u0/uk/K_r3 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [37]),
        .Q(\u0/uk/K_r3 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [38]),
        .Q(\u0/uk/K_r3 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [39]),
        .Q(\u0/uk/K_r3 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [3]),
        .Q(\u0/uk/K_r3 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [40]),
        .Q(\u0/uk/K_r3 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [41]),
        .Q(\u0/uk/K_r3 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [42]),
        .Q(\u0/uk/K_r3 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [43]),
        .Q(\u0/uk/K_r3 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [44]),
        .Q(\u0/uk/K_r3 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [45]),
        .Q(\u0/uk/K_r3 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [46]),
        .Q(\u0/uk/K_r3 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [47]),
        .Q(\u0/uk/K_r3 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [48]),
        .Q(\u0/uk/K_r3 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [49]),
        .Q(\u0/uk/K_r3 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [4]),
        .Q(\u0/uk/K_r3 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [50]),
        .Q(\u0/uk/K_r3 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [51]),
        .Q(\u0/uk/K_r3 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [52]),
        .Q(\u0/uk/K_r3 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [53]),
        .Q(\u0/uk/K_r3 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [54]),
        .Q(\u0/uk/K_r3 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [55]),
        .Q(\u0/uk/K_r3 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [5]),
        .Q(\u0/uk/K_r3 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [6]),
        .Q(\u0/uk/K_r3 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [7]),
        .Q(\u0/uk/K_r3 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [8]),
        .Q(\u0/uk/K_r3 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r3_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r2 [9]),
        .Q(\u0/uk/K_r3 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [0]),
        .Q(\u0/uk/K_r4_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [10]),
        .Q(\u0/uk/K_r4_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [11]),
        .Q(\u0/uk/K_r4_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [12]),
        .Q(\u0/uk/K_r4_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [13]),
        .Q(\u0/uk/K_r4_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [14]),
        .Q(\u0/uk/K_r4_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [15]),
        .Q(\u0/uk/K_r4_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [16]),
        .Q(\u0/uk/K_r4_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [17]),
        .Q(\u0/uk/K_r4_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [18]),
        .Q(\u0/uk/K_r4_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [19]),
        .Q(\u0/uk/K_r4_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [1]),
        .Q(\u0/uk/K_r4_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [20]),
        .Q(\u0/uk/K_r4_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [21]),
        .Q(\u0/uk/K_r4_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [22]),
        .Q(\u0/uk/K_r4_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [23]),
        .Q(\u0/uk/K_r4_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [24]),
        .Q(\u0/uk/K_r4_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [25]),
        .Q(\u0/uk/K_r4_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [26]),
        .Q(\u0/uk/K_r4_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [27]),
        .Q(\u0/uk/K_r4_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [28]),
        .Q(\u0/uk/K_r4_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [29]),
        .Q(\u0/uk/K_r4_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [2]),
        .Q(\u0/uk/K_r4_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [30]),
        .Q(\u0/uk/K_r4_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [31]),
        .Q(\u0/uk/K_r4_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [32]),
        .Q(\u0/uk/K_r4_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [33]),
        .Q(\u0/uk/K_r4_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [34]),
        .Q(\u0/uk/p_50_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [35]),
        .Q(\u0/uk/K_r4_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [36]),
        .Q(\u0/uk/K_r4_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [37]),
        .Q(\u0/uk/K_r4_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [38]),
        .Q(\u0/uk/K_r4_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [39]),
        .Q(\u0/uk/K_r4_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [3]),
        .Q(\u0/uk/K_r4_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [40]),
        .Q(\u0/uk/p_49_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [41]),
        .Q(\u0/uk/K_r4_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [42]),
        .Q(\u0/uk/K_r4_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [43]),
        .Q(\u0/uk/p_44_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [44]),
        .Q(\u0/uk/K_r4_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [45]),
        .Q(\u0/uk/K_r4_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [46]),
        .Q(\u0/uk/p_47_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [47]),
        .Q(\u0/uk/K_r4_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [48]),
        .Q(\u0/uk/K_r4_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [49]),
        .Q(\u0/uk/K_r4_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [4]),
        .Q(\u0/uk/K_r4_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [50]),
        .Q(\u0/uk/K_r4_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [51]),
        .Q(\u0/uk/K_r4_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [52]),
        .Q(\u0/uk/K_r4_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [53]),
        .Q(\u0/uk/p_51_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [54]),
        .Q(\u0/uk/K_r4_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [55]),
        .Q(\u0/uk/K_r4_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [5]),
        .Q(\u0/uk/K_r4_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [6]),
        .Q(\u0/uk/K_r4_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [7]),
        .Q(\u0/uk/K_r4_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [8]),
        .Q(\u0/uk/p_42_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r4_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r3 [9]),
        .Q(\u0/uk/K_r4_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_ ),
        .Q(\u0/uk/K_r5 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[10] ),
        .Q(\u0/uk/K_r5 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[11] ),
        .Q(\u0/uk/K_r5 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[12] ),
        .Q(\u0/uk/K_r5 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[13] ),
        .Q(\u0/uk/K_r5 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[14] ),
        .Q(\u0/uk/K_r5 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[15] ),
        .Q(\u0/uk/K_r5 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[16] ),
        .Q(\u0/uk/K_r5 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[17] ),
        .Q(\u0/uk/K_r5 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[18] ),
        .Q(\u0/uk/K_r5 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[19] ),
        .Q(\u0/uk/K_r5 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[1] ),
        .Q(\u0/uk/K_r5 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[20] ),
        .Q(\u0/uk/K_r5 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[21] ),
        .Q(\u0/uk/K_r5 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[22] ),
        .Q(\u0/uk/K_r5 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[23] ),
        .Q(\u0/uk/K_r5 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[24] ),
        .Q(\u0/uk/K_r5 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[25] ),
        .Q(\u0/uk/K_r5 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[26] ),
        .Q(\u0/uk/K_r5 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[27] ),
        .Q(\u0/uk/K_r5 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[28] ),
        .Q(\u0/uk/K_r5 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[29] ),
        .Q(\u0/uk/K_r5 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[2] ),
        .Q(\u0/uk/K_r5 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[30] ),
        .Q(\u0/uk/K_r5 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[31] ),
        .Q(\u0/uk/K_r5 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[32] ),
        .Q(\u0/uk/K_r5 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[33] ),
        .Q(\u0/uk/K_r5 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_50_in ),
        .Q(\u0/uk/K_r5 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[35] ),
        .Q(\u0/uk/K_r5 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[36] ),
        .Q(\u0/uk/K_r5 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[37] ),
        .Q(\u0/uk/K_r5 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[38] ),
        .Q(\u0/uk/K_r5 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[39] ),
        .Q(\u0/uk/K_r5 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[3] ),
        .Q(\u0/uk/K_r5 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_49_in ),
        .Q(\u0/uk/K_r5 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[41] ),
        .Q(\u0/uk/K_r5 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[42] ),
        .Q(\u0/uk/K_r5 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_44_in ),
        .Q(\u0/uk/K_r5 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[44] ),
        .Q(\u0/uk/K_r5 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[45] ),
        .Q(\u0/uk/K_r5 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_47_in ),
        .Q(\u0/uk/K_r5 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[47] ),
        .Q(\u0/uk/K_r5 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[48] ),
        .Q(\u0/uk/K_r5 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[49] ),
        .Q(\u0/uk/K_r5 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[4] ),
        .Q(\u0/uk/K_r5 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[50] ),
        .Q(\u0/uk/K_r5 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[51] ),
        .Q(\u0/uk/K_r5 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[52] ),
        .Q(\u0/uk/K_r5 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_51_in ),
        .Q(\u0/uk/K_r5 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[54] ),
        .Q(\u0/uk/K_r5 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[55] ),
        .Q(\u0/uk/K_r5 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[5] ),
        .Q(\u0/uk/K_r5 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[6] ),
        .Q(\u0/uk/K_r5 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[7] ),
        .Q(\u0/uk/K_r5 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_42_in ),
        .Q(\u0/uk/K_r5 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r5_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r4_reg_n_0_[9] ),
        .Q(\u0/uk/K_r5 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [0]),
        .Q(\u0/uk/K_r6_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [10]),
        .Q(\u0/uk/K_r6_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [11]),
        .Q(\u0/uk/K_r6_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [12]),
        .Q(\u0/uk/K_r6_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [13]),
        .Q(\u0/uk/p_52_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [14]),
        .Q(\u0/uk/K_r6_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [15]),
        .Q(\u0/uk/K_r6_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [16]),
        .Q(\u0/uk/K_r6_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [17]),
        .Q(\u0/uk/K_r6_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [18]),
        .Q(\u0/uk/K_r6_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [19]),
        .Q(\u0/uk/K_r6_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [1]),
        .Q(\u0/uk/K_r6_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [20]),
        .Q(\u0/uk/K_r6_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [21]),
        .Q(\u0/uk/K_r6_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [22]),
        .Q(\u0/uk/K_r6_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [23]),
        .Q(\u0/uk/K_r6_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [24]),
        .Q(\u0/uk/K_r6_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [25]),
        .Q(\u0/uk/K_r6_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [26]),
        .Q(\u0/uk/K_r6_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [27]),
        .Q(\u0/uk/K_r6_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [28]),
        .Q(\u0/uk/K_r6_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [29]),
        .Q(\u0/uk/K_r6_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [2]),
        .Q(\u0/uk/K_r6_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [30]),
        .Q(\u0/uk/K_r6_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [31]),
        .Q(\u0/uk/K_r6_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [32]),
        .Q(\u0/uk/K_r6_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [33]),
        .Q(\u0/uk/K_r6_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [34]),
        .Q(\u0/uk/K_r6_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [35]),
        .Q(\u0/uk/K_r6_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [36]),
        .Q(\u0/uk/K_r6_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [37]),
        .Q(\u0/uk/K_r6_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [38]),
        .Q(\u0/uk/K_r6_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [39]),
        .Q(\u0/uk/K_r6_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [3]),
        .Q(\u0/uk/K_r6_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [40]),
        .Q(\u0/uk/K_r6_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [41]),
        .Q(\u0/uk/K_r6_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [42]),
        .Q(\u0/uk/p_41_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [43]),
        .Q(\u0/uk/p_45_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [44]),
        .Q(\u0/uk/K_r6_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [45]),
        .Q(\u0/uk/K_r6_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [46]),
        .Q(\u0/uk/K_r6_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [47]),
        .Q(\u0/uk/K_r6_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [48]),
        .Q(\u0/uk/K_r6_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [49]),
        .Q(\u0/uk/p_43_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [4]),
        .Q(\u0/uk/K_r6_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [50]),
        .Q(\u0/uk/K_r6_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [51]),
        .Q(\u0/uk/K_r6_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [52]),
        .Q(\u0/uk/K_r6_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [53]),
        .Q(\u0/uk/K_r6_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [54]),
        .Q(\u0/uk/K_r6_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [55]),
        .Q(\u0/uk/K_r6_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [5]),
        .Q(\u0/uk/K_r6_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [6]),
        .Q(\u0/uk/p_53_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [7]),
        .Q(\u0/uk/K_r6_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [8]),
        .Q(\u0/uk/K_r6_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r6_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r5 [9]),
        .Q(\u0/uk/K_r6_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_ ),
        .Q(\u0/uk/K_r7_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[10] ),
        .Q(\u0/uk/K_r7_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[11] ),
        .Q(\u0/uk/K_r7_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[12] ),
        .Q(\u0/uk/K_r7_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_52_in ),
        .Q(\u0/uk/K_r7_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[14] ),
        .Q(\u0/uk/K_r7_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[15] ),
        .Q(\u0/uk/K_r7_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[16] ),
        .Q(\u0/uk/K_r7_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[17] ),
        .Q(\u0/uk/K_r7_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[18] ),
        .Q(\u0/uk/K_r7_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[19] ),
        .Q(\u0/uk/K_r7_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[1] ),
        .Q(\u0/uk/K_r7_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[20] ),
        .Q(\u0/uk/K_r7_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[21] ),
        .Q(\u0/uk/K_r7_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[22] ),
        .Q(\u0/uk/K_r7_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[23] ),
        .Q(\u0/uk/K_r7_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[24] ),
        .Q(\u0/uk/K_r7_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[25] ),
        .Q(\u0/uk/K_r7_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[26] ),
        .Q(\u0/uk/K_r7_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[27] ),
        .Q(\u0/uk/K_r7_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[28] ),
        .Q(\u0/uk/K_r7_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[29] ),
        .Q(\u0/uk/K_r7_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[2] ),
        .Q(\u0/uk/K_r7_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[30] ),
        .Q(\u0/uk/K_r7_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[31] ),
        .Q(\u0/uk/K_r7_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[32] ),
        .Q(\u0/uk/K_r7_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[33] ),
        .Q(\u0/uk/K_r7_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[34] ),
        .Q(\u0/uk/K_r7_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[35] ),
        .Q(\u0/uk/K_r7_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[36] ),
        .Q(\u0/uk/K_r7_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[37] ),
        .Q(\u0/uk/K_r7_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[38] ),
        .Q(\u0/uk/K_r7_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[39] ),
        .Q(\u0/uk/K_r7_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[3] ),
        .Q(\u0/uk/K_r7_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[40] ),
        .Q(\u0/uk/K_r7_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[41] ),
        .Q(\u0/uk/K_r7_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_41_in ),
        .Q(\u0/uk/K_r7_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_45_in ),
        .Q(\u0/uk/K_r7_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[44] ),
        .Q(\u0/uk/p_48_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[45] ),
        .Q(\u0/uk/K_r7_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[46] ),
        .Q(\u0/uk/K_r7_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[47] ),
        .Q(\u0/uk/K_r7_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[48] ),
        .Q(\u0/uk/K_r7_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_43_in ),
        .Q(\u0/uk/K_r7_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[4] ),
        .Q(\u0/uk/K_r7_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[50] ),
        .Q(\u0/uk/K_r7_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[51] ),
        .Q(\u0/uk/K_r7_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[52] ),
        .Q(\u0/uk/K_r7_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[53] ),
        .Q(\u0/uk/K_r7_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[54] ),
        .Q(\u0/uk/K_r7_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[55] ),
        .Q(\u0/uk/K_r7_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[5] ),
        .Q(\u0/uk/K_r7_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_53_in ),
        .Q(\u0/uk/K_r7_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[7] ),
        .Q(\u0/uk/K_r7_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[8] ),
        .Q(\u0/uk/K_r7_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r7_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r6_reg_n_0_[9] ),
        .Q(\u0/uk/K_r7_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_ ),
        .Q(\u0/uk/K_r8 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[10] ),
        .Q(\u0/uk/K_r8 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[11] ),
        .Q(\u0/uk/K_r8 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[12] ),
        .Q(\u0/uk/K_r8 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[13] ),
        .Q(\u0/uk/K_r8 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[14] ),
        .Q(\u0/uk/K_r8 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[15] ),
        .Q(\u0/uk/K_r8 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[16] ),
        .Q(\u0/uk/K_r8 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[17] ),
        .Q(\u0/uk/K_r8 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[18] ),
        .Q(\u0/uk/K_r8 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[19] ),
        .Q(\u0/uk/K_r8 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[1] ),
        .Q(\u0/uk/K_r8 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[20] ),
        .Q(\u0/uk/K_r8 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[21] ),
        .Q(\u0/uk/K_r8 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[22] ),
        .Q(\u0/uk/K_r8 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[23] ),
        .Q(\u0/uk/K_r8 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[24] ),
        .Q(\u0/uk/K_r8 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[25] ),
        .Q(\u0/uk/K_r8 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[26] ),
        .Q(\u0/uk/K_r8 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[27] ),
        .Q(\u0/uk/K_r8 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[28] ),
        .Q(\u0/uk/K_r8 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[29] ),
        .Q(\u0/uk/K_r8 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[2] ),
        .Q(\u0/uk/K_r8 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[30] ),
        .Q(\u0/uk/K_r8 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[31] ),
        .Q(\u0/uk/K_r8 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[32] ),
        .Q(\u0/uk/K_r8 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[33] ),
        .Q(\u0/uk/K_r8 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[34] ),
        .Q(\u0/uk/K_r8 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[35] ),
        .Q(\u0/uk/K_r8 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[36] ),
        .Q(\u0/uk/K_r8 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[37] ),
        .Q(\u0/uk/K_r8 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[38] ),
        .Q(\u0/uk/K_r8 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[39] ),
        .Q(\u0/uk/K_r8 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[3] ),
        .Q(\u0/uk/K_r8 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[40] ),
        .Q(\u0/uk/K_r8 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[41] ),
        .Q(\u0/uk/K_r8 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[42] ),
        .Q(\u0/uk/K_r8 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[43] ),
        .Q(\u0/uk/K_r8 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/p_48_in ),
        .Q(\u0/uk/K_r8 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[45] ),
        .Q(\u0/uk/K_r8 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[46] ),
        .Q(\u0/uk/K_r8 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[47] ),
        .Q(\u0/uk/K_r8 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[48] ),
        .Q(\u0/uk/K_r8 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[49] ),
        .Q(\u0/uk/K_r8 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[4] ),
        .Q(\u0/uk/K_r8 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[50] ),
        .Q(\u0/uk/K_r8 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[51] ),
        .Q(\u0/uk/K_r8 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[52] ),
        .Q(\u0/uk/K_r8 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[53] ),
        .Q(\u0/uk/K_r8 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[54] ),
        .Q(\u0/uk/K_r8 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[55] ),
        .Q(\u0/uk/K_r8 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[5] ),
        .Q(\u0/uk/K_r8 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[6] ),
        .Q(\u0/uk/K_r8 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[7] ),
        .Q(\u0/uk/K_r8 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[8] ),
        .Q(\u0/uk/K_r8 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r8_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r7_reg_n_0_[9] ),
        .Q(\u0/uk/K_r8 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [0]),
        .Q(\u0/uk/K_r9 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [10]),
        .Q(\u0/uk/K_r9 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [11]),
        .Q(\u0/uk/K_r9 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [12]),
        .Q(\u0/uk/K_r9 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [13]),
        .Q(\u0/uk/K_r9 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [14]),
        .Q(\u0/uk/K_r9 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [15]),
        .Q(\u0/uk/K_r9 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [16]),
        .Q(\u0/uk/K_r9 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [17]),
        .Q(\u0/uk/K_r9 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [18]),
        .Q(\u0/uk/K_r9 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [19]),
        .Q(\u0/uk/K_r9 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [1]),
        .Q(\u0/uk/K_r9 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [20]),
        .Q(\u0/uk/K_r9 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [21]),
        .Q(\u0/uk/K_r9 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [22]),
        .Q(\u0/uk/K_r9 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [23]),
        .Q(\u0/uk/K_r9 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [24]),
        .Q(\u0/uk/K_r9 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [25]),
        .Q(\u0/uk/K_r9 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [26]),
        .Q(\u0/uk/K_r9 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [27]),
        .Q(\u0/uk/K_r9 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [28]),
        .Q(\u0/uk/K_r9 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [29]),
        .Q(\u0/uk/K_r9 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [2]),
        .Q(\u0/uk/K_r9 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [30]),
        .Q(\u0/uk/K_r9 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [31]),
        .Q(\u0/uk/K_r9 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [32]),
        .Q(\u0/uk/K_r9 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [33]),
        .Q(\u0/uk/K_r9 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [34]),
        .Q(\u0/uk/K_r9 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [35]),
        .Q(\u0/uk/K_r9 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [36]),
        .Q(\u0/uk/K_r9 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [37]),
        .Q(\u0/uk/K_r9 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [38]),
        .Q(\u0/uk/K_r9 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [39]),
        .Q(\u0/uk/K_r9 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [3]),
        .Q(\u0/uk/K_r9 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [40]),
        .Q(\u0/uk/K_r9 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [41]),
        .Q(\u0/uk/K_r9 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [42]),
        .Q(\u0/uk/K_r9 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [43]),
        .Q(\u0/uk/K_r9 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [44]),
        .Q(\u0/uk/K_r9 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [45]),
        .Q(\u0/uk/K_r9 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [46]),
        .Q(\u0/uk/K_r9 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [47]),
        .Q(\u0/uk/K_r9 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [48]),
        .Q(\u0/uk/K_r9 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [49]),
        .Q(\u0/uk/K_r9 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [4]),
        .Q(\u0/uk/K_r9 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [50]),
        .Q(\u0/uk/K_r9 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [51]),
        .Q(\u0/uk/K_r9 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [52]),
        .Q(\u0/uk/K_r9 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [53]),
        .Q(\u0/uk/K_r9 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [54]),
        .Q(\u0/uk/K_r9 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [55]),
        .Q(\u0/uk/K_r9 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [5]),
        .Q(\u0/uk/K_r9 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [6]),
        .Q(\u0/uk/K_r9 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [7]),
        .Q(\u0/uk/K_r9 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [8]),
        .Q(\u0/uk/K_r9 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u0/uk/K_r9_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u0/uk/K_r8 [9]),
        .Q(\u0/uk/K_r9 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [42]),
        .Q(\u1/L0 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [43]),
        .Q(\u1/L0 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [44]),
        .Q(\u1/L0 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [45]),
        .Q(\u1/L0 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [46]),
        .Q(\u1/L0 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [47]),
        .Q(\u1/L0 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [48]),
        .Q(\u1/L0 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [49]),
        .Q(\u1/L0 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [50]),
        .Q(\u1/L0 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [51]),
        .Q(\u1/L0 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [33]),
        .Q(\u1/L0 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [52]),
        .Q(\u1/L0 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [53]),
        .Q(\u1/L0 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [54]),
        .Q(\u1/L0 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [55]),
        .Q(\u1/L0 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [56]),
        .Q(\u1/L0 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [57]),
        .Q(\u1/L0 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [58]),
        .Q(\u1/L0 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [59]),
        .Q(\u1/L0 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [60]),
        .Q(\u1/L0 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [61]),
        .Q(\u1/L0 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [34]),
        .Q(\u1/L0 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [62]),
        .Q(\u1/L0 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [63]),
        .Q(\u1/L0 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [64]),
        .Q(\u1/L0 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [35]),
        .Q(\u1/L0 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [36]),
        .Q(\u1/L0 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [37]),
        .Q(\u1/L0 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [38]),
        .Q(\u1/L0 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [39]),
        .Q(\u1/L0 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [40]),
        .Q(\u1/L0 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L0_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/IP [41]),
        .Q(\u1/L0 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [10]),
        .Q(\u1/L10 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [11]),
        .Q(\u1/L10 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [12]),
        .Q(\u1/L10 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [13]),
        .Q(\u1/L10 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [14]),
        .Q(\u1/L10 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [15]),
        .Q(\u1/L10 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [16]),
        .Q(\u1/L10 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [17]),
        .Q(\u1/L10 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [18]),
        .Q(\u1/L10 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [19]),
        .Q(\u1/L10 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [1]),
        .Q(\u1/L10 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [20]),
        .Q(\u1/L10 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [21]),
        .Q(\u1/L10 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [22]),
        .Q(\u1/L10 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [23]),
        .Q(\u1/L10 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [24]),
        .Q(\u1/L10 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [25]),
        .Q(\u1/L10 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [26]),
        .Q(\u1/L10 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [27]),
        .Q(\u1/L10 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [28]),
        .Q(\u1/L10 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [29]),
        .Q(\u1/L10 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [2]),
        .Q(\u1/L10 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [30]),
        .Q(\u1/L10 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [31]),
        .Q(\u1/L10 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [32]),
        .Q(\u1/L10 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [3]),
        .Q(\u1/L10 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [4]),
        .Q(\u1/L10 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [5]),
        .Q(\u1/L10 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [6]),
        .Q(\u1/L10 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [7]),
        .Q(\u1/L10 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [8]),
        .Q(\u1/L10 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L10_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R9 [9]),
        .Q(\u1/L10 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_ ),
        .Q(\u1/L11 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[11] ),
        .Q(\u1/L11 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[12] ),
        .Q(\u1/L11 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[13] ),
        .Q(\u1/L11 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[14] ),
        .Q(\u1/L11 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[15] ),
        .Q(\u1/L11 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[16] ),
        .Q(\u1/L11 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[17] ),
        .Q(\u1/L11 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[18] ),
        .Q(\u1/L11 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[19] ),
        .Q(\u1/L11 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[1] ),
        .Q(\u1/L11 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[20] ),
        .Q(\u1/L11 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[21] ),
        .Q(\u1/L11 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[22] ),
        .Q(\u1/L11 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[23] ),
        .Q(\u1/L11 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[24] ),
        .Q(\u1/L11 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[25] ),
        .Q(\u1/L11 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[26] ),
        .Q(\u1/L11 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[27] ),
        .Q(\u1/L11 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[28] ),
        .Q(\u1/L11 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[29] ),
        .Q(\u1/L11 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[2] ),
        .Q(\u1/L11 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[30] ),
        .Q(\u1/L11 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[31] ),
        .Q(\u1/L11 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[32] ),
        .Q(\u1/L11 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[3] ),
        .Q(\u1/L11 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[4] ),
        .Q(\u1/L11 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[5] ),
        .Q(\u1/L11 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[6] ),
        .Q(\u1/L11 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[7] ),
        .Q(\u1/L11 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[8] ),
        .Q(\u1/L11 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L11_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10_reg_n_0_[9] ),
        .Q(\u1/L11 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [10]),
        .Q(\u1/L12 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [11]),
        .Q(\u1/L12 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [12]),
        .Q(\u1/L12 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [13]),
        .Q(\u1/L12 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [14]),
        .Q(\u1/L12 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [15]),
        .Q(\u1/L12 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [16]),
        .Q(\u1/L12 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [17]),
        .Q(\u1/L12 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [18]),
        .Q(\u1/L12 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [19]),
        .Q(\u1/L12 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [1]),
        .Q(\u1/L12 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [20]),
        .Q(\u1/L12 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [21]),
        .Q(\u1/L12 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [22]),
        .Q(\u1/L12 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [23]),
        .Q(\u1/L12 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [24]),
        .Q(\u1/L12 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [25]),
        .Q(\u1/L12 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [26]),
        .Q(\u1/L12 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [27]),
        .Q(\u1/L12 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [28]),
        .Q(\u1/L12 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [29]),
        .Q(\u1/L12 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [2]),
        .Q(\u1/L12 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [30]),
        .Q(\u1/L12 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [31]),
        .Q(\u1/L12 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [32]),
        .Q(\u1/L12 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [3]),
        .Q(\u1/L12 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [4]),
        .Q(\u1/L12 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [5]),
        .Q(\u1/L12 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [6]),
        .Q(\u1/L12 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [7]),
        .Q(\u1/L12 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [8]),
        .Q(\u1/L12 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L12_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R11 [9]),
        .Q(\u1/L12 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [10]),
        .Q(\u1/L13 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [11]),
        .Q(\u1/L13 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [12]),
        .Q(\u1/L13 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [13]),
        .Q(\u1/L13 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [14]),
        .Q(\u1/L13 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [15]),
        .Q(\u1/L13 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [16]),
        .Q(\u1/L13 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [17]),
        .Q(\u1/L13 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [18]),
        .Q(\u1/L13 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [19]),
        .Q(\u1/L13 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [1]),
        .Q(\u1/L13 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [20]),
        .Q(\u1/L13 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [21]),
        .Q(\u1/L13 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [22]),
        .Q(\u1/L13 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [23]),
        .Q(\u1/L13 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [24]),
        .Q(\u1/L13 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [25]),
        .Q(\u1/L13 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [26]),
        .Q(\u1/L13 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [27]),
        .Q(\u1/L13 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [28]),
        .Q(\u1/L13 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [29]),
        .Q(\u1/L13 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [2]),
        .Q(\u1/L13 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [30]),
        .Q(\u1/L13 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [31]),
        .Q(\u1/L13 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [32]),
        .Q(\u1/L13 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [3]),
        .Q(\u1/L13 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [4]),
        .Q(\u1/L13 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [5]),
        .Q(\u1/L13 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [6]),
        .Q(\u1/L13 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [7]),
        .Q(\u1/L13 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [8]),
        .Q(\u1/L13 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L13_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R12 [9]),
        .Q(\u1/L13 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [10]),
        .Q(\u1/L14 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [11]),
        .Q(\u1/L14 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [12]),
        .Q(\u1/L14 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [13]),
        .Q(\u1/L14 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [14]),
        .Q(\u1/L14 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [15]),
        .Q(\u1/L14 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [16]),
        .Q(\u1/L14 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [17]),
        .Q(\u1/L14 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [18]),
        .Q(\u1/L14 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [19]),
        .Q(\u1/L14 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [1]),
        .Q(\u1/L14 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [20]),
        .Q(\u1/L14 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [21]),
        .Q(\u1/L14 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [22]),
        .Q(\u1/L14 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [23]),
        .Q(\u1/L14 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [24]),
        .Q(\u1/L14 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [25]),
        .Q(\u1/L14 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [26]),
        .Q(\u1/L14 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [27]),
        .Q(\u1/L14 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [28]),
        .Q(\u1/L14 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [29]),
        .Q(\u1/L14 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [2]),
        .Q(\u1/L14 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [30]),
        .Q(\u1/L14 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [31]),
        .Q(\u1/L14 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [32]),
        .Q(\u1/L14 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [3]),
        .Q(\u1/L14 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [4]),
        .Q(\u1/L14 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [5]),
        .Q(\u1/L14 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [6]),
        .Q(\u1/L14 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [7]),
        .Q(\u1/L14 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [8]),
        .Q(\u1/L14 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L14_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R13 [9]),
        .Q(\u1/L14 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [10]),
        .Q(\u1/L1 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [11]),
        .Q(\u1/L1 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [12]),
        .Q(\u1/L1 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [13]),
        .Q(\u1/L1 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [14]),
        .Q(\u1/L1 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [15]),
        .Q(\u1/L1 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [16]),
        .Q(\u1/L1 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [17]),
        .Q(\u1/L1 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [18]),
        .Q(\u1/L1 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [19]),
        .Q(\u1/L1 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [1]),
        .Q(\u1/L1 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [20]),
        .Q(\u1/L1 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [21]),
        .Q(\u1/L1 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [22]),
        .Q(\u1/L1 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [23]),
        .Q(\u1/L1 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [24]),
        .Q(\u1/L1 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [25]),
        .Q(\u1/L1 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [26]),
        .Q(\u1/L1 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [27]),
        .Q(\u1/L1 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [28]),
        .Q(\u1/L1 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [29]),
        .Q(\u1/L1 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [2]),
        .Q(\u1/L1 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [30]),
        .Q(\u1/L1 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [31]),
        .Q(\u1/L1 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [32]),
        .Q(\u1/L1 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [3]),
        .Q(\u1/L1 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [4]),
        .Q(\u1/L1 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [5]),
        .Q(\u1/L1 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [6]),
        .Q(\u1/L1 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [7]),
        .Q(\u1/L1 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [8]),
        .Q(\u1/L1 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R0 [9]),
        .Q(\u1/L1 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [10]),
        .Q(\u1/L2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [11]),
        .Q(\u1/L2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [12]),
        .Q(\u1/L2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [13]),
        .Q(\u1/L2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [14]),
        .Q(\u1/L2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [15]),
        .Q(\u1/L2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [16]),
        .Q(\u1/L2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [17]),
        .Q(\u1/L2 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [18]),
        .Q(\u1/L2 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [19]),
        .Q(\u1/L2 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [1]),
        .Q(\u1/L2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [20]),
        .Q(\u1/L2 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [21]),
        .Q(\u1/L2 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [22]),
        .Q(\u1/L2 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [23]),
        .Q(\u1/L2 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [24]),
        .Q(\u1/L2 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [25]),
        .Q(\u1/L2 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [26]),
        .Q(\u1/L2 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [27]),
        .Q(\u1/L2 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [28]),
        .Q(\u1/L2 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [29]),
        .Q(\u1/L2 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [2]),
        .Q(\u1/L2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [30]),
        .Q(\u1/L2 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [31]),
        .Q(\u1/L2 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [32]),
        .Q(\u1/L2 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [3]),
        .Q(\u1/L2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [4]),
        .Q(\u1/L2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [5]),
        .Q(\u1/L2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [6]),
        .Q(\u1/L2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [7]),
        .Q(\u1/L2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [8]),
        .Q(\u1/L2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L2_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R1 [9]),
        .Q(\u1/L2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [10]),
        .Q(\u1/L3 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [11]),
        .Q(\u1/L3 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [12]),
        .Q(\u1/L3 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [13]),
        .Q(\u1/L3 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [14]),
        .Q(\u1/L3 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [15]),
        .Q(\u1/L3 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [16]),
        .Q(\u1/L3 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [17]),
        .Q(\u1/L3 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [18]),
        .Q(\u1/L3 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [19]),
        .Q(\u1/L3 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [1]),
        .Q(\u1/L3 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [20]),
        .Q(\u1/L3 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [21]),
        .Q(\u1/L3 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [22]),
        .Q(\u1/L3 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [23]),
        .Q(\u1/L3 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [24]),
        .Q(\u1/L3 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [25]),
        .Q(\u1/L3 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [26]),
        .Q(\u1/L3 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [27]),
        .Q(\u1/L3 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [28]),
        .Q(\u1/L3 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [29]),
        .Q(\u1/L3 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [2]),
        .Q(\u1/L3 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [30]),
        .Q(\u1/L3 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [31]),
        .Q(\u1/L3 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [32]),
        .Q(\u1/L3 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [3]),
        .Q(\u1/L3 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [4]),
        .Q(\u1/L3 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [5]),
        .Q(\u1/L3 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [6]),
        .Q(\u1/L3 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [7]),
        .Q(\u1/L3 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [8]),
        .Q(\u1/L3 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L3_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R2 [9]),
        .Q(\u1/L3 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [10]),
        .Q(\u1/L4 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [11]),
        .Q(\u1/L4 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [12]),
        .Q(\u1/L4 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [13]),
        .Q(\u1/L4 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [14]),
        .Q(\u1/L4 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [15]),
        .Q(\u1/L4 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [16]),
        .Q(\u1/L4 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [17]),
        .Q(\u1/L4 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [18]),
        .Q(\u1/L4 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [19]),
        .Q(\u1/L4 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [1]),
        .Q(\u1/L4 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [20]),
        .Q(\u1/L4 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [21]),
        .Q(\u1/L4 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [22]),
        .Q(\u1/L4 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [23]),
        .Q(\u1/L4 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [24]),
        .Q(\u1/L4 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [25]),
        .Q(\u1/L4 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [26]),
        .Q(\u1/L4 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [27]),
        .Q(\u1/L4 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [28]),
        .Q(\u1/L4 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [29]),
        .Q(\u1/L4 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [2]),
        .Q(\u1/L4 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [30]),
        .Q(\u1/L4 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [31]),
        .Q(\u1/L4 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [32]),
        .Q(\u1/L4 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [3]),
        .Q(\u1/L4 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [4]),
        .Q(\u1/L4 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [5]),
        .Q(\u1/L4 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [6]),
        .Q(\u1/L4 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [7]),
        .Q(\u1/L4 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [8]),
        .Q(\u1/L4 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L4_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R3 [9]),
        .Q(\u1/L4 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [10]),
        .Q(\u1/L5 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [11]),
        .Q(\u1/L5 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [12]),
        .Q(\u1/L5 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [13]),
        .Q(\u1/L5 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [14]),
        .Q(\u1/L5 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [15]),
        .Q(\u1/L5 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [16]),
        .Q(\u1/L5 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [17]),
        .Q(\u1/L5 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [18]),
        .Q(\u1/L5 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [19]),
        .Q(\u1/L5 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [1]),
        .Q(\u1/L5 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [20]),
        .Q(\u1/L5 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [21]),
        .Q(\u1/L5 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [22]),
        .Q(\u1/L5 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [23]),
        .Q(\u1/L5 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [24]),
        .Q(\u1/L5 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [25]),
        .Q(\u1/L5 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [26]),
        .Q(\u1/L5 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [27]),
        .Q(\u1/L5 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [28]),
        .Q(\u1/L5 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [29]),
        .Q(\u1/L5 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [2]),
        .Q(\u1/L5 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [30]),
        .Q(\u1/L5 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [31]),
        .Q(\u1/L5 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [32]),
        .Q(\u1/L5 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [3]),
        .Q(\u1/L5 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [4]),
        .Q(\u1/L5 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [5]),
        .Q(\u1/L5 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [6]),
        .Q(\u1/L5 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [7]),
        .Q(\u1/L5 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [8]),
        .Q(\u1/L5 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L5_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R4 [9]),
        .Q(\u1/L5 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [10]),
        .Q(\u1/L6 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [11]),
        .Q(\u1/L6 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [12]),
        .Q(\u1/L6 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [13]),
        .Q(\u1/L6 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [14]),
        .Q(\u1/L6 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [15]),
        .Q(\u1/L6 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [16]),
        .Q(\u1/L6 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [17]),
        .Q(\u1/L6 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [18]),
        .Q(\u1/L6 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [19]),
        .Q(\u1/L6 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [1]),
        .Q(\u1/L6 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [20]),
        .Q(\u1/L6 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [21]),
        .Q(\u1/L6 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [22]),
        .Q(\u1/L6 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [23]),
        .Q(\u1/L6 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [24]),
        .Q(\u1/L6 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [25]),
        .Q(\u1/L6 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [26]),
        .Q(\u1/L6 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [27]),
        .Q(\u1/L6 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [28]),
        .Q(\u1/L6 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [29]),
        .Q(\u1/L6 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [2]),
        .Q(\u1/L6 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [30]),
        .Q(\u1/L6 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [31]),
        .Q(\u1/L6 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [32]),
        .Q(\u1/L6 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [3]),
        .Q(\u1/L6 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [4]),
        .Q(\u1/L6 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [5]),
        .Q(\u1/L6 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [6]),
        .Q(\u1/L6 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [7]),
        .Q(\u1/L6 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [8]),
        .Q(\u1/L6 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L6_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R5 [9]),
        .Q(\u1/L6 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [10]),
        .Q(\u1/L7 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [11]),
        .Q(\u1/L7 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [12]),
        .Q(\u1/L7 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [13]),
        .Q(\u1/L7 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [14]),
        .Q(\u1/L7 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [15]),
        .Q(\u1/L7 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [16]),
        .Q(\u1/L7 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [17]),
        .Q(\u1/L7 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [18]),
        .Q(\u1/L7 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [19]),
        .Q(\u1/L7 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [1]),
        .Q(\u1/L7 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [20]),
        .Q(\u1/L7 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [21]),
        .Q(\u1/L7 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [22]),
        .Q(\u1/L7 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [23]),
        .Q(\u1/L7 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [24]),
        .Q(\u1/L7 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [25]),
        .Q(\u1/L7 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [26]),
        .Q(\u1/L7 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [27]),
        .Q(\u1/L7 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [28]),
        .Q(\u1/L7 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [29]),
        .Q(\u1/L7 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [2]),
        .Q(\u1/L7 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [30]),
        .Q(\u1/L7 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [31]),
        .Q(\u1/L7 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [32]),
        .Q(\u1/L7 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [3]),
        .Q(\u1/L7 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [4]),
        .Q(\u1/L7 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [5]),
        .Q(\u1/L7 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [6]),
        .Q(\u1/L7 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [7]),
        .Q(\u1/L7 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [8]),
        .Q(\u1/L7 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L7_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R6 [9]),
        .Q(\u1/L7 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [10]),
        .Q(\u1/L8 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [11]),
        .Q(\u1/L8 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [12]),
        .Q(\u1/L8 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [13]),
        .Q(\u1/L8 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [14]),
        .Q(\u1/L8 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [15]),
        .Q(\u1/L8 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [16]),
        .Q(\u1/L8 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [17]),
        .Q(\u1/L8 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [18]),
        .Q(\u1/L8 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [19]),
        .Q(\u1/L8 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [1]),
        .Q(\u1/L8 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [20]),
        .Q(\u1/L8 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [21]),
        .Q(\u1/L8 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [22]),
        .Q(\u1/L8 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [23]),
        .Q(\u1/L8 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [24]),
        .Q(\u1/L8 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [25]),
        .Q(\u1/L8 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [26]),
        .Q(\u1/L8 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [27]),
        .Q(\u1/L8 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [28]),
        .Q(\u1/L8 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [29]),
        .Q(\u1/L8 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [2]),
        .Q(\u1/L8 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [30]),
        .Q(\u1/L8 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [31]),
        .Q(\u1/L8 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [32]),
        .Q(\u1/L8 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [3]),
        .Q(\u1/L8 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [4]),
        .Q(\u1/L8 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [5]),
        .Q(\u1/L8 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [6]),
        .Q(\u1/L8 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [7]),
        .Q(\u1/L8 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [8]),
        .Q(\u1/L8 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L8_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R7 [9]),
        .Q(\u1/L8 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [10]),
        .Q(\u1/L9 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [11]),
        .Q(\u1/L9 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [12]),
        .Q(\u1/L9 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [13]),
        .Q(\u1/L9 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [14]),
        .Q(\u1/L9 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [15]),
        .Q(\u1/L9 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [16]),
        .Q(\u1/L9 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [17]),
        .Q(\u1/L9 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [18]),
        .Q(\u1/L9 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [19]),
        .Q(\u1/L9 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [1]),
        .Q(\u1/L9 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [20]),
        .Q(\u1/L9 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [21]),
        .Q(\u1/L9 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [22]),
        .Q(\u1/L9 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [23]),
        .Q(\u1/L9 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [24]),
        .Q(\u1/L9 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [25]),
        .Q(\u1/L9 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [26]),
        .Q(\u1/L9 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [27]),
        .Q(\u1/L9 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [28]),
        .Q(\u1/L9 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [29]),
        .Q(\u1/L9 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [2]),
        .Q(\u1/L9 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [30]),
        .Q(\u1/L9 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [31]),
        .Q(\u1/L9 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [32]),
        .Q(\u1/L9 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [3]),
        .Q(\u1/L9 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [4]),
        .Q(\u1/L9 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [5]),
        .Q(\u1/L9 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [6]),
        .Q(\u1/L9 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [7]),
        .Q(\u1/L9 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [8]),
        .Q(\u1/L9 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/L9_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R8 [9]),
        .Q(\u1/L9 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[10]_i_1 
       (.I0(\u1/IP [10]),
        .I1(\u1/out0 [10]),
        .O(\u1/R00 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[11]_i_1 
       (.I0(\u1/IP [11]),
        .I1(\u1/out0 [11]),
        .O(\u1/R00 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[12]_i_1 
       (.I0(\u1/IP [12]),
        .I1(\u1/out0 [12]),
        .O(\u1/R00 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[13]_i_1 
       (.I0(\u1/IP [13]),
        .I1(\u1/out0 [13]),
        .O(\u1/R00 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[14]_i_1 
       (.I0(\u1/IP [14]),
        .I1(\u1/out0 [14]),
        .O(\u1/R00 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[15]_i_1 
       (.I0(\u1/IP [15]),
        .I1(\u1/out0 [15]),
        .O(\u1/R00 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[16]_i_1 
       (.I0(\u1/IP [16]),
        .I1(\u1/out0 [16]),
        .O(\u1/R00 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[17]_i_1 
       (.I0(\u1/IP [17]),
        .I1(\u1/out0 [17]),
        .O(\u1/R00 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[18]_i_1 
       (.I0(\u1/IP [18]),
        .I1(\u1/out0 [18]),
        .O(\u1/R00 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[19]_i_1 
       (.I0(\u1/IP [19]),
        .I1(\u1/out0 [19]),
        .O(\u1/R00 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[1]_i_1 
       (.I0(\u1/IP [1]),
        .I1(\u1/out0 [1]),
        .O(\u1/R00 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[20]_i_1 
       (.I0(\u1/IP [20]),
        .I1(\u1/out0 [20]),
        .O(\u1/R00 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[21]_i_1 
       (.I0(\u1/IP [21]),
        .I1(\u1/out0 [21]),
        .O(\u1/R00 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[22]_i_1 
       (.I0(\u1/IP [22]),
        .I1(\u1/out0 [22]),
        .O(\u1/R00 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[23]_i_1 
       (.I0(\u1/IP [23]),
        .I1(\u1/out0 [23]),
        .O(\u1/R00 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[24]_i_1 
       (.I0(\u1/IP [24]),
        .I1(\u1/out0 [24]),
        .O(\u1/R00 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[25]_i_1 
       (.I0(\u1/IP [25]),
        .I1(\u1/out0 [25]),
        .O(\u1/R00 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[26]_i_1 
       (.I0(\u1/IP [26]),
        .I1(\u1/out0 [26]),
        .O(\u1/R00 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[27]_i_1 
       (.I0(\u1/IP [27]),
        .I1(\u1/out0 [27]),
        .O(\u1/R00 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[28]_i_1 
       (.I0(\u1/IP [28]),
        .I1(\u1/out0 [28]),
        .O(\u1/R00 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[29]_i_1 
       (.I0(\u1/IP [29]),
        .I1(\u1/out0 [29]),
        .O(\u1/R00 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[2]_i_1 
       (.I0(\u1/IP [2]),
        .I1(\u1/out0 [2]),
        .O(\u1/R00 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[30]_i_1 
       (.I0(\u1/IP [30]),
        .I1(\u1/out0 [30]),
        .O(\u1/R00 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[31]_i_1 
       (.I0(\u1/IP [31]),
        .I1(\u1/out0 [31]),
        .O(\u1/R00 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[32]_i_1 
       (.I0(\u1/IP [32]),
        .I1(\u1/out0 [32]),
        .O(\u1/R00 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[3]_i_1 
       (.I0(\u1/IP [3]),
        .I1(\u1/out0 [3]),
        .O(\u1/R00 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[4]_i_1 
       (.I0(\u1/IP [4]),
        .I1(\u1/out0 [4]),
        .O(\u1/R00 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[5]_i_1 
       (.I0(\u1/IP [5]),
        .I1(\u1/out0 [5]),
        .O(\u1/R00 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[6]_i_1 
       (.I0(\u1/IP [6]),
        .I1(\u1/out0 [6]),
        .O(\u1/R00 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[7]_i_1 
       (.I0(\u1/IP [7]),
        .I1(\u1/out0 [7]),
        .O(\u1/R00 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[8]_i_1 
       (.I0(\u1/IP [8]),
        .I1(\u1/out0 [8]),
        .O(\u1/R00 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R0[9]_i_1 
       (.I0(\u1/IP [9]),
        .I1(\u1/out0 [9]),
        .O(\u1/R00 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [22]),
        .Q(\u1/R0 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [21]),
        .Q(\u1/R0 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [20]),
        .Q(\u1/R0 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [19]),
        .Q(\u1/R0 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [18]),
        .Q(\u1/R0 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [17]),
        .Q(\u1/R0 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [16]),
        .Q(\u1/R0 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [15]),
        .Q(\u1/R0 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [14]),
        .Q(\u1/R0 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [13]),
        .Q(\u1/R0 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [31]),
        .Q(\u1/R0 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [12]),
        .Q(\u1/R0 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [11]),
        .Q(\u1/R0 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [10]),
        .Q(\u1/R0 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [9]),
        .Q(\u1/R0 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [8]),
        .Q(\u1/R0 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [7]),
        .Q(\u1/R0 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [6]),
        .Q(\u1/R0 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [5]),
        .Q(\u1/R0 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [4]),
        .Q(\u1/R0 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [3]),
        .Q(\u1/R0 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [30]),
        .Q(\u1/R0 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [2]),
        .Q(\u1/R0 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [1]),
        .Q(\u1/R0 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [0]),
        .Q(\u1/R0 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [29]),
        .Q(\u1/R0 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [28]),
        .Q(\u1/R0 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [27]),
        .Q(\u1/R0 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [26]),
        .Q(\u1/R0 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [25]),
        .Q(\u1/R0 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [24]),
        .Q(\u1/R0 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R0_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R00 [23]),
        .Q(\u1/R0 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[10]_i_1 
       (.I0(\u1/L9 [10]),
        .I1(\u1/out10 [10]),
        .O(\u1/R100 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[11]_i_1 
       (.I0(\u1/L9 [11]),
        .I1(\u1/out10 [11]),
        .O(\u1/R100 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[12]_i_1 
       (.I0(\u1/L9 [12]),
        .I1(\u1/out10 [12]),
        .O(\u1/R100 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[13]_i_1 
       (.I0(\u1/L9 [13]),
        .I1(\u1/out10 [13]),
        .O(\u1/R100 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[14]_i_1 
       (.I0(\u1/L9 [14]),
        .I1(\u1/out10 [14]),
        .O(\u1/R100 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[15]_i_1 
       (.I0(\u1/L9 [15]),
        .I1(\u1/out10 [15]),
        .O(\u1/R100 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[16]_i_1 
       (.I0(\u1/L9 [16]),
        .I1(\u1/out10 [16]),
        .O(\u1/R100 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[17]_i_1 
       (.I0(\u1/L9 [17]),
        .I1(\u1/out10 [17]),
        .O(\u1/R100 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[18]_i_1 
       (.I0(\u1/L9 [18]),
        .I1(\u1/out10 [18]),
        .O(\u1/R100 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[19]_i_1 
       (.I0(\u1/L9 [19]),
        .I1(\u1/out10 [19]),
        .O(\u1/R100 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[1]_i_1 
       (.I0(\u1/L9 [1]),
        .I1(\u1/out10 [1]),
        .O(\u1/R100 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[20]_i_1 
       (.I0(\u1/L9 [20]),
        .I1(\u1/out10 [20]),
        .O(\u1/R100 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[21]_i_1 
       (.I0(\u1/L9 [21]),
        .I1(\u1/out10 [21]),
        .O(\u1/R100 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[22]_i_1 
       (.I0(\u1/L9 [22]),
        .I1(\u1/out10 [22]),
        .O(\u1/R100 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[23]_i_1 
       (.I0(\u1/L9 [23]),
        .I1(\u1/out10 [23]),
        .O(\u1/R100 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[24]_i_1 
       (.I0(\u1/L9 [24]),
        .I1(\u1/out10 [24]),
        .O(\u1/R100 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[25]_i_1 
       (.I0(\u1/L9 [25]),
        .I1(\u1/out10 [25]),
        .O(\u1/R100 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[26]_i_1 
       (.I0(\u1/L9 [26]),
        .I1(\u1/out10 [26]),
        .O(\u1/R100 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[27]_i_1 
       (.I0(\u1/L9 [27]),
        .I1(\u1/out10 [27]),
        .O(\u1/R100 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[28]_i_1 
       (.I0(\u1/L9 [28]),
        .I1(\u1/out10 [28]),
        .O(\u1/R100 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[29]_i_1 
       (.I0(\u1/L9 [29]),
        .I1(\u1/out10 [29]),
        .O(\u1/R100 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[2]_i_1 
       (.I0(\u1/L9 [2]),
        .I1(\u1/out10 [2]),
        .O(\u1/R100 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[30]_i_1 
       (.I0(\u1/L9 [30]),
        .I1(\u1/out10 [30]),
        .O(\u1/R100 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[31]_i_1 
       (.I0(\u1/L9 [31]),
        .I1(\u1/out10 [31]),
        .O(\u1/R100 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[32]_i_1 
       (.I0(\u1/L9 [32]),
        .I1(\u1/out10 [32]),
        .O(\u1/R100 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[3]_i_1 
       (.I0(\u1/L9 [3]),
        .I1(\u1/out10 [3]),
        .O(\u1/R100 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[4]_i_1 
       (.I0(\u1/L9 [4]),
        .I1(\u1/out10 [4]),
        .O(\u1/R100 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[5]_i_1 
       (.I0(\u1/L9 [5]),
        .I1(\u1/out10 [5]),
        .O(\u1/R100 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[6]_i_1 
       (.I0(\u1/L9 [6]),
        .I1(\u1/out10 [6]),
        .O(\u1/R100 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[7]_i_1 
       (.I0(\u1/L9 [7]),
        .I1(\u1/out10 [7]),
        .O(\u1/R100 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[8]_i_1 
       (.I0(\u1/L9 [8]),
        .I1(\u1/out10 [8]),
        .O(\u1/R100 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R10[9]_i_1 
       (.I0(\u1/L9 [9]),
        .I1(\u1/out10 [9]),
        .O(\u1/R100 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [22]),
        .Q(\u1/R10_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [21]),
        .Q(\u1/R10_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [20]),
        .Q(\u1/R10_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [19]),
        .Q(\u1/R10_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [18]),
        .Q(\u1/R10_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [17]),
        .Q(\u1/R10_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [16]),
        .Q(\u1/R10_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [15]),
        .Q(\u1/R10_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [14]),
        .Q(\u1/R10_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [13]),
        .Q(\u1/R10_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [31]),
        .Q(\u1/R10_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [12]),
        .Q(\u1/R10_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [11]),
        .Q(\u1/R10_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [10]),
        .Q(\u1/R10_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [9]),
        .Q(\u1/R10_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [8]),
        .Q(\u1/R10_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [7]),
        .Q(\u1/R10_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [6]),
        .Q(\u1/R10_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [5]),
        .Q(\u1/R10_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [4]),
        .Q(\u1/R10_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [3]),
        .Q(\u1/R10_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [30]),
        .Q(\u1/R10_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [2]),
        .Q(\u1/R10_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [1]),
        .Q(\u1/R10_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [0]),
        .Q(\u1/R10_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [29]),
        .Q(\u1/R10_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [28]),
        .Q(\u1/R10_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [27]),
        .Q(\u1/R10_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [26]),
        .Q(\u1/R10_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [25]),
        .Q(\u1/R10_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [24]),
        .Q(\u1/R10_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R10_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R100 [23]),
        .Q(\u1/R10_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[10]_i_1 
       (.I0(\u1/L10 [10]),
        .I1(\u1/out11 [10]),
        .O(\u1/R110 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[11]_i_1 
       (.I0(\u1/L10 [11]),
        .I1(\u1/out11 [11]),
        .O(\u1/R110 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[12]_i_1 
       (.I0(\u1/L10 [12]),
        .I1(\u1/out11 [12]),
        .O(\u1/R110 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[13]_i_1 
       (.I0(\u1/L10 [13]),
        .I1(\u1/out11 [13]),
        .O(\u1/R110 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[14]_i_1 
       (.I0(\u1/L10 [14]),
        .I1(\u1/out11 [14]),
        .O(\u1/R110 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[15]_i_1 
       (.I0(\u1/L10 [15]),
        .I1(\u1/out11 [15]),
        .O(\u1/R110 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[16]_i_1 
       (.I0(\u1/L10 [16]),
        .I1(\u1/out11 [16]),
        .O(\u1/R110 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[17]_i_1 
       (.I0(\u1/L10 [17]),
        .I1(\u1/out11 [17]),
        .O(\u1/R110 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[18]_i_1 
       (.I0(\u1/L10 [18]),
        .I1(\u1/out11 [18]),
        .O(\u1/R110 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[19]_i_1 
       (.I0(\u1/L10 [19]),
        .I1(\u1/out11 [19]),
        .O(\u1/R110 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[1]_i_1 
       (.I0(\u1/L10 [1]),
        .I1(\u1/out11 [1]),
        .O(\u1/R110 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[20]_i_1 
       (.I0(\u1/L10 [20]),
        .I1(\u1/out11 [20]),
        .O(\u1/R110 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[21]_i_1 
       (.I0(\u1/L10 [21]),
        .I1(\u1/out11 [21]),
        .O(\u1/R110 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[22]_i_1 
       (.I0(\u1/L10 [22]),
        .I1(\u1/out11 [22]),
        .O(\u1/R110 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[23]_i_1 
       (.I0(\u1/L10 [23]),
        .I1(\u1/out11 [23]),
        .O(\u1/R110 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[24]_i_1 
       (.I0(\u1/L10 [24]),
        .I1(\u1/out11 [24]),
        .O(\u1/R110 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[25]_i_1 
       (.I0(\u1/L10 [25]),
        .I1(\u1/out11 [25]),
        .O(\u1/R110 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[26]_i_1 
       (.I0(\u1/L10 [26]),
        .I1(\u1/out11 [26]),
        .O(\u1/R110 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[27]_i_1 
       (.I0(\u1/L10 [27]),
        .I1(\u1/out11 [27]),
        .O(\u1/R110 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[28]_i_1 
       (.I0(\u1/L10 [28]),
        .I1(\u1/out11 [28]),
        .O(\u1/R110 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[29]_i_1 
       (.I0(\u1/L10 [29]),
        .I1(\u1/out11 [29]),
        .O(\u1/R110 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[2]_i_1 
       (.I0(\u1/L10 [2]),
        .I1(\u1/out11 [2]),
        .O(\u1/R110 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[30]_i_1 
       (.I0(\u1/L10 [30]),
        .I1(\u1/out11 [30]),
        .O(\u1/R110 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[31]_i_1 
       (.I0(\u1/L10 [31]),
        .I1(\u1/out11 [31]),
        .O(\u1/R110 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[32]_i_1 
       (.I0(\u1/L10 [32]),
        .I1(\u1/out11 [32]),
        .O(\u1/R110 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[3]_i_1 
       (.I0(\u1/L10 [3]),
        .I1(\u1/out11 [3]),
        .O(\u1/R110 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[4]_i_1 
       (.I0(\u1/L10 [4]),
        .I1(\u1/out11 [4]),
        .O(\u1/R110 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[5]_i_1 
       (.I0(\u1/L10 [5]),
        .I1(\u1/out11 [5]),
        .O(\u1/R110 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[6]_i_1 
       (.I0(\u1/L10 [6]),
        .I1(\u1/out11 [6]),
        .O(\u1/R110 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[7]_i_1 
       (.I0(\u1/L10 [7]),
        .I1(\u1/out11 [7]),
        .O(\u1/R110 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[8]_i_1 
       (.I0(\u1/L10 [8]),
        .I1(\u1/out11 [8]),
        .O(\u1/R110 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R11[9]_i_1 
       (.I0(\u1/L10 [9]),
        .I1(\u1/out11 [9]),
        .O(\u1/R110 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [22]),
        .Q(\u1/R11 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [21]),
        .Q(\u1/R11 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [20]),
        .Q(\u1/R11 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [19]),
        .Q(\u1/R11 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [18]),
        .Q(\u1/R11 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [17]),
        .Q(\u1/R11 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [16]),
        .Q(\u1/R11 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [15]),
        .Q(\u1/R11 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [14]),
        .Q(\u1/R11 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [13]),
        .Q(\u1/R11 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [31]),
        .Q(\u1/R11 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [12]),
        .Q(\u1/R11 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [11]),
        .Q(\u1/R11 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [10]),
        .Q(\u1/R11 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [9]),
        .Q(\u1/R11 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [8]),
        .Q(\u1/R11 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [7]),
        .Q(\u1/R11 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [6]),
        .Q(\u1/R11 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [5]),
        .Q(\u1/R11 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [4]),
        .Q(\u1/R11 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [3]),
        .Q(\u1/R11 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [30]),
        .Q(\u1/R11 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [2]),
        .Q(\u1/R11 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [1]),
        .Q(\u1/R11 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [0]),
        .Q(\u1/R11 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [29]),
        .Q(\u1/R11 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [28]),
        .Q(\u1/R11 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [27]),
        .Q(\u1/R11 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [26]),
        .Q(\u1/R11 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [25]),
        .Q(\u1/R11 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [24]),
        .Q(\u1/R11 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R11_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R110 [23]),
        .Q(\u1/R11 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[10]_i_1 
       (.I0(\u1/L11 [10]),
        .I1(\u1/out12 [10]),
        .O(\u1/R120 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[11]_i_1 
       (.I0(\u1/L11 [11]),
        .I1(\u1/out12 [11]),
        .O(\u1/R120 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[12]_i_1 
       (.I0(\u1/L11 [12]),
        .I1(\u1/out12 [12]),
        .O(\u1/R120 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[13]_i_1 
       (.I0(\u1/L11 [13]),
        .I1(\u1/out12 [13]),
        .O(\u1/R120 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[14]_i_1 
       (.I0(\u1/L11 [14]),
        .I1(\u1/out12 [14]),
        .O(\u1/R120 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[15]_i_1 
       (.I0(\u1/L11 [15]),
        .I1(\u1/out12 [15]),
        .O(\u1/R120 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[16]_i_1 
       (.I0(\u1/L11 [16]),
        .I1(\u1/out12 [16]),
        .O(\u1/R120 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[17]_i_1 
       (.I0(\u1/L11 [17]),
        .I1(\u1/out12 [17]),
        .O(\u1/R120 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[18]_i_1 
       (.I0(\u1/L11 [18]),
        .I1(\u1/out12 [18]),
        .O(\u1/R120 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[19]_i_1 
       (.I0(\u1/L11 [19]),
        .I1(\u1/out12 [19]),
        .O(\u1/R120 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[1]_i_1 
       (.I0(\u1/L11 [1]),
        .I1(\u1/out12 [1]),
        .O(\u1/R120 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[20]_i_1 
       (.I0(\u1/L11 [20]),
        .I1(\u1/out12 [20]),
        .O(\u1/R120 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[21]_i_1 
       (.I0(\u1/L11 [21]),
        .I1(\u1/out12 [21]),
        .O(\u1/R120 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[22]_i_1 
       (.I0(\u1/L11 [22]),
        .I1(\u1/out12 [22]),
        .O(\u1/R120 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[23]_i_1 
       (.I0(\u1/L11 [23]),
        .I1(\u1/out12 [23]),
        .O(\u1/R120 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[24]_i_1 
       (.I0(\u1/L11 [24]),
        .I1(\u1/out12 [24]),
        .O(\u1/R120 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[25]_i_1 
       (.I0(\u1/L11 [25]),
        .I1(\u1/out12 [25]),
        .O(\u1/R120 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[26]_i_1 
       (.I0(\u1/L11 [26]),
        .I1(\u1/out12 [26]),
        .O(\u1/R120 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[27]_i_1 
       (.I0(\u1/L11 [27]),
        .I1(\u1/out12 [27]),
        .O(\u1/R120 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[28]_i_1 
       (.I0(\u1/L11 [28]),
        .I1(\u1/out12 [28]),
        .O(\u1/R120 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[29]_i_1 
       (.I0(\u1/L11 [29]),
        .I1(\u1/out12 [29]),
        .O(\u1/R120 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[2]_i_1 
       (.I0(\u1/L11 [2]),
        .I1(\u1/out12 [2]),
        .O(\u1/R120 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[30]_i_1 
       (.I0(\u1/L11 [30]),
        .I1(\u1/out12 [30]),
        .O(\u1/R120 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[31]_i_1 
       (.I0(\u1/L11 [31]),
        .I1(\u1/out12 [31]),
        .O(\u1/R120 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[32]_i_1 
       (.I0(\u1/L11 [32]),
        .I1(\u1/out12 [32]),
        .O(\u1/R120 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[3]_i_1 
       (.I0(\u1/L11 [3]),
        .I1(\u1/out12 [3]),
        .O(\u1/R120 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[4]_i_1 
       (.I0(\u1/L11 [4]),
        .I1(\u1/out12 [4]),
        .O(\u1/R120 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[5]_i_1 
       (.I0(\u1/L11 [5]),
        .I1(\u1/out12 [5]),
        .O(\u1/R120 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[6]_i_1 
       (.I0(\u1/L11 [6]),
        .I1(\u1/out12 [6]),
        .O(\u1/R120 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[7]_i_1 
       (.I0(\u1/L11 [7]),
        .I1(\u1/out12 [7]),
        .O(\u1/R120 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[8]_i_1 
       (.I0(\u1/L11 [8]),
        .I1(\u1/out12 [8]),
        .O(\u1/R120 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R12[9]_i_1 
       (.I0(\u1/L11 [9]),
        .I1(\u1/out12 [9]),
        .O(\u1/R120 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [22]),
        .Q(\u1/R12 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [21]),
        .Q(\u1/R12 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [20]),
        .Q(\u1/R12 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [19]),
        .Q(\u1/R12 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [18]),
        .Q(\u1/R12 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [17]),
        .Q(\u1/R12 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [16]),
        .Q(\u1/R12 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [15]),
        .Q(\u1/R12 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [14]),
        .Q(\u1/R12 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [13]),
        .Q(\u1/R12 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [31]),
        .Q(\u1/R12 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [12]),
        .Q(\u1/R12 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [11]),
        .Q(\u1/R12 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [10]),
        .Q(\u1/R12 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [9]),
        .Q(\u1/R12 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [8]),
        .Q(\u1/R12 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [7]),
        .Q(\u1/R12 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [6]),
        .Q(\u1/R12 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [5]),
        .Q(\u1/R12 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [4]),
        .Q(\u1/R12 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [3]),
        .Q(\u1/R12 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [30]),
        .Q(\u1/R12 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [2]),
        .Q(\u1/R12 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [1]),
        .Q(\u1/R12 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [0]),
        .Q(\u1/R12 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [29]),
        .Q(\u1/R12 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [28]),
        .Q(\u1/R12 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [27]),
        .Q(\u1/R12 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [26]),
        .Q(\u1/R12 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [25]),
        .Q(\u1/R12 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [24]),
        .Q(\u1/R12 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R12_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R120 [23]),
        .Q(\u1/R12 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[10]_i_1 
       (.I0(\u1/L12 [10]),
        .I1(\u1/out13 [10]),
        .O(\u1/R130 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[11]_i_1 
       (.I0(\u1/L12 [11]),
        .I1(\u1/out13 [11]),
        .O(\u1/R130 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[12]_i_1 
       (.I0(\u1/L12 [12]),
        .I1(\u1/out13 [12]),
        .O(\u1/R130 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[13]_i_1 
       (.I0(\u1/L12 [13]),
        .I1(\u1/out13 [13]),
        .O(\u1/R130 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[14]_i_1 
       (.I0(\u1/L12 [14]),
        .I1(\u1/out13 [14]),
        .O(\u1/R130 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[15]_i_1 
       (.I0(\u1/L12 [15]),
        .I1(\u1/out13 [15]),
        .O(\u1/R130 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[16]_i_1 
       (.I0(\u1/L12 [16]),
        .I1(\u1/out13 [16]),
        .O(\u1/R130 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[17]_i_1 
       (.I0(\u1/L12 [17]),
        .I1(\u1/out13 [17]),
        .O(\u1/R130 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[18]_i_1 
       (.I0(\u1/L12 [18]),
        .I1(\u1/out13 [18]),
        .O(\u1/R130 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[19]_i_1 
       (.I0(\u1/L12 [19]),
        .I1(\u1/out13 [19]),
        .O(\u1/R130 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[1]_i_1 
       (.I0(\u1/L12 [1]),
        .I1(\u1/out13 [1]),
        .O(\u1/R130 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[20]_i_1 
       (.I0(\u1/L12 [20]),
        .I1(\u1/out13 [20]),
        .O(\u1/R130 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[21]_i_1 
       (.I0(\u1/L12 [21]),
        .I1(\u1/out13 [21]),
        .O(\u1/R130 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[22]_i_1 
       (.I0(\u1/L12 [22]),
        .I1(\u1/out13 [22]),
        .O(\u1/R130 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[23]_i_1 
       (.I0(\u1/L12 [23]),
        .I1(\u1/out13 [23]),
        .O(\u1/R130 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[24]_i_1 
       (.I0(\u1/L12 [24]),
        .I1(\u1/out13 [24]),
        .O(\u1/R130 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[25]_i_1 
       (.I0(\u1/L12 [25]),
        .I1(\u1/out13 [25]),
        .O(\u1/R130 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[26]_i_1 
       (.I0(\u1/L12 [26]),
        .I1(\u1/out13 [26]),
        .O(\u1/R130 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[27]_i_1 
       (.I0(\u1/L12 [27]),
        .I1(\u1/out13 [27]),
        .O(\u1/R130 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[28]_i_1 
       (.I0(\u1/L12 [28]),
        .I1(\u1/out13 [28]),
        .O(\u1/R130 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[29]_i_1 
       (.I0(\u1/L12 [29]),
        .I1(\u1/out13 [29]),
        .O(\u1/R130 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[2]_i_1 
       (.I0(\u1/L12 [2]),
        .I1(\u1/out13 [2]),
        .O(\u1/R130 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[30]_i_1 
       (.I0(\u1/L12 [30]),
        .I1(\u1/out13 [30]),
        .O(\u1/R130 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[31]_i_1 
       (.I0(\u1/L12 [31]),
        .I1(\u1/out13 [31]),
        .O(\u1/R130 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[32]_i_1 
       (.I0(\u1/L12 [32]),
        .I1(\u1/out13 [32]),
        .O(\u1/R130 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[3]_i_1 
       (.I0(\u1/L12 [3]),
        .I1(\u1/out13 [3]),
        .O(\u1/R130 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[4]_i_1 
       (.I0(\u1/L12 [4]),
        .I1(\u1/out13 [4]),
        .O(\u1/R130 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[5]_i_1 
       (.I0(\u1/L12 [5]),
        .I1(\u1/out13 [5]),
        .O(\u1/R130 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[6]_i_1 
       (.I0(\u1/L12 [6]),
        .I1(\u1/out13 [6]),
        .O(\u1/R130 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[7]_i_1 
       (.I0(\u1/L12 [7]),
        .I1(\u1/out13 [7]),
        .O(\u1/R130 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[8]_i_1 
       (.I0(\u1/L12 [8]),
        .I1(\u1/out13 [8]),
        .O(\u1/R130 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R13[9]_i_1 
       (.I0(\u1/L12 [9]),
        .I1(\u1/out13 [9]),
        .O(\u1/R130 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [22]),
        .Q(\u1/R13 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [21]),
        .Q(\u1/R13 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [20]),
        .Q(\u1/R13 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [19]),
        .Q(\u1/R13 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [18]),
        .Q(\u1/R13 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [17]),
        .Q(\u1/R13 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [16]),
        .Q(\u1/R13 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [15]),
        .Q(\u1/R13 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [14]),
        .Q(\u1/R13 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [13]),
        .Q(\u1/R13 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [31]),
        .Q(\u1/R13 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [12]),
        .Q(\u1/R13 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [11]),
        .Q(\u1/R13 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [10]),
        .Q(\u1/R13 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [9]),
        .Q(\u1/R13 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [8]),
        .Q(\u1/R13 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [7]),
        .Q(\u1/R13 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [6]),
        .Q(\u1/R13 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [5]),
        .Q(\u1/R13 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [4]),
        .Q(\u1/R13 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [3]),
        .Q(\u1/R13 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [30]),
        .Q(\u1/R13 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [2]),
        .Q(\u1/R13 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [1]),
        .Q(\u1/R13 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [0]),
        .Q(\u1/R13 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [29]),
        .Q(\u1/R13 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [28]),
        .Q(\u1/R13 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [27]),
        .Q(\u1/R13 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [26]),
        .Q(\u1/R13 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [25]),
        .Q(\u1/R13 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [24]),
        .Q(\u1/R13 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R13_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R130 [23]),
        .Q(\u1/R13 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[10]_i_1 
       (.I0(\u1/L13 [10]),
        .I1(\u1/out14 [10]),
        .O(\u1/R140 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[11]_i_1 
       (.I0(\u1/L13 [11]),
        .I1(\u1/out14 [11]),
        .O(\u1/R140 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[12]_i_1 
       (.I0(\u1/L13 [12]),
        .I1(\u1/out14 [12]),
        .O(\u1/R140 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[13]_i_1 
       (.I0(\u1/L13 [13]),
        .I1(\u1/out14 [13]),
        .O(\u1/R140 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[14]_i_1 
       (.I0(\u1/L13 [14]),
        .I1(\u1/out14 [14]),
        .O(\u1/R140 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[15]_i_1 
       (.I0(\u1/L13 [15]),
        .I1(\u1/out14 [15]),
        .O(\u1/R140 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[16]_i_1 
       (.I0(\u1/L13 [16]),
        .I1(\u1/out14 [16]),
        .O(\u1/R140 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[17]_i_1 
       (.I0(\u1/L13 [17]),
        .I1(\u1/out14 [17]),
        .O(\u1/R140 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[18]_i_1 
       (.I0(\u1/L13 [18]),
        .I1(\u1/out14 [18]),
        .O(\u1/R140 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[19]_i_1 
       (.I0(\u1/L13 [19]),
        .I1(\u1/out14 [19]),
        .O(\u1/R140 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[1]_i_1 
       (.I0(\u1/L13 [1]),
        .I1(\u1/out14 [1]),
        .O(\u1/R140 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[20]_i_1 
       (.I0(\u1/L13 [20]),
        .I1(\u1/out14 [20]),
        .O(\u1/R140 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[21]_i_1 
       (.I0(\u1/L13 [21]),
        .I1(\u1/out14 [21]),
        .O(\u1/R140 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[22]_i_1 
       (.I0(\u1/L13 [22]),
        .I1(\u1/out14 [22]),
        .O(\u1/R140 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[23]_i_1 
       (.I0(\u1/L13 [23]),
        .I1(\u1/out14 [23]),
        .O(\u1/R140 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[24]_i_1 
       (.I0(\u1/L13 [24]),
        .I1(\u1/out14 [24]),
        .O(\u1/R140 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[25]_i_1 
       (.I0(\u1/L13 [25]),
        .I1(\u1/out14 [25]),
        .O(\u1/R140 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[26]_i_1 
       (.I0(\u1/L13 [26]),
        .I1(\u1/out14 [26]),
        .O(\u1/R140 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[27]_i_1 
       (.I0(\u1/L13 [27]),
        .I1(\u1/out14 [27]),
        .O(\u1/R140 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[28]_i_1 
       (.I0(\u1/L13 [28]),
        .I1(\u1/out14 [28]),
        .O(\u1/R140 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[29]_i_1 
       (.I0(\u1/L13 [29]),
        .I1(\u1/out14 [29]),
        .O(\u1/R140 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[2]_i_1 
       (.I0(\u1/L13 [2]),
        .I1(\u1/out14 [2]),
        .O(\u1/R140 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[30]_i_1 
       (.I0(\u1/L13 [30]),
        .I1(\u1/out14 [30]),
        .O(\u1/R140 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[31]_i_1 
       (.I0(\u1/L13 [31]),
        .I1(\u1/out14 [31]),
        .O(\u1/R140 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[32]_i_1 
       (.I0(\u1/L13 [32]),
        .I1(\u1/out14 [32]),
        .O(\u1/R140 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[3]_i_1 
       (.I0(\u1/L13 [3]),
        .I1(\u1/out14 [3]),
        .O(\u1/R140 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[4]_i_1 
       (.I0(\u1/L13 [4]),
        .I1(\u1/out14 [4]),
        .O(\u1/R140 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[5]_i_1 
       (.I0(\u1/L13 [5]),
        .I1(\u1/out14 [5]),
        .O(\u1/R140 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[6]_i_1 
       (.I0(\u1/L13 [6]),
        .I1(\u1/out14 [6]),
        .O(\u1/R140 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[7]_i_1 
       (.I0(\u1/L13 [7]),
        .I1(\u1/out14 [7]),
        .O(\u1/R140 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[8]_i_1 
       (.I0(\u1/L13 [8]),
        .I1(\u1/out14 [8]),
        .O(\u1/R140 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R14[9]_i_1 
       (.I0(\u1/L13 [9]),
        .I1(\u1/out14 [9]),
        .O(\u1/R140 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [22]),
        .Q(\u1/FP [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [21]),
        .Q(\u1/FP [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [20]),
        .Q(\u1/FP [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [19]),
        .Q(\u1/FP [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [18]),
        .Q(\u1/FP [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [17]),
        .Q(\u1/FP [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [16]),
        .Q(\u1/FP [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [15]),
        .Q(\u1/FP [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [14]),
        .Q(\u1/FP [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [13]),
        .Q(\u1/FP [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [31]),
        .Q(\u1/FP [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [12]),
        .Q(\u1/FP [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [11]),
        .Q(\u1/FP [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [10]),
        .Q(\u1/FP [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [9]),
        .Q(\u1/FP [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [8]),
        .Q(\u1/FP [56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [7]),
        .Q(\u1/FP [57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [6]),
        .Q(\u1/FP [58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [5]),
        .Q(\u1/FP [59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [4]),
        .Q(\u1/FP [60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [3]),
        .Q(\u1/FP [61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [30]),
        .Q(\u1/FP [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [2]),
        .Q(\u1/FP [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [1]),
        .Q(\u1/FP [63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [0]),
        .Q(\u1/FP [64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [29]),
        .Q(\u1/FP [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [28]),
        .Q(\u1/FP [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [27]),
        .Q(\u1/FP [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [26]),
        .Q(\u1/FP [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [25]),
        .Q(\u1/FP [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [24]),
        .Q(\u1/FP [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R14_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R140 [23]),
        .Q(\u1/FP [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[10]_i_1 
       (.I0(\u1/L0 [10]),
        .I1(\u1/out1 [10]),
        .O(\u1/R10 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[11]_i_1 
       (.I0(\u1/L0 [11]),
        .I1(\u1/out1 [11]),
        .O(\u1/R10 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[12]_i_1 
       (.I0(\u1/L0 [12]),
        .I1(\u1/out1 [12]),
        .O(\u1/R10 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[13]_i_1 
       (.I0(\u1/L0 [13]),
        .I1(\u1/out1 [13]),
        .O(\u1/R10 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[14]_i_1 
       (.I0(\u1/L0 [14]),
        .I1(\u1/out1 [14]),
        .O(\u1/R10 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[15]_i_1 
       (.I0(\u1/L0 [15]),
        .I1(\u1/out1 [15]),
        .O(\u1/R10 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[16]_i_1 
       (.I0(\u1/L0 [16]),
        .I1(\u1/out1 [16]),
        .O(\u1/R10 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[17]_i_1 
       (.I0(\u1/L0 [17]),
        .I1(\u1/out1 [17]),
        .O(\u1/R10 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[18]_i_1 
       (.I0(\u1/L0 [18]),
        .I1(\u1/out1 [18]),
        .O(\u1/R10 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[19]_i_1 
       (.I0(\u1/L0 [19]),
        .I1(\u1/out1 [19]),
        .O(\u1/R10 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[1]_i_1 
       (.I0(\u1/L0 [1]),
        .I1(\u1/out1 [1]),
        .O(\u1/R10 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[20]_i_1 
       (.I0(\u1/L0 [20]),
        .I1(\u1/out1 [20]),
        .O(\u1/R10 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[21]_i_1 
       (.I0(\u1/L0 [21]),
        .I1(\u1/out1 [21]),
        .O(\u1/R10 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[22]_i_1 
       (.I0(\u1/L0 [22]),
        .I1(\u1/out1 [22]),
        .O(\u1/R10 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[23]_i_1 
       (.I0(\u1/L0 [23]),
        .I1(\u1/out1 [23]),
        .O(\u1/R10 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[24]_i_1 
       (.I0(\u1/L0 [24]),
        .I1(\u1/out1 [24]),
        .O(\u1/R10 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[25]_i_1 
       (.I0(\u1/L0 [25]),
        .I1(\u1/out1 [25]),
        .O(\u1/R10 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[26]_i_1 
       (.I0(\u1/L0 [26]),
        .I1(\u1/out1 [26]),
        .O(\u1/R10 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[27]_i_1 
       (.I0(\u1/L0 [27]),
        .I1(\u1/out1 [27]),
        .O(\u1/R10 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[28]_i_1 
       (.I0(\u1/L0 [28]),
        .I1(\u1/out1 [28]),
        .O(\u1/R10 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[29]_i_1 
       (.I0(\u1/L0 [29]),
        .I1(\u1/out1 [29]),
        .O(\u1/R10 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[2]_i_1 
       (.I0(\u1/L0 [2]),
        .I1(\u1/out1 [2]),
        .O(\u1/R10 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[30]_i_1 
       (.I0(\u1/L0 [30]),
        .I1(\u1/out1 [30]),
        .O(\u1/R10 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[31]_i_1 
       (.I0(\u1/L0 [31]),
        .I1(\u1/out1 [31]),
        .O(\u1/R10 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[32]_i_1 
       (.I0(\u1/L0 [32]),
        .I1(\u1/out1 [32]),
        .O(\u1/R10 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[3]_i_1 
       (.I0(\u1/L0 [3]),
        .I1(\u1/out1 [3]),
        .O(\u1/R10 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[4]_i_1 
       (.I0(\u1/L0 [4]),
        .I1(\u1/out1 [4]),
        .O(\u1/R10 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[5]_i_1 
       (.I0(\u1/L0 [5]),
        .I1(\u1/out1 [5]),
        .O(\u1/R10 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[6]_i_1 
       (.I0(\u1/L0 [6]),
        .I1(\u1/out1 [6]),
        .O(\u1/R10 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[7]_i_1 
       (.I0(\u1/L0 [7]),
        .I1(\u1/out1 [7]),
        .O(\u1/R10 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[8]_i_1 
       (.I0(\u1/L0 [8]),
        .I1(\u1/out1 [8]),
        .O(\u1/R10 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R1[9]_i_1 
       (.I0(\u1/L0 [9]),
        .I1(\u1/out1 [9]),
        .O(\u1/R10 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [22]),
        .Q(\u1/R1 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [21]),
        .Q(\u1/R1 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [20]),
        .Q(\u1/R1 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [19]),
        .Q(\u1/R1 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [18]),
        .Q(\u1/R1 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [17]),
        .Q(\u1/R1 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [16]),
        .Q(\u1/R1 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [15]),
        .Q(\u1/R1 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [14]),
        .Q(\u1/R1 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [13]),
        .Q(\u1/R1 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [31]),
        .Q(\u1/R1 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [12]),
        .Q(\u1/R1 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [11]),
        .Q(\u1/R1 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [10]),
        .Q(\u1/R1 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [9]),
        .Q(\u1/R1 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [8]),
        .Q(\u1/R1 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [7]),
        .Q(\u1/R1 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [6]),
        .Q(\u1/R1 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [5]),
        .Q(\u1/R1 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [4]),
        .Q(\u1/R1 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [3]),
        .Q(\u1/R1 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [30]),
        .Q(\u1/R1 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [2]),
        .Q(\u1/R1 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [1]),
        .Q(\u1/R1 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [0]),
        .Q(\u1/R1 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [29]),
        .Q(\u1/R1 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [28]),
        .Q(\u1/R1 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [27]),
        .Q(\u1/R1 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [26]),
        .Q(\u1/R1 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [25]),
        .Q(\u1/R1 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [24]),
        .Q(\u1/R1 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R10 [23]),
        .Q(\u1/R1 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[10]_i_1 
       (.I0(\u1/L1 [10]),
        .I1(\u1/out2 [10]),
        .O(\u1/R20 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[11]_i_1 
       (.I0(\u1/L1 [11]),
        .I1(\u1/out2 [11]),
        .O(\u1/R20 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[12]_i_1 
       (.I0(\u1/L1 [12]),
        .I1(\u1/out2 [12]),
        .O(\u1/R20 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[13]_i_1 
       (.I0(\u1/L1 [13]),
        .I1(\u1/out2 [13]),
        .O(\u1/R20 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[14]_i_1 
       (.I0(\u1/L1 [14]),
        .I1(\u1/out2 [14]),
        .O(\u1/R20 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[15]_i_1 
       (.I0(\u1/L1 [15]),
        .I1(\u1/out2 [15]),
        .O(\u1/R20 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[16]_i_1 
       (.I0(\u1/L1 [16]),
        .I1(\u1/out2 [16]),
        .O(\u1/R20 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[17]_i_1 
       (.I0(\u1/L1 [17]),
        .I1(\u1/out2 [17]),
        .O(\u1/R20 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[18]_i_1 
       (.I0(\u1/L1 [18]),
        .I1(\u1/out2 [18]),
        .O(\u1/R20 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[19]_i_1 
       (.I0(\u1/L1 [19]),
        .I1(\u1/out2 [19]),
        .O(\u1/R20 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[1]_i_1 
       (.I0(\u1/L1 [1]),
        .I1(\u1/out2 [1]),
        .O(\u1/R20 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[20]_i_1 
       (.I0(\u1/L1 [20]),
        .I1(\u1/out2 [20]),
        .O(\u1/R20 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[21]_i_1 
       (.I0(\u1/L1 [21]),
        .I1(\u1/out2 [21]),
        .O(\u1/R20 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[22]_i_1 
       (.I0(\u1/L1 [22]),
        .I1(\u1/out2 [22]),
        .O(\u1/R20 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[23]_i_1 
       (.I0(\u1/L1 [23]),
        .I1(\u1/out2 [23]),
        .O(\u1/R20 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[24]_i_1 
       (.I0(\u1/L1 [24]),
        .I1(\u1/out2 [24]),
        .O(\u1/R20 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[25]_i_1 
       (.I0(\u1/L1 [25]),
        .I1(\u1/out2 [25]),
        .O(\u1/R20 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[26]_i_1 
       (.I0(\u1/L1 [26]),
        .I1(\u1/out2 [26]),
        .O(\u1/R20 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[27]_i_1 
       (.I0(\u1/L1 [27]),
        .I1(\u1/out2 [27]),
        .O(\u1/R20 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[28]_i_1 
       (.I0(\u1/L1 [28]),
        .I1(\u1/out2 [28]),
        .O(\u1/R20 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[29]_i_1 
       (.I0(\u1/L1 [29]),
        .I1(\u1/out2 [29]),
        .O(\u1/R20 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[2]_i_1 
       (.I0(\u1/L1 [2]),
        .I1(\u1/out2 [2]),
        .O(\u1/R20 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[30]_i_1 
       (.I0(\u1/L1 [30]),
        .I1(\u1/out2 [30]),
        .O(\u1/R20 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[31]_i_1 
       (.I0(\u1/L1 [31]),
        .I1(\u1/out2 [31]),
        .O(\u1/R20 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[32]_i_1 
       (.I0(\u1/L1 [32]),
        .I1(\u1/out2 [32]),
        .O(\u1/R20 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[3]_i_1 
       (.I0(\u1/L1 [3]),
        .I1(\u1/out2 [3]),
        .O(\u1/R20 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[4]_i_1 
       (.I0(\u1/L1 [4]),
        .I1(\u1/out2 [4]),
        .O(\u1/R20 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[5]_i_1 
       (.I0(\u1/L1 [5]),
        .I1(\u1/out2 [5]),
        .O(\u1/R20 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[6]_i_1 
       (.I0(\u1/L1 [6]),
        .I1(\u1/out2 [6]),
        .O(\u1/R20 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[7]_i_1 
       (.I0(\u1/L1 [7]),
        .I1(\u1/out2 [7]),
        .O(\u1/R20 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[8]_i_1 
       (.I0(\u1/L1 [8]),
        .I1(\u1/out2 [8]),
        .O(\u1/R20 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R2[9]_i_1 
       (.I0(\u1/L1 [9]),
        .I1(\u1/out2 [9]),
        .O(\u1/R20 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [22]),
        .Q(\u1/R2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [21]),
        .Q(\u1/R2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [20]),
        .Q(\u1/R2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [19]),
        .Q(\u1/R2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [18]),
        .Q(\u1/R2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [17]),
        .Q(\u1/R2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [16]),
        .Q(\u1/R2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [15]),
        .Q(\u1/R2 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [14]),
        .Q(\u1/R2 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [13]),
        .Q(\u1/R2 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [31]),
        .Q(\u1/R2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [12]),
        .Q(\u1/R2 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [11]),
        .Q(\u1/R2 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [10]),
        .Q(\u1/R2 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [9]),
        .Q(\u1/R2 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [8]),
        .Q(\u1/R2 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [7]),
        .Q(\u1/R2 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [6]),
        .Q(\u1/R2 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [5]),
        .Q(\u1/R2 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [4]),
        .Q(\u1/R2 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [3]),
        .Q(\u1/R2 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [30]),
        .Q(\u1/R2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [2]),
        .Q(\u1/R2 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [1]),
        .Q(\u1/R2 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [0]),
        .Q(\u1/R2 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [29]),
        .Q(\u1/R2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [28]),
        .Q(\u1/R2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [27]),
        .Q(\u1/R2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [26]),
        .Q(\u1/R2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [25]),
        .Q(\u1/R2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [24]),
        .Q(\u1/R2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R2_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R20 [23]),
        .Q(\u1/R2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[10]_i_1 
       (.I0(\u1/L2 [10]),
        .I1(\u1/out3 [10]),
        .O(\u1/R30 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[11]_i_1 
       (.I0(\u1/L2 [11]),
        .I1(\u1/out3 [11]),
        .O(\u1/R30 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[12]_i_1 
       (.I0(\u1/L2 [12]),
        .I1(\u1/out3 [12]),
        .O(\u1/R30 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[13]_i_1 
       (.I0(\u1/L2 [13]),
        .I1(\u1/out3 [13]),
        .O(\u1/R30 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[14]_i_1 
       (.I0(\u1/L2 [14]),
        .I1(\u1/out3 [14]),
        .O(\u1/R30 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[15]_i_1 
       (.I0(\u1/L2 [15]),
        .I1(\u1/out3 [15]),
        .O(\u1/R30 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[16]_i_1 
       (.I0(\u1/L2 [16]),
        .I1(\u1/out3 [16]),
        .O(\u1/R30 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[17]_i_1 
       (.I0(\u1/L2 [17]),
        .I1(\u1/out3 [17]),
        .O(\u1/R30 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[18]_i_1 
       (.I0(\u1/L2 [18]),
        .I1(\u1/out3 [18]),
        .O(\u1/R30 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[19]_i_1 
       (.I0(\u1/L2 [19]),
        .I1(\u1/out3 [19]),
        .O(\u1/R30 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[1]_i_1 
       (.I0(\u1/L2 [1]),
        .I1(\u1/out3 [1]),
        .O(\u1/R30 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[20]_i_1 
       (.I0(\u1/L2 [20]),
        .I1(\u1/out3 [20]),
        .O(\u1/R30 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[21]_i_1 
       (.I0(\u1/L2 [21]),
        .I1(\u1/out3 [21]),
        .O(\u1/R30 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[22]_i_1 
       (.I0(\u1/L2 [22]),
        .I1(\u1/out3 [22]),
        .O(\u1/R30 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[23]_i_1 
       (.I0(\u1/L2 [23]),
        .I1(\u1/out3 [23]),
        .O(\u1/R30 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[24]_i_1 
       (.I0(\u1/L2 [24]),
        .I1(\u1/out3 [24]),
        .O(\u1/R30 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[25]_i_1 
       (.I0(\u1/L2 [25]),
        .I1(\u1/out3 [25]),
        .O(\u1/R30 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[26]_i_1 
       (.I0(\u1/L2 [26]),
        .I1(\u1/out3 [26]),
        .O(\u1/R30 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[27]_i_1 
       (.I0(\u1/L2 [27]),
        .I1(\u1/out3 [27]),
        .O(\u1/R30 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[28]_i_1 
       (.I0(\u1/L2 [28]),
        .I1(\u1/out3 [28]),
        .O(\u1/R30 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[29]_i_1 
       (.I0(\u1/L2 [29]),
        .I1(\u1/out3 [29]),
        .O(\u1/R30 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[2]_i_1 
       (.I0(\u1/L2 [2]),
        .I1(\u1/out3 [2]),
        .O(\u1/R30 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[30]_i_1 
       (.I0(\u1/L2 [30]),
        .I1(\u1/out3 [30]),
        .O(\u1/R30 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[31]_i_1 
       (.I0(\u1/L2 [31]),
        .I1(\u1/out3 [31]),
        .O(\u1/R30 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[32]_i_1 
       (.I0(\u1/L2 [32]),
        .I1(\u1/out3 [32]),
        .O(\u1/R30 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[3]_i_1 
       (.I0(\u1/L2 [3]),
        .I1(\u1/out3 [3]),
        .O(\u1/R30 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[4]_i_1 
       (.I0(\u1/L2 [4]),
        .I1(\u1/out3 [4]),
        .O(\u1/R30 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[5]_i_1 
       (.I0(\u1/L2 [5]),
        .I1(\u1/out3 [5]),
        .O(\u1/R30 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[6]_i_1 
       (.I0(\u1/L2 [6]),
        .I1(\u1/out3 [6]),
        .O(\u1/R30 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[7]_i_1 
       (.I0(\u1/L2 [7]),
        .I1(\u1/out3 [7]),
        .O(\u1/R30 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[8]_i_1 
       (.I0(\u1/L2 [8]),
        .I1(\u1/out3 [8]),
        .O(\u1/R30 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R3[9]_i_1 
       (.I0(\u1/L2 [9]),
        .I1(\u1/out3 [9]),
        .O(\u1/R30 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [22]),
        .Q(\u1/R3 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [21]),
        .Q(\u1/R3 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [20]),
        .Q(\u1/R3 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [19]),
        .Q(\u1/R3 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [18]),
        .Q(\u1/R3 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [17]),
        .Q(\u1/R3 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [16]),
        .Q(\u1/R3 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [15]),
        .Q(\u1/R3 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [14]),
        .Q(\u1/R3 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [13]),
        .Q(\u1/R3 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [31]),
        .Q(\u1/R3 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [12]),
        .Q(\u1/R3 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [11]),
        .Q(\u1/R3 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [10]),
        .Q(\u1/R3 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [9]),
        .Q(\u1/R3 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [8]),
        .Q(\u1/R3 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [7]),
        .Q(\u1/R3 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [6]),
        .Q(\u1/R3 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [5]),
        .Q(\u1/R3 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [4]),
        .Q(\u1/R3 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [3]),
        .Q(\u1/R3 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [30]),
        .Q(\u1/R3 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [2]),
        .Q(\u1/R3 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [1]),
        .Q(\u1/R3 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [0]),
        .Q(\u1/R3 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [29]),
        .Q(\u1/R3 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [28]),
        .Q(\u1/R3 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [27]),
        .Q(\u1/R3 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [26]),
        .Q(\u1/R3 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [25]),
        .Q(\u1/R3 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [24]),
        .Q(\u1/R3 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R3_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R30 [23]),
        .Q(\u1/R3 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[10]_i_1 
       (.I0(\u1/L3 [10]),
        .I1(\u1/out4 [10]),
        .O(\u1/R40 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[11]_i_1 
       (.I0(\u1/L3 [11]),
        .I1(\u1/out4 [11]),
        .O(\u1/R40 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[12]_i_1 
       (.I0(\u1/L3 [12]),
        .I1(\u1/out4 [12]),
        .O(\u1/R40 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[13]_i_1 
       (.I0(\u1/L3 [13]),
        .I1(\u1/out4 [13]),
        .O(\u1/R40 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[14]_i_1 
       (.I0(\u1/L3 [14]),
        .I1(\u1/out4 [14]),
        .O(\u1/R40 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[15]_i_1 
       (.I0(\u1/L3 [15]),
        .I1(\u1/out4 [15]),
        .O(\u1/R40 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[16]_i_1 
       (.I0(\u1/L3 [16]),
        .I1(\u1/out4 [16]),
        .O(\u1/R40 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[17]_i_1 
       (.I0(\u1/L3 [17]),
        .I1(\u1/out4 [17]),
        .O(\u1/R40 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[18]_i_1 
       (.I0(\u1/L3 [18]),
        .I1(\u1/out4 [18]),
        .O(\u1/R40 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[19]_i_1 
       (.I0(\u1/L3 [19]),
        .I1(\u1/out4 [19]),
        .O(\u1/R40 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[1]_i_1 
       (.I0(\u1/L3 [1]),
        .I1(\u1/out4 [1]),
        .O(\u1/R40 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[20]_i_1 
       (.I0(\u1/L3 [20]),
        .I1(\u1/out4 [20]),
        .O(\u1/R40 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[21]_i_1 
       (.I0(\u1/L3 [21]),
        .I1(\u1/out4 [21]),
        .O(\u1/R40 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[22]_i_1 
       (.I0(\u1/L3 [22]),
        .I1(\u1/out4 [22]),
        .O(\u1/R40 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[23]_i_1 
       (.I0(\u1/L3 [23]),
        .I1(\u1/out4 [23]),
        .O(\u1/R40 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[24]_i_1 
       (.I0(\u1/L3 [24]),
        .I1(\u1/out4 [24]),
        .O(\u1/R40 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[25]_i_1 
       (.I0(\u1/L3 [25]),
        .I1(\u1/out4 [25]),
        .O(\u1/R40 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[26]_i_1 
       (.I0(\u1/L3 [26]),
        .I1(\u1/out4 [26]),
        .O(\u1/R40 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[27]_i_1 
       (.I0(\u1/L3 [27]),
        .I1(\u1/out4 [27]),
        .O(\u1/R40 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[28]_i_1 
       (.I0(\u1/L3 [28]),
        .I1(\u1/out4 [28]),
        .O(\u1/R40 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[29]_i_1 
       (.I0(\u1/L3 [29]),
        .I1(\u1/out4 [29]),
        .O(\u1/R40 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[2]_i_1 
       (.I0(\u1/L3 [2]),
        .I1(\u1/out4 [2]),
        .O(\u1/R40 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[30]_i_1 
       (.I0(\u1/L3 [30]),
        .I1(\u1/out4 [30]),
        .O(\u1/R40 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[31]_i_1 
       (.I0(\u1/L3 [31]),
        .I1(\u1/out4 [31]),
        .O(\u1/R40 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[32]_i_1 
       (.I0(\u1/L3 [32]),
        .I1(\u1/out4 [32]),
        .O(\u1/R40 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[3]_i_1 
       (.I0(\u1/L3 [3]),
        .I1(\u1/out4 [3]),
        .O(\u1/R40 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[4]_i_1 
       (.I0(\u1/L3 [4]),
        .I1(\u1/out4 [4]),
        .O(\u1/R40 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[5]_i_1 
       (.I0(\u1/L3 [5]),
        .I1(\u1/out4 [5]),
        .O(\u1/R40 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[6]_i_1 
       (.I0(\u1/L3 [6]),
        .I1(\u1/out4 [6]),
        .O(\u1/R40 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[7]_i_1 
       (.I0(\u1/L3 [7]),
        .I1(\u1/out4 [7]),
        .O(\u1/R40 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[8]_i_1 
       (.I0(\u1/L3 [8]),
        .I1(\u1/out4 [8]),
        .O(\u1/R40 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R4[9]_i_1 
       (.I0(\u1/L3 [9]),
        .I1(\u1/out4 [9]),
        .O(\u1/R40 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [22]),
        .Q(\u1/R4 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [21]),
        .Q(\u1/R4 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [20]),
        .Q(\u1/R4 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [19]),
        .Q(\u1/R4 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [18]),
        .Q(\u1/R4 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [17]),
        .Q(\u1/R4 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [16]),
        .Q(\u1/R4 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [15]),
        .Q(\u1/R4 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [14]),
        .Q(\u1/R4 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [13]),
        .Q(\u1/R4 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [31]),
        .Q(\u1/R4 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [12]),
        .Q(\u1/R4 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [11]),
        .Q(\u1/R4 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [10]),
        .Q(\u1/R4 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [9]),
        .Q(\u1/R4 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [8]),
        .Q(\u1/R4 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [7]),
        .Q(\u1/R4 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [6]),
        .Q(\u1/R4 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [5]),
        .Q(\u1/R4 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [4]),
        .Q(\u1/R4 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [3]),
        .Q(\u1/R4 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [30]),
        .Q(\u1/R4 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [2]),
        .Q(\u1/R4 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [1]),
        .Q(\u1/R4 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [0]),
        .Q(\u1/R4 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [29]),
        .Q(\u1/R4 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [28]),
        .Q(\u1/R4 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [27]),
        .Q(\u1/R4 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [26]),
        .Q(\u1/R4 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [25]),
        .Q(\u1/R4 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [24]),
        .Q(\u1/R4 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R4_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R40 [23]),
        .Q(\u1/R4 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[10]_i_1 
       (.I0(\u1/L4 [10]),
        .I1(\u1/out5 [10]),
        .O(\u1/R50 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[11]_i_1 
       (.I0(\u1/L4 [11]),
        .I1(\u1/out5 [11]),
        .O(\u1/R50 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[12]_i_1 
       (.I0(\u1/L4 [12]),
        .I1(\u1/out5 [12]),
        .O(\u1/R50 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[13]_i_1 
       (.I0(\u1/L4 [13]),
        .I1(\u1/out5 [13]),
        .O(\u1/R50 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[14]_i_1 
       (.I0(\u1/L4 [14]),
        .I1(\u1/out5 [14]),
        .O(\u1/R50 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[15]_i_1 
       (.I0(\u1/L4 [15]),
        .I1(\u1/out5 [15]),
        .O(\u1/R50 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[16]_i_1 
       (.I0(\u1/L4 [16]),
        .I1(\u1/out5 [16]),
        .O(\u1/R50 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[17]_i_1 
       (.I0(\u1/L4 [17]),
        .I1(\u1/out5 [17]),
        .O(\u1/R50 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[18]_i_1 
       (.I0(\u1/L4 [18]),
        .I1(\u1/out5 [18]),
        .O(\u1/R50 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[19]_i_1 
       (.I0(\u1/L4 [19]),
        .I1(\u1/out5 [19]),
        .O(\u1/R50 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[1]_i_1 
       (.I0(\u1/L4 [1]),
        .I1(\u1/out5 [1]),
        .O(\u1/R50 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[20]_i_1 
       (.I0(\u1/L4 [20]),
        .I1(\u1/out5 [20]),
        .O(\u1/R50 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[21]_i_1 
       (.I0(\u1/L4 [21]),
        .I1(\u1/out5 [21]),
        .O(\u1/R50 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[22]_i_1 
       (.I0(\u1/L4 [22]),
        .I1(\u1/out5 [22]),
        .O(\u1/R50 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[23]_i_1 
       (.I0(\u1/L4 [23]),
        .I1(\u1/out5 [23]),
        .O(\u1/R50 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[24]_i_1 
       (.I0(\u1/L4 [24]),
        .I1(\u1/out5 [24]),
        .O(\u1/R50 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[25]_i_1 
       (.I0(\u1/L4 [25]),
        .I1(\u1/out5 [25]),
        .O(\u1/R50 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[26]_i_1 
       (.I0(\u1/L4 [26]),
        .I1(\u1/out5 [26]),
        .O(\u1/R50 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[27]_i_1 
       (.I0(\u1/L4 [27]),
        .I1(\u1/out5 [27]),
        .O(\u1/R50 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[28]_i_1 
       (.I0(\u1/L4 [28]),
        .I1(\u1/out5 [28]),
        .O(\u1/R50 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[29]_i_1 
       (.I0(\u1/L4 [29]),
        .I1(\u1/out5 [29]),
        .O(\u1/R50 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[2]_i_1 
       (.I0(\u1/L4 [2]),
        .I1(\u1/out5 [2]),
        .O(\u1/R50 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[30]_i_1 
       (.I0(\u1/L4 [30]),
        .I1(\u1/out5 [30]),
        .O(\u1/R50 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[31]_i_1 
       (.I0(\u1/L4 [31]),
        .I1(\u1/out5 [31]),
        .O(\u1/R50 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[32]_i_1 
       (.I0(\u1/L4 [32]),
        .I1(\u1/out5 [32]),
        .O(\u1/R50 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[3]_i_1 
       (.I0(\u1/L4 [3]),
        .I1(\u1/out5 [3]),
        .O(\u1/R50 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[4]_i_1 
       (.I0(\u1/L4 [4]),
        .I1(\u1/out5 [4]),
        .O(\u1/R50 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[5]_i_1 
       (.I0(\u1/L4 [5]),
        .I1(\u1/out5 [5]),
        .O(\u1/R50 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[6]_i_1 
       (.I0(\u1/L4 [6]),
        .I1(\u1/out5 [6]),
        .O(\u1/R50 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[7]_i_1 
       (.I0(\u1/L4 [7]),
        .I1(\u1/out5 [7]),
        .O(\u1/R50 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[8]_i_1 
       (.I0(\u1/L4 [8]),
        .I1(\u1/out5 [8]),
        .O(\u1/R50 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R5[9]_i_1 
       (.I0(\u1/L4 [9]),
        .I1(\u1/out5 [9]),
        .O(\u1/R50 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [22]),
        .Q(\u1/R5 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [21]),
        .Q(\u1/R5 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [20]),
        .Q(\u1/R5 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [19]),
        .Q(\u1/R5 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [18]),
        .Q(\u1/R5 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [17]),
        .Q(\u1/R5 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [16]),
        .Q(\u1/R5 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [15]),
        .Q(\u1/R5 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [14]),
        .Q(\u1/R5 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [13]),
        .Q(\u1/R5 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [31]),
        .Q(\u1/R5 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [12]),
        .Q(\u1/R5 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [11]),
        .Q(\u1/R5 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [10]),
        .Q(\u1/R5 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [9]),
        .Q(\u1/R5 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [8]),
        .Q(\u1/R5 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [7]),
        .Q(\u1/R5 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [6]),
        .Q(\u1/R5 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [5]),
        .Q(\u1/R5 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [4]),
        .Q(\u1/R5 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [3]),
        .Q(\u1/R5 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [30]),
        .Q(\u1/R5 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [2]),
        .Q(\u1/R5 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [1]),
        .Q(\u1/R5 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [0]),
        .Q(\u1/R5 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [29]),
        .Q(\u1/R5 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [28]),
        .Q(\u1/R5 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [27]),
        .Q(\u1/R5 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [26]),
        .Q(\u1/R5 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [25]),
        .Q(\u1/R5 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [24]),
        .Q(\u1/R5 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R5_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R50 [23]),
        .Q(\u1/R5 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[10]_i_1 
       (.I0(\u1/L5 [10]),
        .I1(\u1/out6 [10]),
        .O(\u1/R60 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[11]_i_1 
       (.I0(\u1/L5 [11]),
        .I1(\u1/out6 [11]),
        .O(\u1/R60 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[12]_i_1 
       (.I0(\u1/L5 [12]),
        .I1(\u1/out6 [12]),
        .O(\u1/R60 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[13]_i_1 
       (.I0(\u1/L5 [13]),
        .I1(\u1/out6 [13]),
        .O(\u1/R60 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[14]_i_1 
       (.I0(\u1/L5 [14]),
        .I1(\u1/out6 [14]),
        .O(\u1/R60 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[15]_i_1 
       (.I0(\u1/L5 [15]),
        .I1(\u1/out6 [15]),
        .O(\u1/R60 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[16]_i_1 
       (.I0(\u1/L5 [16]),
        .I1(\u1/out6 [16]),
        .O(\u1/R60 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[17]_i_1 
       (.I0(\u1/L5 [17]),
        .I1(\u1/out6 [17]),
        .O(\u1/R60 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[18]_i_1 
       (.I0(\u1/L5 [18]),
        .I1(\u1/out6 [18]),
        .O(\u1/R60 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[19]_i_1 
       (.I0(\u1/L5 [19]),
        .I1(\u1/out6 [19]),
        .O(\u1/R60 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[1]_i_1 
       (.I0(\u1/L5 [1]),
        .I1(\u1/out6 [1]),
        .O(\u1/R60 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[20]_i_1 
       (.I0(\u1/L5 [20]),
        .I1(\u1/out6 [20]),
        .O(\u1/R60 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[21]_i_1 
       (.I0(\u1/L5 [21]),
        .I1(\u1/out6 [21]),
        .O(\u1/R60 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[22]_i_1 
       (.I0(\u1/L5 [22]),
        .I1(\u1/out6 [22]),
        .O(\u1/R60 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[23]_i_1 
       (.I0(\u1/L5 [23]),
        .I1(\u1/out6 [23]),
        .O(\u1/R60 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[24]_i_1 
       (.I0(\u1/L5 [24]),
        .I1(\u1/out6 [24]),
        .O(\u1/R60 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[25]_i_1 
       (.I0(\u1/L5 [25]),
        .I1(\u1/out6 [25]),
        .O(\u1/R60 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[26]_i_1 
       (.I0(\u1/L5 [26]),
        .I1(\u1/out6 [26]),
        .O(\u1/R60 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[27]_i_1 
       (.I0(\u1/L5 [27]),
        .I1(\u1/out6 [27]),
        .O(\u1/R60 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[28]_i_1 
       (.I0(\u1/L5 [28]),
        .I1(\u1/out6 [28]),
        .O(\u1/R60 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[29]_i_1 
       (.I0(\u1/L5 [29]),
        .I1(\u1/out6 [29]),
        .O(\u1/R60 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[2]_i_1 
       (.I0(\u1/L5 [2]),
        .I1(\u1/out6 [2]),
        .O(\u1/R60 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[30]_i_1 
       (.I0(\u1/L5 [30]),
        .I1(\u1/out6 [30]),
        .O(\u1/R60 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[31]_i_1 
       (.I0(\u1/L5 [31]),
        .I1(\u1/out6 [31]),
        .O(\u1/R60 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[32]_i_1 
       (.I0(\u1/L5 [32]),
        .I1(\u1/out6 [32]),
        .O(\u1/R60 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[3]_i_1 
       (.I0(\u1/L5 [3]),
        .I1(\u1/out6 [3]),
        .O(\u1/R60 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[4]_i_1 
       (.I0(\u1/L5 [4]),
        .I1(\u1/out6 [4]),
        .O(\u1/R60 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[5]_i_1 
       (.I0(\u1/L5 [5]),
        .I1(\u1/out6 [5]),
        .O(\u1/R60 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[6]_i_1 
       (.I0(\u1/L5 [6]),
        .I1(\u1/out6 [6]),
        .O(\u1/R60 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[7]_i_1 
       (.I0(\u1/L5 [7]),
        .I1(\u1/out6 [7]),
        .O(\u1/R60 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[8]_i_1 
       (.I0(\u1/L5 [8]),
        .I1(\u1/out6 [8]),
        .O(\u1/R60 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R6[9]_i_1 
       (.I0(\u1/L5 [9]),
        .I1(\u1/out6 [9]),
        .O(\u1/R60 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [22]),
        .Q(\u1/R6 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [21]),
        .Q(\u1/R6 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [20]),
        .Q(\u1/R6 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [19]),
        .Q(\u1/R6 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [18]),
        .Q(\u1/R6 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [17]),
        .Q(\u1/R6 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [16]),
        .Q(\u1/R6 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [15]),
        .Q(\u1/R6 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [14]),
        .Q(\u1/R6 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [13]),
        .Q(\u1/R6 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [31]),
        .Q(\u1/R6 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [12]),
        .Q(\u1/R6 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [11]),
        .Q(\u1/R6 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [10]),
        .Q(\u1/R6 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [9]),
        .Q(\u1/R6 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [8]),
        .Q(\u1/R6 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [7]),
        .Q(\u1/R6 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [6]),
        .Q(\u1/R6 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [5]),
        .Q(\u1/R6 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [4]),
        .Q(\u1/R6 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [3]),
        .Q(\u1/R6 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [30]),
        .Q(\u1/R6 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [2]),
        .Q(\u1/R6 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [1]),
        .Q(\u1/R6 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [0]),
        .Q(\u1/R6 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [29]),
        .Q(\u1/R6 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [28]),
        .Q(\u1/R6 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [27]),
        .Q(\u1/R6 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [26]),
        .Q(\u1/R6 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [25]),
        .Q(\u1/R6 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [24]),
        .Q(\u1/R6 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R6_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R60 [23]),
        .Q(\u1/R6 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[10]_i_1 
       (.I0(\u1/L6 [10]),
        .I1(\u1/out7 [10]),
        .O(\u1/R70 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[11]_i_1 
       (.I0(\u1/L6 [11]),
        .I1(\u1/out7 [11]),
        .O(\u1/R70 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[12]_i_1 
       (.I0(\u1/L6 [12]),
        .I1(\u1/out7 [12]),
        .O(\u1/R70 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[13]_i_1 
       (.I0(\u1/L6 [13]),
        .I1(\u1/out7 [13]),
        .O(\u1/R70 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[14]_i_1 
       (.I0(\u1/L6 [14]),
        .I1(\u1/out7 [14]),
        .O(\u1/R70 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[15]_i_1 
       (.I0(\u1/L6 [15]),
        .I1(\u1/out7 [15]),
        .O(\u1/R70 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[16]_i_1 
       (.I0(\u1/L6 [16]),
        .I1(\u1/out7 [16]),
        .O(\u1/R70 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[17]_i_1 
       (.I0(\u1/L6 [17]),
        .I1(\u1/out7 [17]),
        .O(\u1/R70 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[18]_i_1 
       (.I0(\u1/L6 [18]),
        .I1(\u1/out7 [18]),
        .O(\u1/R70 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[19]_i_1 
       (.I0(\u1/L6 [19]),
        .I1(\u1/out7 [19]),
        .O(\u1/R70 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[1]_i_1 
       (.I0(\u1/L6 [1]),
        .I1(\u1/out7 [1]),
        .O(\u1/R70 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[20]_i_1 
       (.I0(\u1/L6 [20]),
        .I1(\u1/out7 [20]),
        .O(\u1/R70 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[21]_i_1 
       (.I0(\u1/L6 [21]),
        .I1(\u1/out7 [21]),
        .O(\u1/R70 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[22]_i_1 
       (.I0(\u1/L6 [22]),
        .I1(\u1/out7 [22]),
        .O(\u1/R70 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[23]_i_1 
       (.I0(\u1/L6 [23]),
        .I1(\u1/out7 [23]),
        .O(\u1/R70 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[24]_i_1 
       (.I0(\u1/L6 [24]),
        .I1(\u1/out7 [24]),
        .O(\u1/R70 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[25]_i_1 
       (.I0(\u1/L6 [25]),
        .I1(\u1/out7 [25]),
        .O(\u1/R70 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[26]_i_1 
       (.I0(\u1/L6 [26]),
        .I1(\u1/out7 [26]),
        .O(\u1/R70 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[27]_i_1 
       (.I0(\u1/L6 [27]),
        .I1(\u1/out7 [27]),
        .O(\u1/R70 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[28]_i_1 
       (.I0(\u1/L6 [28]),
        .I1(\u1/out7 [28]),
        .O(\u1/R70 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[29]_i_1 
       (.I0(\u1/L6 [29]),
        .I1(\u1/out7 [29]),
        .O(\u1/R70 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[2]_i_1 
       (.I0(\u1/L6 [2]),
        .I1(\u1/out7 [2]),
        .O(\u1/R70 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[30]_i_1 
       (.I0(\u1/L6 [30]),
        .I1(\u1/out7 [30]),
        .O(\u1/R70 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[31]_i_1 
       (.I0(\u1/L6 [31]),
        .I1(\u1/out7 [31]),
        .O(\u1/R70 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[32]_i_1 
       (.I0(\u1/L6 [32]),
        .I1(\u1/out7 [32]),
        .O(\u1/R70 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[3]_i_1 
       (.I0(\u1/L6 [3]),
        .I1(\u1/out7 [3]),
        .O(\u1/R70 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[4]_i_1 
       (.I0(\u1/L6 [4]),
        .I1(\u1/out7 [4]),
        .O(\u1/R70 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[5]_i_1 
       (.I0(\u1/L6 [5]),
        .I1(\u1/out7 [5]),
        .O(\u1/R70 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[6]_i_1 
       (.I0(\u1/L6 [6]),
        .I1(\u1/out7 [6]),
        .O(\u1/R70 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[7]_i_1 
       (.I0(\u1/L6 [7]),
        .I1(\u1/out7 [7]),
        .O(\u1/R70 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[8]_i_1 
       (.I0(\u1/L6 [8]),
        .I1(\u1/out7 [8]),
        .O(\u1/R70 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R7[9]_i_1 
       (.I0(\u1/L6 [9]),
        .I1(\u1/out7 [9]),
        .O(\u1/R70 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [22]),
        .Q(\u1/R7 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [21]),
        .Q(\u1/R7 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [20]),
        .Q(\u1/R7 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [19]),
        .Q(\u1/R7 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [18]),
        .Q(\u1/R7 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [17]),
        .Q(\u1/R7 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [16]),
        .Q(\u1/R7 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [15]),
        .Q(\u1/R7 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [14]),
        .Q(\u1/R7 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [13]),
        .Q(\u1/R7 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [31]),
        .Q(\u1/R7 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [12]),
        .Q(\u1/R7 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [11]),
        .Q(\u1/R7 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [10]),
        .Q(\u1/R7 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [9]),
        .Q(\u1/R7 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [8]),
        .Q(\u1/R7 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [7]),
        .Q(\u1/R7 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [6]),
        .Q(\u1/R7 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [5]),
        .Q(\u1/R7 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [4]),
        .Q(\u1/R7 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [3]),
        .Q(\u1/R7 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [30]),
        .Q(\u1/R7 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [2]),
        .Q(\u1/R7 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [1]),
        .Q(\u1/R7 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [0]),
        .Q(\u1/R7 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [29]),
        .Q(\u1/R7 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [28]),
        .Q(\u1/R7 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [27]),
        .Q(\u1/R7 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [26]),
        .Q(\u1/R7 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [25]),
        .Q(\u1/R7 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [24]),
        .Q(\u1/R7 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R7_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R70 [23]),
        .Q(\u1/R7 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[10]_i_1 
       (.I0(\u1/L7 [10]),
        .I1(\u1/out8 [10]),
        .O(\u1/R80 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[11]_i_1 
       (.I0(\u1/L7 [11]),
        .I1(\u1/out8 [11]),
        .O(\u1/R80 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[12]_i_1 
       (.I0(\u1/L7 [12]),
        .I1(\u1/out8 [12]),
        .O(\u1/R80 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[13]_i_1 
       (.I0(\u1/L7 [13]),
        .I1(\u1/out8 [13]),
        .O(\u1/R80 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[14]_i_1 
       (.I0(\u1/L7 [14]),
        .I1(\u1/out8 [14]),
        .O(\u1/R80 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[15]_i_1 
       (.I0(\u1/L7 [15]),
        .I1(\u1/out8 [15]),
        .O(\u1/R80 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[16]_i_1 
       (.I0(\u1/L7 [16]),
        .I1(\u1/out8 [16]),
        .O(\u1/R80 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[17]_i_1 
       (.I0(\u1/L7 [17]),
        .I1(\u1/out8 [17]),
        .O(\u1/R80 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[18]_i_1 
       (.I0(\u1/L7 [18]),
        .I1(\u1/out8 [18]),
        .O(\u1/R80 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[19]_i_1 
       (.I0(\u1/L7 [19]),
        .I1(\u1/out8 [19]),
        .O(\u1/R80 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[1]_i_1 
       (.I0(\u1/L7 [1]),
        .I1(\u1/out8 [1]),
        .O(\u1/R80 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[20]_i_1 
       (.I0(\u1/L7 [20]),
        .I1(\u1/out8 [20]),
        .O(\u1/R80 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[21]_i_1 
       (.I0(\u1/L7 [21]),
        .I1(\u1/out8 [21]),
        .O(\u1/R80 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[22]_i_1 
       (.I0(\u1/L7 [22]),
        .I1(\u1/out8 [22]),
        .O(\u1/R80 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[23]_i_1 
       (.I0(\u1/L7 [23]),
        .I1(\u1/out8 [23]),
        .O(\u1/R80 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[24]_i_1 
       (.I0(\u1/L7 [24]),
        .I1(\u1/out8 [24]),
        .O(\u1/R80 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[25]_i_1 
       (.I0(\u1/L7 [25]),
        .I1(\u1/out8 [25]),
        .O(\u1/R80 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[26]_i_1 
       (.I0(\u1/L7 [26]),
        .I1(\u1/out8 [26]),
        .O(\u1/R80 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[27]_i_1 
       (.I0(\u1/L7 [27]),
        .I1(\u1/out8 [27]),
        .O(\u1/R80 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[28]_i_1 
       (.I0(\u1/L7 [28]),
        .I1(\u1/out8 [28]),
        .O(\u1/R80 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[29]_i_1 
       (.I0(\u1/L7 [29]),
        .I1(\u1/out8 [29]),
        .O(\u1/R80 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[2]_i_1 
       (.I0(\u1/L7 [2]),
        .I1(\u1/out8 [2]),
        .O(\u1/R80 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[30]_i_1 
       (.I0(\u1/L7 [30]),
        .I1(\u1/out8 [30]),
        .O(\u1/R80 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[31]_i_1 
       (.I0(\u1/L7 [31]),
        .I1(\u1/out8 [31]),
        .O(\u1/R80 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[32]_i_1 
       (.I0(\u1/L7 [32]),
        .I1(\u1/out8 [32]),
        .O(\u1/R80 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[3]_i_1 
       (.I0(\u1/L7 [3]),
        .I1(\u1/out8 [3]),
        .O(\u1/R80 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[4]_i_1 
       (.I0(\u1/L7 [4]),
        .I1(\u1/out8 [4]),
        .O(\u1/R80 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[5]_i_1 
       (.I0(\u1/L7 [5]),
        .I1(\u1/out8 [5]),
        .O(\u1/R80 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[6]_i_1 
       (.I0(\u1/L7 [6]),
        .I1(\u1/out8 [6]),
        .O(\u1/R80 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[7]_i_1 
       (.I0(\u1/L7 [7]),
        .I1(\u1/out8 [7]),
        .O(\u1/R80 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[8]_i_1 
       (.I0(\u1/L7 [8]),
        .I1(\u1/out8 [8]),
        .O(\u1/R80 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R8[9]_i_1 
       (.I0(\u1/L7 [9]),
        .I1(\u1/out8 [9]),
        .O(\u1/R80 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [22]),
        .Q(\u1/R8 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [21]),
        .Q(\u1/R8 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [20]),
        .Q(\u1/R8 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [19]),
        .Q(\u1/R8 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [18]),
        .Q(\u1/R8 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [17]),
        .Q(\u1/R8 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [16]),
        .Q(\u1/R8 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [15]),
        .Q(\u1/R8 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [14]),
        .Q(\u1/R8 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [13]),
        .Q(\u1/R8 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [31]),
        .Q(\u1/R8 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [12]),
        .Q(\u1/R8 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [11]),
        .Q(\u1/R8 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [10]),
        .Q(\u1/R8 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [9]),
        .Q(\u1/R8 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [8]),
        .Q(\u1/R8 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [7]),
        .Q(\u1/R8 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [6]),
        .Q(\u1/R8 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [5]),
        .Q(\u1/R8 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [4]),
        .Q(\u1/R8 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [3]),
        .Q(\u1/R8 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [30]),
        .Q(\u1/R8 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [2]),
        .Q(\u1/R8 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [1]),
        .Q(\u1/R8 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [0]),
        .Q(\u1/R8 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [29]),
        .Q(\u1/R8 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [28]),
        .Q(\u1/R8 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [27]),
        .Q(\u1/R8 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [26]),
        .Q(\u1/R8 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [25]),
        .Q(\u1/R8 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [24]),
        .Q(\u1/R8 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R8_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R80 [23]),
        .Q(\u1/R8 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[10]_i_1 
       (.I0(\u1/L8 [10]),
        .I1(\u1/out9 [10]),
        .O(\u1/R90 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[11]_i_1 
       (.I0(\u1/L8 [11]),
        .I1(\u1/out9 [11]),
        .O(\u1/R90 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[12]_i_1 
       (.I0(\u1/L8 [12]),
        .I1(\u1/out9 [12]),
        .O(\u1/R90 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[13]_i_1 
       (.I0(\u1/L8 [13]),
        .I1(\u1/out9 [13]),
        .O(\u1/R90 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[14]_i_1 
       (.I0(\u1/L8 [14]),
        .I1(\u1/out9 [14]),
        .O(\u1/R90 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[15]_i_1 
       (.I0(\u1/L8 [15]),
        .I1(\u1/out9 [15]),
        .O(\u1/R90 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[16]_i_1 
       (.I0(\u1/L8 [16]),
        .I1(\u1/out9 [16]),
        .O(\u1/R90 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[17]_i_1 
       (.I0(\u1/L8 [17]),
        .I1(\u1/out9 [17]),
        .O(\u1/R90 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[18]_i_1 
       (.I0(\u1/L8 [18]),
        .I1(\u1/out9 [18]),
        .O(\u1/R90 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[19]_i_1 
       (.I0(\u1/L8 [19]),
        .I1(\u1/out9 [19]),
        .O(\u1/R90 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[1]_i_1 
       (.I0(\u1/L8 [1]),
        .I1(\u1/out9 [1]),
        .O(\u1/R90 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[20]_i_1 
       (.I0(\u1/L8 [20]),
        .I1(\u1/out9 [20]),
        .O(\u1/R90 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[21]_i_1 
       (.I0(\u1/L8 [21]),
        .I1(\u1/out9 [21]),
        .O(\u1/R90 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[22]_i_1 
       (.I0(\u1/L8 [22]),
        .I1(\u1/out9 [22]),
        .O(\u1/R90 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[23]_i_1 
       (.I0(\u1/L8 [23]),
        .I1(\u1/out9 [23]),
        .O(\u1/R90 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[24]_i_1 
       (.I0(\u1/L8 [24]),
        .I1(\u1/out9 [24]),
        .O(\u1/R90 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[25]_i_1 
       (.I0(\u1/L8 [25]),
        .I1(\u1/out9 [25]),
        .O(\u1/R90 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[26]_i_1 
       (.I0(\u1/L8 [26]),
        .I1(\u1/out9 [26]),
        .O(\u1/R90 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[27]_i_1 
       (.I0(\u1/L8 [27]),
        .I1(\u1/out9 [27]),
        .O(\u1/R90 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[28]_i_1 
       (.I0(\u1/L8 [28]),
        .I1(\u1/out9 [28]),
        .O(\u1/R90 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[29]_i_1 
       (.I0(\u1/L8 [29]),
        .I1(\u1/out9 [29]),
        .O(\u1/R90 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[2]_i_1 
       (.I0(\u1/L8 [2]),
        .I1(\u1/out9 [2]),
        .O(\u1/R90 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[30]_i_1 
       (.I0(\u1/L8 [30]),
        .I1(\u1/out9 [30]),
        .O(\u1/R90 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[31]_i_1 
       (.I0(\u1/L8 [31]),
        .I1(\u1/out9 [31]),
        .O(\u1/R90 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[32]_i_1 
       (.I0(\u1/L8 [32]),
        .I1(\u1/out9 [32]),
        .O(\u1/R90 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[3]_i_1 
       (.I0(\u1/L8 [3]),
        .I1(\u1/out9 [3]),
        .O(\u1/R90 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[4]_i_1 
       (.I0(\u1/L8 [4]),
        .I1(\u1/out9 [4]),
        .O(\u1/R90 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[5]_i_1 
       (.I0(\u1/L8 [5]),
        .I1(\u1/out9 [5]),
        .O(\u1/R90 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[6]_i_1 
       (.I0(\u1/L8 [6]),
        .I1(\u1/out9 [6]),
        .O(\u1/R90 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[7]_i_1 
       (.I0(\u1/L8 [7]),
        .I1(\u1/out9 [7]),
        .O(\u1/R90 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[8]_i_1 
       (.I0(\u1/L8 [8]),
        .I1(\u1/out9 [8]),
        .O(\u1/R90 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/R9[9]_i_1 
       (.I0(\u1/L8 [9]),
        .I1(\u1/out9 [9]),
        .O(\u1/R90 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [22]),
        .Q(\u1/R9 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [21]),
        .Q(\u1/R9 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [20]),
        .Q(\u1/R9 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [19]),
        .Q(\u1/R9 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [18]),
        .Q(\u1/R9 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [17]),
        .Q(\u1/R9 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [16]),
        .Q(\u1/R9 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [15]),
        .Q(\u1/R9 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [14]),
        .Q(\u1/R9 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [13]),
        .Q(\u1/R9 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [31]),
        .Q(\u1/R9 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [12]),
        .Q(\u1/R9 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [11]),
        .Q(\u1/R9 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [10]),
        .Q(\u1/R9 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [9]),
        .Q(\u1/R9 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [8]),
        .Q(\u1/R9 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [7]),
        .Q(\u1/R9 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [6]),
        .Q(\u1/R9 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [5]),
        .Q(\u1/R9 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [4]),
        .Q(\u1/R9 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [3]),
        .Q(\u1/R9 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [30]),
        .Q(\u1/R9 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [2]),
        .Q(\u1/R9 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [1]),
        .Q(\u1/R9 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [0]),
        .Q(\u1/R9 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [29]),
        .Q(\u1/R9 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [28]),
        .Q(\u1/R9 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [27]),
        .Q(\u1/R9 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [26]),
        .Q(\u1/R9 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [25]),
        .Q(\u1/R9 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [24]),
        .Q(\u1/R9 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/R9_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/R90 [23]),
        .Q(\u1/R9 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[0]),
        .Q(\u1/IP [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[10]),
        .Q(\u1/IP [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[11]),
        .Q(\u1/IP [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[12]),
        .Q(\u1/IP [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[13]),
        .Q(\u1/IP [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[14]),
        .Q(\u1/IP [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[15]),
        .Q(\u1/IP [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[16]),
        .Q(\u1/IP [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[17]),
        .Q(\u1/IP [59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[18]),
        .Q(\u1/IP [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[19]),
        .Q(\u1/IP [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[1]),
        .Q(\u1/IP [57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[20]),
        .Q(\u1/IP [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[21]),
        .Q(\u1/IP [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[22]),
        .Q(\u1/IP [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[23]),
        .Q(\u1/IP [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[24]),
        .Q(\u1/IP [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[25]),
        .Q(\u1/IP [60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[26]),
        .Q(\u1/IP [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[27]),
        .Q(\u1/IP [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[28]),
        .Q(\u1/IP [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[29]),
        .Q(\u1/IP [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[2]),
        .Q(\u1/IP [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[30]),
        .Q(\u1/IP [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[31]),
        .Q(\u1/IP [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[32]),
        .Q(\u1/IP [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[33]),
        .Q(\u1/IP [61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[34]),
        .Q(\u1/IP [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[35]),
        .Q(\u1/IP [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[36]),
        .Q(\u1/IP [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[37]),
        .Q(\u1/IP [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[38]),
        .Q(\u1/IP [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[39]),
        .Q(\u1/IP [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[3]),
        .Q(\u1/IP [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[40]),
        .Q(\u1/IP [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[41]),
        .Q(\u1/IP [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[42]),
        .Q(\u1/IP [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[43]),
        .Q(\u1/IP [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[44]),
        .Q(\u1/IP [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[45]),
        .Q(\u1/IP [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[46]),
        .Q(\u1/IP [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[47]),
        .Q(\u1/IP [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[48]),
        .Q(\u1/IP [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[49]),
        .Q(\u1/IP [63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[4]),
        .Q(\u1/IP [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[50]),
        .Q(\u1/IP [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[51]),
        .Q(\u1/IP [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[52]),
        .Q(\u1/IP [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[53]),
        .Q(\u1/IP [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[54]),
        .Q(\u1/IP [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[55]),
        .Q(\u1/IP [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[56]),
        .Q(\u1/IP [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[57]),
        .Q(\u1/IP [64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[58]),
        .Q(\u1/IP [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[59]),
        .Q(\u1/IP [56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[5]),
        .Q(\u1/IP [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[60]),
        .Q(\u1/IP [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[61]),
        .Q(\u1/IP [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[62]),
        .Q(\u1/IP [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[63]),
        .Q(\u1/IP [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[6]),
        .Q(\u1/IP [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[7]),
        .Q(\u1/IP [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[8]),
        .Q(\u1/IP [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desIn_r_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage1_out[9]),
        .Q(\u1/IP [58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[0]_i_1 
       (.I0(\u1/out15 [25]),
        .I1(\u1/L14 [25]),
        .O(\u1/FP [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[10]_i_1 
       (.I0(\u1/out15 [18]),
        .I1(\u1/L14 [18]),
        .O(\u1/FP [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[12]_i_1 
       (.I0(\u1/out15 [10]),
        .I1(\u1/L14 [10]),
        .O(\u1/FP [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[14]_i_1 
       (.I0(\u1/out15 [2]),
        .I1(\u1/L14 [2]),
        .O(\u1/FP [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[16]_i_1 
       (.I0(\u1/out15 [27]),
        .I1(\u1/L14 [27]),
        .O(\u1/FP [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[18]_i_1 
       (.I0(\u1/out15 [19]),
        .I1(\u1/L14 [19]),
        .O(\u1/FP [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[20]_i_1 
       (.I0(\u1/out15 [11]),
        .I1(\u1/L14 [11]),
        .O(\u1/FP [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[22]_i_1 
       (.I0(\u1/out15 [3]),
        .I1(\u1/L14 [3]),
        .O(\u1/FP [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[24]_i_1 
       (.I0(\u1/out15 [28]),
        .I1(\u1/L14 [28]),
        .O(\u1/FP [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[26]_i_1 
       (.I0(\u1/out15 [20]),
        .I1(\u1/L14 [20]),
        .O(\u1/FP [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[28]_i_1 
       (.I0(\u1/out15 [12]),
        .I1(\u1/L14 [12]),
        .O(\u1/FP [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[2]_i_1 
       (.I0(\u1/out15 [17]),
        .I1(\u1/L14 [17]),
        .O(\u1/FP [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[30]_i_1 
       (.I0(\u1/out15 [4]),
        .I1(\u1/L14 [4]),
        .O(\u1/FP [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[32]_i_1 
       (.I0(\u1/out15 [29]),
        .I1(\u1/L14 [29]),
        .O(\u1/FP [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[34]_i_1 
       (.I0(\u1/out15 [21]),
        .I1(\u1/L14 [21]),
        .O(\u1/FP [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[36]_i_1 
       (.I0(\u1/out15 [13]),
        .I1(\u1/L14 [13]),
        .O(\u1/FP [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[38]_i_1 
       (.I0(\u1/out15 [5]),
        .I1(\u1/L14 [5]),
        .O(\u1/FP [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[40]_i_1 
       (.I0(\u1/out15 [30]),
        .I1(\u1/L14 [30]),
        .O(\u1/FP [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[42]_i_1 
       (.I0(\u1/out15 [22]),
        .I1(\u1/L14 [22]),
        .O(\u1/FP [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[44]_i_1 
       (.I0(\u1/out15 [14]),
        .I1(\u1/L14 [14]),
        .O(\u1/FP [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[46]_i_1 
       (.I0(\u1/out15 [6]),
        .I1(\u1/L14 [6]),
        .O(\u1/FP [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[48]_i_1 
       (.I0(\u1/out15 [31]),
        .I1(\u1/L14 [31]),
        .O(\u1/FP [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[4]_i_1 
       (.I0(\u1/out15 [9]),
        .I1(\u1/L14 [9]),
        .O(\u1/FP [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[50]_i_1 
       (.I0(\u1/out15 [23]),
        .I1(\u1/L14 [23]),
        .O(\u1/FP [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[52]_i_1 
       (.I0(\u1/out15 [15]),
        .I1(\u1/L14 [15]),
        .O(\u1/FP [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[54]_i_1 
       (.I0(\u1/out15 [7]),
        .I1(\u1/L14 [7]),
        .O(\u1/FP [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[56]_i_1 
       (.I0(\u1/out15 [32]),
        .I1(\u1/L14 [32]),
        .O(\u1/FP [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[58]_i_1 
       (.I0(\u1/out15 [24]),
        .I1(\u1/L14 [24]),
        .O(\u1/FP [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[60]_i_1 
       (.I0(\u1/out15 [16]),
        .I1(\u1/L14 [16]),
        .O(\u1/FP [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[62]_i_1 
       (.I0(\u1/out15 [8]),
        .I1(\u1/L14 [8]),
        .O(\u1/FP [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[6]_i_1 
       (.I0(\u1/out15 [1]),
        .I1(\u1/L14 [1]),
        .O(\u1/FP [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u1/desOut[8]_i_1 
       (.I0(\u1/out15 [26]),
        .I1(\u1/L14 [26]),
        .O(\u1/FP [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [25]),
        .Q(stage2_out[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [18]),
        .Q(stage2_out[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [50]),
        .Q(stage2_out[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [10]),
        .Q(stage2_out[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [42]),
        .Q(stage2_out[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [2]),
        .Q(stage2_out[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [34]),
        .Q(stage2_out[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [27]),
        .Q(stage2_out[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [59]),
        .Q(stage2_out[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [19]),
        .Q(stage2_out[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [51]),
        .Q(stage2_out[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [57]),
        .Q(stage2_out[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [11]),
        .Q(stage2_out[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [43]),
        .Q(stage2_out[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [3]),
        .Q(stage2_out[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [35]),
        .Q(stage2_out[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [28]),
        .Q(stage2_out[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [60]),
        .Q(stage2_out[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [20]),
        .Q(stage2_out[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [52]),
        .Q(stage2_out[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [12]),
        .Q(stage2_out[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [44]),
        .Q(stage2_out[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [17]),
        .Q(stage2_out[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [4]),
        .Q(stage2_out[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [36]),
        .Q(stage2_out[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [29]),
        .Q(stage2_out[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [61]),
        .Q(stage2_out[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [21]),
        .Q(stage2_out[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [53]),
        .Q(stage2_out[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [13]),
        .Q(stage2_out[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [45]),
        .Q(stage2_out[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [5]),
        .Q(stage2_out[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [37]),
        .Q(stage2_out[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [49]),
        .Q(stage2_out[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [30]),
        .Q(stage2_out[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [62]),
        .Q(stage2_out[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [22]),
        .Q(stage2_out[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [54]),
        .Q(stage2_out[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [14]),
        .Q(stage2_out[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [46]),
        .Q(stage2_out[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [6]),
        .Q(stage2_out[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [38]),
        .Q(stage2_out[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [31]),
        .Q(stage2_out[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [63]),
        .Q(stage2_out[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [9]),
        .Q(stage2_out[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [23]),
        .Q(stage2_out[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [55]),
        .Q(stage2_out[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [15]),
        .Q(stage2_out[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [47]),
        .Q(stage2_out[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [7]),
        .Q(stage2_out[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [39]),
        .Q(stage2_out[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [32]),
        .Q(stage2_out[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [64]),
        .Q(stage2_out[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [24]),
        .Q(stage2_out[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [56]),
        .Q(stage2_out[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [41]),
        .Q(stage2_out[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [16]),
        .Q(stage2_out[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [48]),
        .Q(stage2_out[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [8]),
        .Q(stage2_out[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [40]),
        .Q(stage2_out[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [1]),
        .Q(stage2_out[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [33]),
        .Q(stage2_out[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [26]),
        .Q(stage2_out[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/desOut_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/FP [58]),
        .Q(stage2_out[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(key_b_r_reg),
        .Q(\u1/key_r [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][10]_srl16_n_0 ),
        .Q(\u1/key_r [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][11]_srl16_n_0 ),
        .Q(\u1/key_r [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][12]_srl16_n_0 ),
        .Q(\u1/key_r [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][13]_srl16_n_0 ),
        .Q(\u1/key_r [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][14]_srl16_n_0 ),
        .Q(\u1/key_r [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][15]_srl16_n_0 ),
        .Q(\u1/key_r [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][16]_srl16_n_0 ),
        .Q(\u1/key_r [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][17]_srl16_n_0 ),
        .Q(\u1/key_r [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][18]_srl16_n_0 ),
        .Q(\u1/key_r [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][19]_srl16_n_0 ),
        .Q(\u1/key_r [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][1]_srl16_n_0 ),
        .Q(\u1/key_r [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][20]_srl16_n_0 ),
        .Q(\u1/key_r [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][21]_srl16_n_0 ),
        .Q(\u1/key_r [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][22]_srl16_n_0 ),
        .Q(\u1/key_r [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][23]_srl16_n_0 ),
        .Q(\u1/key_r [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][24]_srl16_n_0 ),
        .Q(\u1/key_r [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][25]_srl16_n_0 ),
        .Q(\u1/key_r [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][26]_srl16_n_0 ),
        .Q(\u1/key_r [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][27]_srl16_n_0 ),
        .Q(\u1/key_r [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][28]_srl16_n_0 ),
        .Q(\u1/key_r [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][29]_srl16_n_0 ),
        .Q(\u1/key_r [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][2]_srl16_n_0 ),
        .Q(\u1/key_r [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][30]_srl16_n_0 ),
        .Q(\u1/key_r [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][31]_srl16_n_0 ),
        .Q(\u1/key_r [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][32]_srl16_n_0 ),
        .Q(\u1/key_r [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][33]_srl16_n_0 ),
        .Q(\u1/key_r [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][34]_srl16_n_0 ),
        .Q(\u1/key_r [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][35]_srl16_n_0 ),
        .Q(\u1/key_r [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][36]_srl16_n_0 ),
        .Q(\u1/key_r [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][37]_srl16_n_0 ),
        .Q(\u1/key_r [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][38]_srl16_n_0 ),
        .Q(\u1/key_r [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][39]_srl16_n_0 ),
        .Q(\u1/key_r [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][3]_srl16_n_0 ),
        .Q(\u1/key_r [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][40]_srl16_n_0 ),
        .Q(\u1/key_r [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][41]_srl16_n_0 ),
        .Q(\u1/key_r [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][42]_srl16_n_0 ),
        .Q(\u1/key_r [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][43]_srl16_n_0 ),
        .Q(\u1/key_r [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][44]_srl16_n_0 ),
        .Q(\u1/key_r [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][45]_srl16_n_0 ),
        .Q(\u1/key_r [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][46]_srl16_n_0 ),
        .Q(\u1/key_r [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][47]_srl16_n_0 ),
        .Q(\u1/key_r [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][48]_srl16_n_0 ),
        .Q(\u1/key_r [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][49]_srl16_n_0 ),
        .Q(\u1/key_r [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][4]_srl16_n_0 ),
        .Q(\u1/key_r [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][50]_srl16_n_0 ),
        .Q(\u1/key_r [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][51]_srl16_n_0 ),
        .Q(\u1/key_r [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][52]_srl16_n_0 ),
        .Q(\u1/key_r [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][53]_srl16_n_0 ),
        .Q(\u1/key_r [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][54]_srl16_n_0 ),
        .Q(\u1/key_r [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][55]_srl16_n_0 ),
        .Q(\u1/key_r [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][5]_srl16_n_0 ),
        .Q(\u1/key_r [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][6]_srl16_n_0 ),
        .Q(\u1/key_r [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][7]_srl16_n_0 ),
        .Q(\u1/key_r [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][8]_srl16_n_0 ),
        .Q(\u1/key_r [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/key_r_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_b_r_reg[16][9]_srl16_n_0 ),
        .Q(\u1/key_r [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [0]),
        .Q(\u1/uk/K_r0_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [10]),
        .Q(\u1/uk/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [11]),
        .Q(\u1/uk/p_14_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [12]),
        .Q(\u1/uk/p_38_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [13]),
        .Q(\u1/uk/p_7_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [14]),
        .Q(\u1/uk/p_36_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [15]),
        .Q(\u1/uk/p_25_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [16]),
        .Q(\u1/uk/p_27_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [17]),
        .Q(\u1/uk/K_r0_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [18]),
        .Q(\u1/uk/p_37_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [19]),
        .Q(\u1/uk/K_r0_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [1]),
        .Q(\u1/uk/K_r0_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [20]),
        .Q(\u1/uk/p_2_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [21]),
        .Q(\u1/uk/p_24_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [22]),
        .Q(\u1/uk/K_r0_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [23]),
        .Q(\u1/uk/p_30_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [24]),
        .Q(\u1/uk/p_3_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [25]),
        .Q(\u1/uk/K_r0_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [26]),
        .Q(\u1/uk/p_9_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [27]),
        .Q(\u1/uk/p_5_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [28]),
        .Q(\u1/uk/p_20_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [29]),
        .Q(\u1/uk/p_31_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [2]),
        .Q(\u1/uk/K_r0_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [30]),
        .Q(\u1/uk/p_22_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [31]),
        .Q(\u1/uk/K_r0_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [32]),
        .Q(\u1/uk/K_r0_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [33]),
        .Q(\u1/uk/p_39_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [34]),
        .Q(\u1/uk/p_6_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [35]),
        .Q(\u1/uk/K_r0_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [36]),
        .Q(\u1/uk/K_r0_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [37]),
        .Q(\u1/uk/p_26_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [38]),
        .Q(\u1/uk/p_18_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [39]),
        .Q(\u1/uk/p_12_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [3]),
        .Q(\u1/uk/p_11_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [40]),
        .Q(\u1/uk/p_8_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [41]),
        .Q(\u1/uk/p_13_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [42]),
        .Q(\u1/uk/p_29_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [43]),
        .Q(\u1/uk/p_17_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [44]),
        .Q(\u1/uk/p_19_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [45]),
        .Q(\u1/uk/p_33_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [46]),
        .Q(\u1/uk/p_1_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [47]),
        .Q(\u1/uk/p_15_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [48]),
        .Q(\u1/uk/p_4_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [49]),
        .Q(\u1/uk/p_34_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [4]),
        .Q(\u1/uk/K_r0_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [50]),
        .Q(\u1/uk/p_28_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [51]),
        .Q(\u1/uk/p_35_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [52]),
        .Q(\u1/uk/K_r0_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [53]),
        .Q(\u1/uk/K_r0_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [54]),
        .Q(\u1/uk/p_40_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [55]),
        .Q(\u1/uk/K_r0_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [5]),
        .Q(\u1/uk/p_10_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [6]),
        .Q(\u1/uk/p_16_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [7]),
        .Q(\u1/uk/p_21_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [8]),
        .Q(\u1/uk/p_32_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r0_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/key_r [9]),
        .Q(\u1/uk/p_23_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [0]),
        .Q(\u1/uk/K_r10 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [10]),
        .Q(\u1/uk/K_r10 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [11]),
        .Q(\u1/uk/K_r10 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [12]),
        .Q(\u1/uk/K_r10 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [13]),
        .Q(\u1/uk/K_r10 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [14]),
        .Q(\u1/uk/K_r10 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [15]),
        .Q(\u1/uk/K_r10 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [16]),
        .Q(\u1/uk/K_r10 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [17]),
        .Q(\u1/uk/K_r10 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [18]),
        .Q(\u1/uk/K_r10 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [19]),
        .Q(\u1/uk/K_r10 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [1]),
        .Q(\u1/uk/K_r10 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [20]),
        .Q(\u1/uk/K_r10 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [21]),
        .Q(\u1/uk/K_r10 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [22]),
        .Q(\u1/uk/K_r10 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [23]),
        .Q(\u1/uk/K_r10 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [24]),
        .Q(\u1/uk/K_r10 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [25]),
        .Q(\u1/uk/K_r10 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [26]),
        .Q(\u1/uk/K_r10 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [27]),
        .Q(\u1/uk/K_r10 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [28]),
        .Q(\u1/uk/K_r10 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [29]),
        .Q(\u1/uk/K_r10 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [2]),
        .Q(\u1/uk/K_r10 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [30]),
        .Q(\u1/uk/K_r10 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [31]),
        .Q(\u1/uk/K_r10 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [32]),
        .Q(\u1/uk/K_r10 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [33]),
        .Q(\u1/uk/K_r10 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [34]),
        .Q(\u1/uk/K_r10 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [35]),
        .Q(\u1/uk/K_r10 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [36]),
        .Q(\u1/uk/K_r10 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [37]),
        .Q(\u1/uk/K_r10 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [38]),
        .Q(\u1/uk/K_r10 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [39]),
        .Q(\u1/uk/K_r10 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [3]),
        .Q(\u1/uk/K_r10 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [40]),
        .Q(\u1/uk/K_r10 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [41]),
        .Q(\u1/uk/K_r10 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [42]),
        .Q(\u1/uk/K_r10 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [43]),
        .Q(\u1/uk/K_r10 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [44]),
        .Q(\u1/uk/K_r10 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [45]),
        .Q(\u1/uk/K_r10 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [46]),
        .Q(\u1/uk/K_r10 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [47]),
        .Q(\u1/uk/K_r10 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [48]),
        .Q(\u1/uk/K_r10 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [49]),
        .Q(\u1/uk/K_r10 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [4]),
        .Q(\u1/uk/K_r10 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [50]),
        .Q(\u1/uk/K_r10 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [51]),
        .Q(\u1/uk/K_r10 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [52]),
        .Q(\u1/uk/K_r10 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [53]),
        .Q(\u1/uk/K_r10 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [54]),
        .Q(\u1/uk/K_r10 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [55]),
        .Q(\u1/uk/K_r10 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [5]),
        .Q(\u1/uk/K_r10 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [6]),
        .Q(\u1/uk/K_r10 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [7]),
        .Q(\u1/uk/K_r10 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [8]),
        .Q(\u1/uk/K_r10 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r10_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r9 [9]),
        .Q(\u1/uk/K_r10 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [0]),
        .Q(\u1/uk/K_r11 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [10]),
        .Q(\u1/uk/K_r11 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [11]),
        .Q(\u1/uk/K_r11 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [12]),
        .Q(\u1/uk/K_r11 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [13]),
        .Q(\u1/uk/K_r11 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [14]),
        .Q(\u1/uk/K_r11 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [15]),
        .Q(\u1/uk/K_r11 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [16]),
        .Q(\u1/uk/K_r11 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [17]),
        .Q(\u1/uk/K_r11 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [18]),
        .Q(\u1/uk/K_r11 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [19]),
        .Q(\u1/uk/K_r11 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [1]),
        .Q(\u1/uk/K_r11 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [20]),
        .Q(\u1/uk/K_r11 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [21]),
        .Q(\u1/uk/K_r11 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [22]),
        .Q(\u1/uk/K_r11 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [23]),
        .Q(\u1/uk/K_r11 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [24]),
        .Q(\u1/uk/K_r11 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [25]),
        .Q(\u1/uk/K_r11 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [26]),
        .Q(\u1/uk/K_r11 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [27]),
        .Q(\u1/uk/K_r11 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [28]),
        .Q(\u1/uk/K_r11 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [29]),
        .Q(\u1/uk/K_r11 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [2]),
        .Q(\u1/uk/K_r11 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [30]),
        .Q(\u1/uk/K_r11 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [31]),
        .Q(\u1/uk/K_r11 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [32]),
        .Q(\u1/uk/K_r11 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [33]),
        .Q(\u1/uk/K_r11 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [34]),
        .Q(\u1/uk/K_r11 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [35]),
        .Q(\u1/uk/K_r11 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [36]),
        .Q(\u1/uk/K_r11 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [37]),
        .Q(\u1/uk/K_r11 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [38]),
        .Q(\u1/uk/K_r11 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [39]),
        .Q(\u1/uk/K_r11 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [3]),
        .Q(\u1/uk/K_r11 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [40]),
        .Q(\u1/uk/K_r11 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [41]),
        .Q(\u1/uk/K_r11 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [42]),
        .Q(\u1/uk/K_r11 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [43]),
        .Q(\u1/uk/K_r11 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [44]),
        .Q(\u1/uk/K_r11 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [45]),
        .Q(\u1/uk/K_r11 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [46]),
        .Q(\u1/uk/K_r11 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [47]),
        .Q(\u1/uk/K_r11 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [48]),
        .Q(\u1/uk/K_r11 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [49]),
        .Q(\u1/uk/K_r11 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [4]),
        .Q(\u1/uk/K_r11 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [50]),
        .Q(\u1/uk/K_r11 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [51]),
        .Q(\u1/uk/K_r11 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [52]),
        .Q(\u1/uk/K_r11 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [53]),
        .Q(\u1/uk/K_r11 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [54]),
        .Q(\u1/uk/K_r11 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [55]),
        .Q(\u1/uk/K_r11 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [5]),
        .Q(\u1/uk/K_r11 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [6]),
        .Q(\u1/uk/K_r11 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [7]),
        .Q(\u1/uk/K_r11 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [8]),
        .Q(\u1/uk/K_r11 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r11_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r10 [9]),
        .Q(\u1/uk/K_r11 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [0]),
        .Q(\u1/uk/K_r12 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [10]),
        .Q(\u1/uk/K_r12 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [11]),
        .Q(\u1/uk/K_r12 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [12]),
        .Q(\u1/uk/K_r12 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [13]),
        .Q(\u1/uk/K_r12 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [14]),
        .Q(\u1/uk/K_r12 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [15]),
        .Q(\u1/uk/K_r12 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [16]),
        .Q(\u1/uk/K_r12 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [17]),
        .Q(\u1/uk/K_r12 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [18]),
        .Q(\u1/uk/K_r12 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [19]),
        .Q(\u1/uk/K_r12 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [1]),
        .Q(\u1/uk/K_r12 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [20]),
        .Q(\u1/uk/K_r12 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [21]),
        .Q(\u1/uk/K_r12 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [22]),
        .Q(\u1/uk/K_r12 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [23]),
        .Q(\u1/uk/K_r12 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [24]),
        .Q(\u1/uk/K_r12 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [25]),
        .Q(\u1/uk/K_r12 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [26]),
        .Q(\u1/uk/K_r12 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [27]),
        .Q(\u1/uk/K_r12 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [28]),
        .Q(\u1/uk/K_r12 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [29]),
        .Q(\u1/uk/K_r12 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [2]),
        .Q(\u1/uk/K_r12 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [30]),
        .Q(\u1/uk/K_r12 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [31]),
        .Q(\u1/uk/K_r12 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [32]),
        .Q(\u1/uk/K_r12 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [33]),
        .Q(\u1/uk/K_r12 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [34]),
        .Q(\u1/uk/K_r12 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [35]),
        .Q(\u1/uk/K_r12 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [36]),
        .Q(\u1/uk/K_r12 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [37]),
        .Q(\u1/uk/K_r12 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [38]),
        .Q(\u1/uk/K_r12 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [39]),
        .Q(\u1/uk/K_r12 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [3]),
        .Q(\u1/uk/K_r12 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [40]),
        .Q(\u1/uk/K_r12 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [41]),
        .Q(\u1/uk/K_r12 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [42]),
        .Q(\u1/uk/K_r12 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [43]),
        .Q(\u1/uk/K_r12 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [44]),
        .Q(\u1/uk/K_r12 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [45]),
        .Q(\u1/uk/K_r12 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [46]),
        .Q(\u1/uk/K_r12 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [47]),
        .Q(\u1/uk/K_r12 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [48]),
        .Q(\u1/uk/K_r12 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [49]),
        .Q(\u1/uk/K_r12 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [4]),
        .Q(\u1/uk/K_r12 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [50]),
        .Q(\u1/uk/K_r12 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [51]),
        .Q(\u1/uk/K_r12 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [52]),
        .Q(\u1/uk/K_r12 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [53]),
        .Q(\u1/uk/K_r12 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [54]),
        .Q(\u1/uk/K_r12 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [55]),
        .Q(\u1/uk/K_r12 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [5]),
        .Q(\u1/uk/K_r12 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [6]),
        .Q(\u1/uk/K_r12 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [7]),
        .Q(\u1/uk/K_r12 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [8]),
        .Q(\u1/uk/K_r12 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r12_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r11 [9]),
        .Q(\u1/uk/K_r12 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [0]),
        .Q(\u1/uk/K_r13 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [10]),
        .Q(\u1/uk/K_r13 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [11]),
        .Q(\u1/uk/K_r13 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [12]),
        .Q(\u1/uk/K_r13 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [13]),
        .Q(\u1/uk/K_r13 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [14]),
        .Q(\u1/uk/K_r13 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [15]),
        .Q(\u1/uk/K_r13 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [16]),
        .Q(\u1/uk/K_r13 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [17]),
        .Q(\u1/uk/K_r13 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [18]),
        .Q(\u1/uk/K_r13 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [19]),
        .Q(\u1/uk/K_r13 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [1]),
        .Q(\u1/uk/K_r13 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [20]),
        .Q(\u1/uk/K_r13 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [21]),
        .Q(\u1/uk/K_r13 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [22]),
        .Q(\u1/uk/K_r13 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [23]),
        .Q(\u1/uk/K_r13 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [24]),
        .Q(\u1/uk/K_r13 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [25]),
        .Q(\u1/uk/K_r13 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [26]),
        .Q(\u1/uk/K_r13 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [27]),
        .Q(\u1/uk/K_r13 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [28]),
        .Q(\u1/uk/K_r13 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [29]),
        .Q(\u1/uk/K_r13 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [2]),
        .Q(\u1/uk/K_r13 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [30]),
        .Q(\u1/uk/K_r13 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [31]),
        .Q(\u1/uk/K_r13 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [32]),
        .Q(\u1/uk/K_r13 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [33]),
        .Q(\u1/uk/K_r13 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [34]),
        .Q(\u1/uk/K_r13 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [35]),
        .Q(\u1/uk/K_r13 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [36]),
        .Q(\u1/uk/K_r13 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [37]),
        .Q(\u1/uk/K_r13 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [38]),
        .Q(\u1/uk/K_r13 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [39]),
        .Q(\u1/uk/K_r13 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [3]),
        .Q(\u1/uk/K_r13 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [40]),
        .Q(\u1/uk/K_r13 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [41]),
        .Q(\u1/uk/K_r13 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [42]),
        .Q(\u1/uk/K_r13 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [43]),
        .Q(\u1/uk/K_r13 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [44]),
        .Q(\u1/uk/K_r13 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [45]),
        .Q(\u1/uk/K_r13 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [46]),
        .Q(\u1/uk/K_r13 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [47]),
        .Q(\u1/uk/K_r13 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [48]),
        .Q(\u1/uk/K_r13 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [49]),
        .Q(\u1/uk/K_r13 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [4]),
        .Q(\u1/uk/K_r13 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [50]),
        .Q(\u1/uk/K_r13 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [51]),
        .Q(\u1/uk/K_r13 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [52]),
        .Q(\u1/uk/K_r13 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [53]),
        .Q(\u1/uk/K_r13 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [54]),
        .Q(\u1/uk/K_r13 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [55]),
        .Q(\u1/uk/K_r13 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [5]),
        .Q(\u1/uk/K_r13 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [6]),
        .Q(\u1/uk/K_r13 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [7]),
        .Q(\u1/uk/K_r13 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [8]),
        .Q(\u1/uk/K_r13 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r13_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r12 [9]),
        .Q(\u1/uk/K_r13 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [0]),
        .Q(\u1/uk/K_r14_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [10]),
        .Q(\u1/uk/K_r14_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [11]),
        .Q(\u1/uk/K_r14_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [12]),
        .Q(\u1/uk/K_r14_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [13]),
        .Q(\u1/uk/K_r14_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [14]),
        .Q(\u1/uk/K_r14_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [15]),
        .Q(\u1/uk/K_r14_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [16]),
        .Q(\u1/uk/K_r14_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [17]),
        .Q(\u1/uk/K_r14_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [18]),
        .Q(\u1/uk/K_r14_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [19]),
        .Q(\u1/uk/K_r14_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [1]),
        .Q(\u1/uk/K_r14_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [20]),
        .Q(\u1/uk/K_r14_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [21]),
        .Q(\u1/uk/K_r14_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [22]),
        .Q(\u1/uk/K_r14_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [23]),
        .Q(\u1/uk/K_r14_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [24]),
        .Q(\u1/uk/K_r14_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [25]),
        .Q(\u1/uk/K_r14_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [26]),
        .Q(\u1/uk/K_r14_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [27]),
        .Q(\u1/uk/K_r14_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [28]),
        .Q(\u1/uk/K_r14_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [29]),
        .Q(\u1/uk/K_r14_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [2]),
        .Q(\u1/uk/K_r14_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [30]),
        .Q(\u1/uk/K_r14_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [31]),
        .Q(\u1/uk/K_r14_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [32]),
        .Q(\u1/uk/K_r14_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [33]),
        .Q(\u1/uk/K_r14_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [34]),
        .Q(\u1/uk/K_r14_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [35]),
        .Q(\u1/uk/K_r14_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [36]),
        .Q(\u1/uk/K_r14_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [37]),
        .Q(\u1/uk/K_r14_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [38]),
        .Q(\u1/uk/K_r14_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [39]),
        .Q(\u1/uk/K_r14_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [3]),
        .Q(\u1/uk/K_r14_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [40]),
        .Q(\u1/uk/K_r14_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [41]),
        .Q(\u1/uk/K_r14_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [42]),
        .Q(\u1/uk/K_r14_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [43]),
        .Q(\u1/uk/K_r14_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [44]),
        .Q(\u1/uk/K_r14_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [45]),
        .Q(\u1/uk/K_r14_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [46]),
        .Q(\u1/uk/K_r14_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [47]),
        .Q(\u1/uk/K_r14_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [48]),
        .Q(\u1/uk/K_r14_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [49]),
        .Q(\u1/uk/K_r14_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [4]),
        .Q(\u1/uk/K_r14_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [50]),
        .Q(\u1/uk/K_r14_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [51]),
        .Q(\u1/uk/K_r14_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [52]),
        .Q(\u1/uk/K_r14_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [53]),
        .Q(\u1/uk/K_r14_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [54]),
        .Q(\u1/uk/K_r14_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [55]),
        .Q(\u1/uk/K_r14_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [5]),
        .Q(\u1/uk/K_r14_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [6]),
        .Q(\u1/uk/K_r14_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [7]),
        .Q(\u1/uk/K_r14_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [8]),
        .Q(\u1/uk/K_r14_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r14_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r13 [9]),
        .Q(\u1/uk/K_r14_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_ ),
        .Q(\u1/uk/K_r1 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_0_in ),
        .Q(\u1/uk/K_r1 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_14_in ),
        .Q(\u1/uk/K_r1 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_38_in ),
        .Q(\u1/uk/K_r1 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_7_in ),
        .Q(\u1/uk/K_r1 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_36_in ),
        .Q(\u1/uk/K_r1 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_25_in ),
        .Q(\u1/uk/K_r1 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_27_in ),
        .Q(\u1/uk/K_r1 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[17] ),
        .Q(\u1/uk/K_r1 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_37_in ),
        .Q(\u1/uk/K_r1 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[19] ),
        .Q(\u1/uk/K_r1 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[1] ),
        .Q(\u1/uk/K_r1 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_2_in ),
        .Q(\u1/uk/K_r1 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_24_in ),
        .Q(\u1/uk/K_r1 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[22] ),
        .Q(\u1/uk/K_r1 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_30_in ),
        .Q(\u1/uk/K_r1 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_3_in ),
        .Q(\u1/uk/K_r1 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[25] ),
        .Q(\u1/uk/K_r1 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_9_in ),
        .Q(\u1/uk/K_r1 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_5_in ),
        .Q(\u1/uk/K_r1 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_20_in ),
        .Q(\u1/uk/K_r1 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_31_in ),
        .Q(\u1/uk/K_r1 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[2] ),
        .Q(\u1/uk/K_r1 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_22_in ),
        .Q(\u1/uk/K_r1 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[31] ),
        .Q(\u1/uk/K_r1 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[32] ),
        .Q(\u1/uk/K_r1 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_39_in ),
        .Q(\u1/uk/K_r1 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_6_in ),
        .Q(\u1/uk/K_r1 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[35] ),
        .Q(\u1/uk/K_r1 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[36] ),
        .Q(\u1/uk/K_r1 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_26_in ),
        .Q(\u1/uk/K_r1 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_18_in ),
        .Q(\u1/uk/K_r1 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_12_in ),
        .Q(\u1/uk/K_r1 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_11_in ),
        .Q(\u1/uk/K_r1 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_8_in ),
        .Q(\u1/uk/K_r1 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_13_in ),
        .Q(\u1/uk/K_r1 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_29_in ),
        .Q(\u1/uk/K_r1 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_17_in ),
        .Q(\u1/uk/K_r1 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_19_in ),
        .Q(\u1/uk/K_r1 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_33_in ),
        .Q(\u1/uk/K_r1 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_1_in ),
        .Q(\u1/uk/K_r1 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_15_in ),
        .Q(\u1/uk/K_r1 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_4_in ),
        .Q(\u1/uk/K_r1 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_34_in ),
        .Q(\u1/uk/K_r1 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[4] ),
        .Q(\u1/uk/K_r1 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_28_in ),
        .Q(\u1/uk/K_r1 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_35_in ),
        .Q(\u1/uk/K_r1 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[52] ),
        .Q(\u1/uk/K_r1 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[53] ),
        .Q(\u1/uk/K_r1 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_40_in ),
        .Q(\u1/uk/K_r1 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r0_reg_n_0_[55] ),
        .Q(\u1/uk/K_r1 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_10_in ),
        .Q(\u1/uk/K_r1 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_16_in ),
        .Q(\u1/uk/K_r1 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_21_in ),
        .Q(\u1/uk/K_r1 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_32_in ),
        .Q(\u1/uk/K_r1 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_23_in ),
        .Q(\u1/uk/K_r1 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [0]),
        .Q(\u1/uk/K_r2 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [10]),
        .Q(\u1/uk/K_r2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [11]),
        .Q(\u1/uk/K_r2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [12]),
        .Q(\u1/uk/K_r2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [13]),
        .Q(\u1/uk/K_r2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [14]),
        .Q(\u1/uk/K_r2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [15]),
        .Q(\u1/uk/K_r2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [16]),
        .Q(\u1/uk/K_r2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [17]),
        .Q(\u1/uk/K_r2 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [18]),
        .Q(\u1/uk/K_r2 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [19]),
        .Q(\u1/uk/K_r2 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [1]),
        .Q(\u1/uk/K_r2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [20]),
        .Q(\u1/uk/K_r2 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [21]),
        .Q(\u1/uk/K_r2 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [22]),
        .Q(\u1/uk/K_r2 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [23]),
        .Q(\u1/uk/K_r2 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [24]),
        .Q(\u1/uk/K_r2 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [25]),
        .Q(\u1/uk/K_r2 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [26]),
        .Q(\u1/uk/K_r2 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [27]),
        .Q(\u1/uk/K_r2 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [28]),
        .Q(\u1/uk/K_r2 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [29]),
        .Q(\u1/uk/K_r2 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [2]),
        .Q(\u1/uk/K_r2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [30]),
        .Q(\u1/uk/K_r2 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [31]),
        .Q(\u1/uk/K_r2 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [32]),
        .Q(\u1/uk/K_r2 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [33]),
        .Q(\u1/uk/K_r2 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [34]),
        .Q(\u1/uk/K_r2 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [35]),
        .Q(\u1/uk/K_r2 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [36]),
        .Q(\u1/uk/K_r2 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [37]),
        .Q(\u1/uk/K_r2 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [38]),
        .Q(\u1/uk/K_r2 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [39]),
        .Q(\u1/uk/K_r2 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [3]),
        .Q(\u1/uk/K_r2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [40]),
        .Q(\u1/uk/K_r2 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [41]),
        .Q(\u1/uk/K_r2 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [42]),
        .Q(\u1/uk/K_r2 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [43]),
        .Q(\u1/uk/K_r2 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [44]),
        .Q(\u1/uk/K_r2 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [45]),
        .Q(\u1/uk/K_r2 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [46]),
        .Q(\u1/uk/K_r2 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [47]),
        .Q(\u1/uk/K_r2 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [48]),
        .Q(\u1/uk/K_r2 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [49]),
        .Q(\u1/uk/K_r2 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [4]),
        .Q(\u1/uk/K_r2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [50]),
        .Q(\u1/uk/K_r2 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [51]),
        .Q(\u1/uk/K_r2 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [52]),
        .Q(\u1/uk/K_r2 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [53]),
        .Q(\u1/uk/K_r2 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [54]),
        .Q(\u1/uk/K_r2 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [55]),
        .Q(\u1/uk/K_r2 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [5]),
        .Q(\u1/uk/K_r2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [6]),
        .Q(\u1/uk/K_r2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [7]),
        .Q(\u1/uk/K_r2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [8]),
        .Q(\u1/uk/K_r2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r2_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r1 [9]),
        .Q(\u1/uk/K_r2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [0]),
        .Q(\u1/uk/K_r3 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [10]),
        .Q(\u1/uk/K_r3 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [11]),
        .Q(\u1/uk/K_r3 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [12]),
        .Q(\u1/uk/K_r3 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [13]),
        .Q(\u1/uk/K_r3 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [14]),
        .Q(\u1/uk/K_r3 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [15]),
        .Q(\u1/uk/K_r3 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [16]),
        .Q(\u1/uk/K_r3 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [17]),
        .Q(\u1/uk/K_r3 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [18]),
        .Q(\u1/uk/K_r3 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [19]),
        .Q(\u1/uk/K_r3 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [1]),
        .Q(\u1/uk/K_r3 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [20]),
        .Q(\u1/uk/K_r3 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [21]),
        .Q(\u1/uk/K_r3 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [22]),
        .Q(\u1/uk/K_r3 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [23]),
        .Q(\u1/uk/K_r3 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [24]),
        .Q(\u1/uk/K_r3 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [25]),
        .Q(\u1/uk/K_r3 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [26]),
        .Q(\u1/uk/K_r3 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [27]),
        .Q(\u1/uk/K_r3 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [28]),
        .Q(\u1/uk/K_r3 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [29]),
        .Q(\u1/uk/K_r3 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [2]),
        .Q(\u1/uk/K_r3 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [30]),
        .Q(\u1/uk/K_r3 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [31]),
        .Q(\u1/uk/K_r3 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [32]),
        .Q(\u1/uk/K_r3 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [33]),
        .Q(\u1/uk/K_r3 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [34]),
        .Q(\u1/uk/K_r3 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [35]),
        .Q(\u1/uk/K_r3 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [36]),
        .Q(\u1/uk/K_r3 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [37]),
        .Q(\u1/uk/K_r3 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [38]),
        .Q(\u1/uk/K_r3 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [39]),
        .Q(\u1/uk/K_r3 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [3]),
        .Q(\u1/uk/K_r3 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [40]),
        .Q(\u1/uk/K_r3 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [41]),
        .Q(\u1/uk/K_r3 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [42]),
        .Q(\u1/uk/K_r3 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [43]),
        .Q(\u1/uk/K_r3 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [44]),
        .Q(\u1/uk/K_r3 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [45]),
        .Q(\u1/uk/K_r3 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [46]),
        .Q(\u1/uk/K_r3 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [47]),
        .Q(\u1/uk/K_r3 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [48]),
        .Q(\u1/uk/K_r3 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [49]),
        .Q(\u1/uk/K_r3 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [4]),
        .Q(\u1/uk/K_r3 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [50]),
        .Q(\u1/uk/K_r3 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [51]),
        .Q(\u1/uk/K_r3 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [52]),
        .Q(\u1/uk/K_r3 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [53]),
        .Q(\u1/uk/K_r3 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [54]),
        .Q(\u1/uk/K_r3 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [55]),
        .Q(\u1/uk/K_r3 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [5]),
        .Q(\u1/uk/K_r3 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [6]),
        .Q(\u1/uk/K_r3 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [7]),
        .Q(\u1/uk/K_r3 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [8]),
        .Q(\u1/uk/K_r3 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r3_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r2 [9]),
        .Q(\u1/uk/K_r3 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [0]),
        .Q(\u1/uk/K_r4_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [10]),
        .Q(\u1/uk/K_r4_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [11]),
        .Q(\u1/uk/K_r4_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [12]),
        .Q(\u1/uk/K_r4_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [13]),
        .Q(\u1/uk/K_r4_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [14]),
        .Q(\u1/uk/K_r4_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [15]),
        .Q(\u1/uk/K_r4_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [16]),
        .Q(\u1/uk/K_r4_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [17]),
        .Q(\u1/uk/K_r4_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [18]),
        .Q(\u1/uk/K_r4_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [19]),
        .Q(\u1/uk/K_r4_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [1]),
        .Q(\u1/uk/K_r4_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [20]),
        .Q(\u1/uk/K_r4_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [21]),
        .Q(\u1/uk/K_r4_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [22]),
        .Q(\u1/uk/K_r4_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [23]),
        .Q(\u1/uk/K_r4_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [24]),
        .Q(\u1/uk/K_r4_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [25]),
        .Q(\u1/uk/K_r4_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [26]),
        .Q(\u1/uk/K_r4_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [27]),
        .Q(\u1/uk/K_r4_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [28]),
        .Q(\u1/uk/K_r4_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [29]),
        .Q(\u1/uk/K_r4_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [2]),
        .Q(\u1/uk/K_r4_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [30]),
        .Q(\u1/uk/K_r4_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [31]),
        .Q(\u1/uk/K_r4_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [32]),
        .Q(\u1/uk/K_r4_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [33]),
        .Q(\u1/uk/K_r4_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [34]),
        .Q(\u1/uk/p_50_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [35]),
        .Q(\u1/uk/K_r4_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [36]),
        .Q(\u1/uk/K_r4_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [37]),
        .Q(\u1/uk/K_r4_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [38]),
        .Q(\u1/uk/K_r4_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [39]),
        .Q(\u1/uk/K_r4_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [3]),
        .Q(\u1/uk/K_r4_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [40]),
        .Q(\u1/uk/p_49_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [41]),
        .Q(\u1/uk/K_r4_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [42]),
        .Q(\u1/uk/K_r4_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [43]),
        .Q(\u1/uk/p_44_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [44]),
        .Q(\u1/uk/K_r4_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [45]),
        .Q(\u1/uk/K_r4_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [46]),
        .Q(\u1/uk/p_47_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [47]),
        .Q(\u1/uk/K_r4_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [48]),
        .Q(\u1/uk/K_r4_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [49]),
        .Q(\u1/uk/K_r4_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [4]),
        .Q(\u1/uk/K_r4_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [50]),
        .Q(\u1/uk/K_r4_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [51]),
        .Q(\u1/uk/K_r4_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [52]),
        .Q(\u1/uk/K_r4_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [53]),
        .Q(\u1/uk/p_51_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [54]),
        .Q(\u1/uk/K_r4_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [55]),
        .Q(\u1/uk/K_r4_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [5]),
        .Q(\u1/uk/K_r4_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [6]),
        .Q(\u1/uk/K_r4_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [7]),
        .Q(\u1/uk/K_r4_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [8]),
        .Q(\u1/uk/p_42_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r4_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r3 [9]),
        .Q(\u1/uk/K_r4_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_ ),
        .Q(\u1/uk/K_r5 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[10] ),
        .Q(\u1/uk/K_r5 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[11] ),
        .Q(\u1/uk/K_r5 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[12] ),
        .Q(\u1/uk/K_r5 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[13] ),
        .Q(\u1/uk/K_r5 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[14] ),
        .Q(\u1/uk/K_r5 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[15] ),
        .Q(\u1/uk/K_r5 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[16] ),
        .Q(\u1/uk/K_r5 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[17] ),
        .Q(\u1/uk/K_r5 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[18] ),
        .Q(\u1/uk/K_r5 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[19] ),
        .Q(\u1/uk/K_r5 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[1] ),
        .Q(\u1/uk/K_r5 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[20] ),
        .Q(\u1/uk/K_r5 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[21] ),
        .Q(\u1/uk/K_r5 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[22] ),
        .Q(\u1/uk/K_r5 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[23] ),
        .Q(\u1/uk/K_r5 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[24] ),
        .Q(\u1/uk/K_r5 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[25] ),
        .Q(\u1/uk/K_r5 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[26] ),
        .Q(\u1/uk/K_r5 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[27] ),
        .Q(\u1/uk/K_r5 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[28] ),
        .Q(\u1/uk/K_r5 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[29] ),
        .Q(\u1/uk/K_r5 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[2] ),
        .Q(\u1/uk/K_r5 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[30] ),
        .Q(\u1/uk/K_r5 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[31] ),
        .Q(\u1/uk/K_r5 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[32] ),
        .Q(\u1/uk/K_r5 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[33] ),
        .Q(\u1/uk/K_r5 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_50_in ),
        .Q(\u1/uk/K_r5 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[35] ),
        .Q(\u1/uk/K_r5 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[36] ),
        .Q(\u1/uk/K_r5 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[37] ),
        .Q(\u1/uk/K_r5 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[38] ),
        .Q(\u1/uk/K_r5 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[39] ),
        .Q(\u1/uk/K_r5 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[3] ),
        .Q(\u1/uk/K_r5 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_49_in ),
        .Q(\u1/uk/K_r5 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[41] ),
        .Q(\u1/uk/K_r5 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[42] ),
        .Q(\u1/uk/K_r5 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_44_in ),
        .Q(\u1/uk/K_r5 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[44] ),
        .Q(\u1/uk/K_r5 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[45] ),
        .Q(\u1/uk/K_r5 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_47_in ),
        .Q(\u1/uk/K_r5 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[47] ),
        .Q(\u1/uk/K_r5 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[48] ),
        .Q(\u1/uk/K_r5 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[49] ),
        .Q(\u1/uk/K_r5 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[4] ),
        .Q(\u1/uk/K_r5 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[50] ),
        .Q(\u1/uk/K_r5 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[51] ),
        .Q(\u1/uk/K_r5 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[52] ),
        .Q(\u1/uk/K_r5 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_51_in ),
        .Q(\u1/uk/K_r5 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[54] ),
        .Q(\u1/uk/K_r5 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[55] ),
        .Q(\u1/uk/K_r5 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[5] ),
        .Q(\u1/uk/K_r5 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[6] ),
        .Q(\u1/uk/K_r5 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[7] ),
        .Q(\u1/uk/K_r5 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_42_in ),
        .Q(\u1/uk/K_r5 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r5_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r4_reg_n_0_[9] ),
        .Q(\u1/uk/K_r5 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [0]),
        .Q(\u1/uk/K_r6_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [10]),
        .Q(\u1/uk/K_r6_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [11]),
        .Q(\u1/uk/K_r6_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [12]),
        .Q(\u1/uk/K_r6_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [13]),
        .Q(\u1/uk/p_52_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [14]),
        .Q(\u1/uk/K_r6_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [15]),
        .Q(\u1/uk/K_r6_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [16]),
        .Q(\u1/uk/K_r6_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [17]),
        .Q(\u1/uk/K_r6_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [18]),
        .Q(\u1/uk/K_r6_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [19]),
        .Q(\u1/uk/K_r6_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [1]),
        .Q(\u1/uk/K_r6_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [20]),
        .Q(\u1/uk/K_r6_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [21]),
        .Q(\u1/uk/K_r6_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [22]),
        .Q(\u1/uk/K_r6_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [23]),
        .Q(\u1/uk/K_r6_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [24]),
        .Q(\u1/uk/K_r6_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [25]),
        .Q(\u1/uk/K_r6_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [26]),
        .Q(\u1/uk/K_r6_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [27]),
        .Q(\u1/uk/K_r6_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [28]),
        .Q(\u1/uk/K_r6_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [29]),
        .Q(\u1/uk/K_r6_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [2]),
        .Q(\u1/uk/K_r6_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [30]),
        .Q(\u1/uk/K_r6_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [31]),
        .Q(\u1/uk/K_r6_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [32]),
        .Q(\u1/uk/K_r6_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [33]),
        .Q(\u1/uk/K_r6_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [34]),
        .Q(\u1/uk/K_r6_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [35]),
        .Q(\u1/uk/K_r6_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [36]),
        .Q(\u1/uk/K_r6_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [37]),
        .Q(\u1/uk/K_r6_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [38]),
        .Q(\u1/uk/K_r6_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [39]),
        .Q(\u1/uk/K_r6_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [3]),
        .Q(\u1/uk/K_r6_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [40]),
        .Q(\u1/uk/K_r6_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [41]),
        .Q(\u1/uk/K_r6_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [42]),
        .Q(\u1/uk/p_41_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [43]),
        .Q(\u1/uk/p_45_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [44]),
        .Q(\u1/uk/K_r6_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [45]),
        .Q(\u1/uk/K_r6_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [46]),
        .Q(\u1/uk/K_r6_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [47]),
        .Q(\u1/uk/K_r6_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [48]),
        .Q(\u1/uk/K_r6_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [49]),
        .Q(\u1/uk/p_43_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [4]),
        .Q(\u1/uk/K_r6_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [50]),
        .Q(\u1/uk/K_r6_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [51]),
        .Q(\u1/uk/K_r6_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [52]),
        .Q(\u1/uk/K_r6_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [53]),
        .Q(\u1/uk/K_r6_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [54]),
        .Q(\u1/uk/K_r6_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [55]),
        .Q(\u1/uk/K_r6_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [5]),
        .Q(\u1/uk/K_r6_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [6]),
        .Q(\u1/uk/p_53_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [7]),
        .Q(\u1/uk/K_r6_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [8]),
        .Q(\u1/uk/K_r6_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r6_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r5 [9]),
        .Q(\u1/uk/K_r6_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_ ),
        .Q(\u1/uk/K_r7_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[10] ),
        .Q(\u1/uk/K_r7_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[11] ),
        .Q(\u1/uk/K_r7_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[12] ),
        .Q(\u1/uk/K_r7_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_52_in ),
        .Q(\u1/uk/K_r7_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[14] ),
        .Q(\u1/uk/K_r7_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[15] ),
        .Q(\u1/uk/K_r7_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[16] ),
        .Q(\u1/uk/K_r7_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[17] ),
        .Q(\u1/uk/K_r7_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[18] ),
        .Q(\u1/uk/K_r7_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[19] ),
        .Q(\u1/uk/K_r7_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[1] ),
        .Q(\u1/uk/K_r7_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[20] ),
        .Q(\u1/uk/K_r7_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[21] ),
        .Q(\u1/uk/K_r7_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[22] ),
        .Q(\u1/uk/K_r7_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[23] ),
        .Q(\u1/uk/K_r7_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[24] ),
        .Q(\u1/uk/K_r7_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[25] ),
        .Q(\u1/uk/K_r7_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[26] ),
        .Q(\u1/uk/K_r7_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[27] ),
        .Q(\u1/uk/K_r7_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[28] ),
        .Q(\u1/uk/K_r7_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[29] ),
        .Q(\u1/uk/K_r7_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[2] ),
        .Q(\u1/uk/K_r7_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[30] ),
        .Q(\u1/uk/K_r7_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[31] ),
        .Q(\u1/uk/K_r7_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[32] ),
        .Q(\u1/uk/K_r7_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[33] ),
        .Q(\u1/uk/K_r7_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[34] ),
        .Q(\u1/uk/K_r7_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[35] ),
        .Q(\u1/uk/K_r7_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[36] ),
        .Q(\u1/uk/K_r7_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[37] ),
        .Q(\u1/uk/K_r7_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[38] ),
        .Q(\u1/uk/K_r7_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[39] ),
        .Q(\u1/uk/K_r7_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[3] ),
        .Q(\u1/uk/K_r7_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[40] ),
        .Q(\u1/uk/K_r7_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[41] ),
        .Q(\u1/uk/K_r7_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_41_in ),
        .Q(\u1/uk/K_r7_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_45_in ),
        .Q(\u1/uk/K_r7_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[44] ),
        .Q(\u1/uk/p_48_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[45] ),
        .Q(\u1/uk/K_r7_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[46] ),
        .Q(\u1/uk/K_r7_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[47] ),
        .Q(\u1/uk/K_r7_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[48] ),
        .Q(\u1/uk/K_r7_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_43_in ),
        .Q(\u1/uk/K_r7_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[4] ),
        .Q(\u1/uk/K_r7_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[50] ),
        .Q(\u1/uk/K_r7_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[51] ),
        .Q(\u1/uk/K_r7_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[52] ),
        .Q(\u1/uk/K_r7_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[53] ),
        .Q(\u1/uk/K_r7_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[54] ),
        .Q(\u1/uk/K_r7_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[55] ),
        .Q(\u1/uk/K_r7_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[5] ),
        .Q(\u1/uk/K_r7_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_53_in ),
        .Q(\u1/uk/K_r7_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[7] ),
        .Q(\u1/uk/K_r7_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[8] ),
        .Q(\u1/uk/K_r7_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r7_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r6_reg_n_0_[9] ),
        .Q(\u1/uk/K_r7_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_ ),
        .Q(\u1/uk/K_r8 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[10] ),
        .Q(\u1/uk/K_r8 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[11] ),
        .Q(\u1/uk/K_r8 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[12] ),
        .Q(\u1/uk/K_r8 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[13] ),
        .Q(\u1/uk/K_r8 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[14] ),
        .Q(\u1/uk/K_r8 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[15] ),
        .Q(\u1/uk/K_r8 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[16] ),
        .Q(\u1/uk/K_r8 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[17] ),
        .Q(\u1/uk/K_r8 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[18] ),
        .Q(\u1/uk/K_r8 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[19] ),
        .Q(\u1/uk/K_r8 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[1] ),
        .Q(\u1/uk/K_r8 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[20] ),
        .Q(\u1/uk/K_r8 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[21] ),
        .Q(\u1/uk/K_r8 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[22] ),
        .Q(\u1/uk/K_r8 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[23] ),
        .Q(\u1/uk/K_r8 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[24] ),
        .Q(\u1/uk/K_r8 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[25] ),
        .Q(\u1/uk/K_r8 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[26] ),
        .Q(\u1/uk/K_r8 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[27] ),
        .Q(\u1/uk/K_r8 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[28] ),
        .Q(\u1/uk/K_r8 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[29] ),
        .Q(\u1/uk/K_r8 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[2] ),
        .Q(\u1/uk/K_r8 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[30] ),
        .Q(\u1/uk/K_r8 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[31] ),
        .Q(\u1/uk/K_r8 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[32] ),
        .Q(\u1/uk/K_r8 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[33] ),
        .Q(\u1/uk/K_r8 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[34] ),
        .Q(\u1/uk/K_r8 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[35] ),
        .Q(\u1/uk/K_r8 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[36] ),
        .Q(\u1/uk/K_r8 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[37] ),
        .Q(\u1/uk/K_r8 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[38] ),
        .Q(\u1/uk/K_r8 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[39] ),
        .Q(\u1/uk/K_r8 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[3] ),
        .Q(\u1/uk/K_r8 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[40] ),
        .Q(\u1/uk/K_r8 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[41] ),
        .Q(\u1/uk/K_r8 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[42] ),
        .Q(\u1/uk/K_r8 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[43] ),
        .Q(\u1/uk/K_r8 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/p_48_in ),
        .Q(\u1/uk/K_r8 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[45] ),
        .Q(\u1/uk/K_r8 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[46] ),
        .Q(\u1/uk/K_r8 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[47] ),
        .Q(\u1/uk/K_r8 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[48] ),
        .Q(\u1/uk/K_r8 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[49] ),
        .Q(\u1/uk/K_r8 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[4] ),
        .Q(\u1/uk/K_r8 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[50] ),
        .Q(\u1/uk/K_r8 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[51] ),
        .Q(\u1/uk/K_r8 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[52] ),
        .Q(\u1/uk/K_r8 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[53] ),
        .Q(\u1/uk/K_r8 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[54] ),
        .Q(\u1/uk/K_r8 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[55] ),
        .Q(\u1/uk/K_r8 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[5] ),
        .Q(\u1/uk/K_r8 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[6] ),
        .Q(\u1/uk/K_r8 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[7] ),
        .Q(\u1/uk/K_r8 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[8] ),
        .Q(\u1/uk/K_r8 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r8_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r7_reg_n_0_[9] ),
        .Q(\u1/uk/K_r8 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [0]),
        .Q(\u1/uk/K_r9 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [10]),
        .Q(\u1/uk/K_r9 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [11]),
        .Q(\u1/uk/K_r9 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [12]),
        .Q(\u1/uk/K_r9 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [13]),
        .Q(\u1/uk/K_r9 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [14]),
        .Q(\u1/uk/K_r9 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [15]),
        .Q(\u1/uk/K_r9 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [16]),
        .Q(\u1/uk/K_r9 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [17]),
        .Q(\u1/uk/K_r9 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [18]),
        .Q(\u1/uk/K_r9 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [19]),
        .Q(\u1/uk/K_r9 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [1]),
        .Q(\u1/uk/K_r9 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [20]),
        .Q(\u1/uk/K_r9 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [21]),
        .Q(\u1/uk/K_r9 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [22]),
        .Q(\u1/uk/K_r9 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [23]),
        .Q(\u1/uk/K_r9 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [24]),
        .Q(\u1/uk/K_r9 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [25]),
        .Q(\u1/uk/K_r9 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [26]),
        .Q(\u1/uk/K_r9 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [27]),
        .Q(\u1/uk/K_r9 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [28]),
        .Q(\u1/uk/K_r9 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [29]),
        .Q(\u1/uk/K_r9 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [2]),
        .Q(\u1/uk/K_r9 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [30]),
        .Q(\u1/uk/K_r9 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [31]),
        .Q(\u1/uk/K_r9 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [32]),
        .Q(\u1/uk/K_r9 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [33]),
        .Q(\u1/uk/K_r9 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [34]),
        .Q(\u1/uk/K_r9 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [35]),
        .Q(\u1/uk/K_r9 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [36]),
        .Q(\u1/uk/K_r9 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [37]),
        .Q(\u1/uk/K_r9 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [38]),
        .Q(\u1/uk/K_r9 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [39]),
        .Q(\u1/uk/K_r9 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [3]),
        .Q(\u1/uk/K_r9 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [40]),
        .Q(\u1/uk/K_r9 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [41]),
        .Q(\u1/uk/K_r9 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [42]),
        .Q(\u1/uk/K_r9 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [43]),
        .Q(\u1/uk/K_r9 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [44]),
        .Q(\u1/uk/K_r9 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [45]),
        .Q(\u1/uk/K_r9 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [46]),
        .Q(\u1/uk/K_r9 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [47]),
        .Q(\u1/uk/K_r9 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [48]),
        .Q(\u1/uk/K_r9 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [49]),
        .Q(\u1/uk/K_r9 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [4]),
        .Q(\u1/uk/K_r9 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [50]),
        .Q(\u1/uk/K_r9 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [51]),
        .Q(\u1/uk/K_r9 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [52]),
        .Q(\u1/uk/K_r9 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [53]),
        .Q(\u1/uk/K_r9 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [54]),
        .Q(\u1/uk/K_r9 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [55]),
        .Q(\u1/uk/K_r9 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [5]),
        .Q(\u1/uk/K_r9 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [6]),
        .Q(\u1/uk/K_r9 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [7]),
        .Q(\u1/uk/K_r9 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [8]),
        .Q(\u1/uk/K_r9 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u1/uk/K_r9_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u1/uk/K_r8 [9]),
        .Q(\u1/uk/K_r9 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [42]),
        .Q(\u2/L0 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [43]),
        .Q(\u2/L0 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [44]),
        .Q(\u2/L0 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [45]),
        .Q(\u2/L0 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [46]),
        .Q(\u2/L0 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [47]),
        .Q(\u2/L0 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [48]),
        .Q(\u2/L0 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [49]),
        .Q(\u2/L0 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [50]),
        .Q(\u2/L0 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [51]),
        .Q(\u2/L0 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [33]),
        .Q(\u2/L0 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [52]),
        .Q(\u2/L0 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [53]),
        .Q(\u2/L0 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [54]),
        .Q(\u2/L0 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [55]),
        .Q(\u2/L0 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [56]),
        .Q(\u2/L0 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [57]),
        .Q(\u2/L0 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [58]),
        .Q(\u2/L0 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [59]),
        .Q(\u2/L0 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [60]),
        .Q(\u2/L0 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [61]),
        .Q(\u2/L0 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [34]),
        .Q(\u2/L0 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [62]),
        .Q(\u2/L0 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [63]),
        .Q(\u2/L0 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [64]),
        .Q(\u2/L0 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [35]),
        .Q(\u2/L0 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [36]),
        .Q(\u2/L0 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [37]),
        .Q(\u2/L0 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [38]),
        .Q(\u2/L0 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [39]),
        .Q(\u2/L0 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [40]),
        .Q(\u2/L0 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L0_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/IP [41]),
        .Q(\u2/L0 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [10]),
        .Q(\u2/L10 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [11]),
        .Q(\u2/L10 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [12]),
        .Q(\u2/L10 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [13]),
        .Q(\u2/L10 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [14]),
        .Q(\u2/L10 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [15]),
        .Q(\u2/L10 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [16]),
        .Q(\u2/L10 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [17]),
        .Q(\u2/L10 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [18]),
        .Q(\u2/L10 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [19]),
        .Q(\u2/L10 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [1]),
        .Q(\u2/L10 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [20]),
        .Q(\u2/L10 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [21]),
        .Q(\u2/L10 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [22]),
        .Q(\u2/L10 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [23]),
        .Q(\u2/L10 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [24]),
        .Q(\u2/L10 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [25]),
        .Q(\u2/L10 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [26]),
        .Q(\u2/L10 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [27]),
        .Q(\u2/L10 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [28]),
        .Q(\u2/L10 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [29]),
        .Q(\u2/L10 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [2]),
        .Q(\u2/L10 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [30]),
        .Q(\u2/L10 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [31]),
        .Q(\u2/L10 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [32]),
        .Q(\u2/L10 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [3]),
        .Q(\u2/L10 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [4]),
        .Q(\u2/L10 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [5]),
        .Q(\u2/L10 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [6]),
        .Q(\u2/L10 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [7]),
        .Q(\u2/L10 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [8]),
        .Q(\u2/L10 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L10_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R9 [9]),
        .Q(\u2/L10 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_ ),
        .Q(\u2/L11 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[11] ),
        .Q(\u2/L11 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[12] ),
        .Q(\u2/L11 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[13] ),
        .Q(\u2/L11 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[14] ),
        .Q(\u2/L11 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[15] ),
        .Q(\u2/L11 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[16] ),
        .Q(\u2/L11 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[17] ),
        .Q(\u2/L11 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[18] ),
        .Q(\u2/L11 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[19] ),
        .Q(\u2/L11 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[1] ),
        .Q(\u2/L11 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[20] ),
        .Q(\u2/L11 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[21] ),
        .Q(\u2/L11 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[22] ),
        .Q(\u2/L11 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[23] ),
        .Q(\u2/L11 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[24] ),
        .Q(\u2/L11 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[25] ),
        .Q(\u2/L11 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[26] ),
        .Q(\u2/L11 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[27] ),
        .Q(\u2/L11 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[28] ),
        .Q(\u2/L11 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[29] ),
        .Q(\u2/L11 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[2] ),
        .Q(\u2/L11 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[30] ),
        .Q(\u2/L11 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[31] ),
        .Q(\u2/L11 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[32] ),
        .Q(\u2/L11 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[3] ),
        .Q(\u2/L11 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[4] ),
        .Q(\u2/L11 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[5] ),
        .Q(\u2/L11 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[6] ),
        .Q(\u2/L11 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[7] ),
        .Q(\u2/L11 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[8] ),
        .Q(\u2/L11 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L11_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10_reg_n_0_[9] ),
        .Q(\u2/L11 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [10]),
        .Q(\u2/L12 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [11]),
        .Q(\u2/L12 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [12]),
        .Q(\u2/L12 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [13]),
        .Q(\u2/L12 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [14]),
        .Q(\u2/L12 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [15]),
        .Q(\u2/L12 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [16]),
        .Q(\u2/L12 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [17]),
        .Q(\u2/L12 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [18]),
        .Q(\u2/L12 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [19]),
        .Q(\u2/L12 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [1]),
        .Q(\u2/L12 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [20]),
        .Q(\u2/L12 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [21]),
        .Q(\u2/L12 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [22]),
        .Q(\u2/L12 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [23]),
        .Q(\u2/L12 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [24]),
        .Q(\u2/L12 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [25]),
        .Q(\u2/L12 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [26]),
        .Q(\u2/L12 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [27]),
        .Q(\u2/L12 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [28]),
        .Q(\u2/L12 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [29]),
        .Q(\u2/L12 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [2]),
        .Q(\u2/L12 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [30]),
        .Q(\u2/L12 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [31]),
        .Q(\u2/L12 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [32]),
        .Q(\u2/L12 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [3]),
        .Q(\u2/L12 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [4]),
        .Q(\u2/L12 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [5]),
        .Q(\u2/L12 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [6]),
        .Q(\u2/L12 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [7]),
        .Q(\u2/L12 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [8]),
        .Q(\u2/L12 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L12_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R11 [9]),
        .Q(\u2/L12 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [10]),
        .Q(\u2/L13 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [11]),
        .Q(\u2/L13 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [12]),
        .Q(\u2/L13 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [13]),
        .Q(\u2/L13 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [14]),
        .Q(\u2/L13 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [15]),
        .Q(\u2/L13 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [16]),
        .Q(\u2/L13 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [17]),
        .Q(\u2/L13 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [18]),
        .Q(\u2/L13 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [19]),
        .Q(\u2/L13 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [1]),
        .Q(\u2/L13 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [20]),
        .Q(\u2/L13 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [21]),
        .Q(\u2/L13 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [22]),
        .Q(\u2/L13 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [23]),
        .Q(\u2/L13 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [24]),
        .Q(\u2/L13 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [25]),
        .Q(\u2/L13 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [26]),
        .Q(\u2/L13 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [27]),
        .Q(\u2/L13 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [28]),
        .Q(\u2/L13 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [29]),
        .Q(\u2/L13 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [2]),
        .Q(\u2/L13 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [30]),
        .Q(\u2/L13 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [31]),
        .Q(\u2/L13 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [32]),
        .Q(\u2/L13 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [3]),
        .Q(\u2/L13 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [4]),
        .Q(\u2/L13 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [5]),
        .Q(\u2/L13 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [6]),
        .Q(\u2/L13 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [7]),
        .Q(\u2/L13 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [8]),
        .Q(\u2/L13 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L13_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R12 [9]),
        .Q(\u2/L13 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [10]),
        .Q(\u2/L14 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [11]),
        .Q(\u2/L14 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [12]),
        .Q(\u2/L14 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [13]),
        .Q(\u2/L14 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [14]),
        .Q(\u2/L14 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [15]),
        .Q(\u2/L14 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [16]),
        .Q(\u2/L14 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [17]),
        .Q(\u2/L14 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [18]),
        .Q(\u2/L14 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [19]),
        .Q(\u2/L14 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [1]),
        .Q(\u2/L14 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [20]),
        .Q(\u2/L14 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [21]),
        .Q(\u2/L14 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [22]),
        .Q(\u2/L14 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [23]),
        .Q(\u2/L14 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [24]),
        .Q(\u2/L14 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [25]),
        .Q(\u2/L14 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [26]),
        .Q(\u2/L14 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [27]),
        .Q(\u2/L14 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [28]),
        .Q(\u2/L14 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [29]),
        .Q(\u2/L14 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [2]),
        .Q(\u2/L14 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [30]),
        .Q(\u2/L14 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [31]),
        .Q(\u2/L14 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [32]),
        .Q(\u2/L14 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [3]),
        .Q(\u2/L14 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [4]),
        .Q(\u2/L14 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [5]),
        .Q(\u2/L14 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [6]),
        .Q(\u2/L14 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [7]),
        .Q(\u2/L14 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [8]),
        .Q(\u2/L14 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L14_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R13 [9]),
        .Q(\u2/L14 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [10]),
        .Q(\u2/L1 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [11]),
        .Q(\u2/L1 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [12]),
        .Q(\u2/L1 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [13]),
        .Q(\u2/L1 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [14]),
        .Q(\u2/L1 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [15]),
        .Q(\u2/L1 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [16]),
        .Q(\u2/L1 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [17]),
        .Q(\u2/L1 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [18]),
        .Q(\u2/L1 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [19]),
        .Q(\u2/L1 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [1]),
        .Q(\u2/L1 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [20]),
        .Q(\u2/L1 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [21]),
        .Q(\u2/L1 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [22]),
        .Q(\u2/L1 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [23]),
        .Q(\u2/L1 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [24]),
        .Q(\u2/L1 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [25]),
        .Q(\u2/L1 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [26]),
        .Q(\u2/L1 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [27]),
        .Q(\u2/L1 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [28]),
        .Q(\u2/L1 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [29]),
        .Q(\u2/L1 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [2]),
        .Q(\u2/L1 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [30]),
        .Q(\u2/L1 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [31]),
        .Q(\u2/L1 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [32]),
        .Q(\u2/L1 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [3]),
        .Q(\u2/L1 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [4]),
        .Q(\u2/L1 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [5]),
        .Q(\u2/L1 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [6]),
        .Q(\u2/L1 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [7]),
        .Q(\u2/L1 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [8]),
        .Q(\u2/L1 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R0 [9]),
        .Q(\u2/L1 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [10]),
        .Q(\u2/L2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [11]),
        .Q(\u2/L2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [12]),
        .Q(\u2/L2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [13]),
        .Q(\u2/L2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [14]),
        .Q(\u2/L2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [15]),
        .Q(\u2/L2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [16]),
        .Q(\u2/L2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [17]),
        .Q(\u2/L2 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [18]),
        .Q(\u2/L2 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [19]),
        .Q(\u2/L2 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [1]),
        .Q(\u2/L2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [20]),
        .Q(\u2/L2 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [21]),
        .Q(\u2/L2 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [22]),
        .Q(\u2/L2 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [23]),
        .Q(\u2/L2 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [24]),
        .Q(\u2/L2 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [25]),
        .Q(\u2/L2 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [26]),
        .Q(\u2/L2 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [27]),
        .Q(\u2/L2 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [28]),
        .Q(\u2/L2 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [29]),
        .Q(\u2/L2 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [2]),
        .Q(\u2/L2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [30]),
        .Q(\u2/L2 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [31]),
        .Q(\u2/L2 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [32]),
        .Q(\u2/L2 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [3]),
        .Q(\u2/L2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [4]),
        .Q(\u2/L2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [5]),
        .Q(\u2/L2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [6]),
        .Q(\u2/L2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [7]),
        .Q(\u2/L2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [8]),
        .Q(\u2/L2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L2_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R1 [9]),
        .Q(\u2/L2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [10]),
        .Q(\u2/L3 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [11]),
        .Q(\u2/L3 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [12]),
        .Q(\u2/L3 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [13]),
        .Q(\u2/L3 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [14]),
        .Q(\u2/L3 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [15]),
        .Q(\u2/L3 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [16]),
        .Q(\u2/L3 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [17]),
        .Q(\u2/L3 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [18]),
        .Q(\u2/L3 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [19]),
        .Q(\u2/L3 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [1]),
        .Q(\u2/L3 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [20]),
        .Q(\u2/L3 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [21]),
        .Q(\u2/L3 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [22]),
        .Q(\u2/L3 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [23]),
        .Q(\u2/L3 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [24]),
        .Q(\u2/L3 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [25]),
        .Q(\u2/L3 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [26]),
        .Q(\u2/L3 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [27]),
        .Q(\u2/L3 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [28]),
        .Q(\u2/L3 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [29]),
        .Q(\u2/L3 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [2]),
        .Q(\u2/L3 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [30]),
        .Q(\u2/L3 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [31]),
        .Q(\u2/L3 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [32]),
        .Q(\u2/L3 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [3]),
        .Q(\u2/L3 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [4]),
        .Q(\u2/L3 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [5]),
        .Q(\u2/L3 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [6]),
        .Q(\u2/L3 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [7]),
        .Q(\u2/L3 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [8]),
        .Q(\u2/L3 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L3_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R2 [9]),
        .Q(\u2/L3 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [10]),
        .Q(\u2/L4 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [11]),
        .Q(\u2/L4 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [12]),
        .Q(\u2/L4 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [13]),
        .Q(\u2/L4 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [14]),
        .Q(\u2/L4 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [15]),
        .Q(\u2/L4 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [16]),
        .Q(\u2/L4 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [17]),
        .Q(\u2/L4 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [18]),
        .Q(\u2/L4 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [19]),
        .Q(\u2/L4 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [1]),
        .Q(\u2/L4 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [20]),
        .Q(\u2/L4 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [21]),
        .Q(\u2/L4 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [22]),
        .Q(\u2/L4 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [23]),
        .Q(\u2/L4 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [24]),
        .Q(\u2/L4 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [25]),
        .Q(\u2/L4 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [26]),
        .Q(\u2/L4 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [27]),
        .Q(\u2/L4 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [28]),
        .Q(\u2/L4 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [29]),
        .Q(\u2/L4 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [2]),
        .Q(\u2/L4 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [30]),
        .Q(\u2/L4 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [31]),
        .Q(\u2/L4 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [32]),
        .Q(\u2/L4 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [3]),
        .Q(\u2/L4 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [4]),
        .Q(\u2/L4 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [5]),
        .Q(\u2/L4 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [6]),
        .Q(\u2/L4 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [7]),
        .Q(\u2/L4 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [8]),
        .Q(\u2/L4 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L4_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R3 [9]),
        .Q(\u2/L4 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [10]),
        .Q(\u2/L5 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [11]),
        .Q(\u2/L5 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [12]),
        .Q(\u2/L5 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [13]),
        .Q(\u2/L5 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [14]),
        .Q(\u2/L5 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [15]),
        .Q(\u2/L5 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [16]),
        .Q(\u2/L5 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [17]),
        .Q(\u2/L5 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [18]),
        .Q(\u2/L5 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [19]),
        .Q(\u2/L5 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [1]),
        .Q(\u2/L5 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [20]),
        .Q(\u2/L5 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [21]),
        .Q(\u2/L5 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [22]),
        .Q(\u2/L5 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [23]),
        .Q(\u2/L5 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [24]),
        .Q(\u2/L5 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [25]),
        .Q(\u2/L5 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [26]),
        .Q(\u2/L5 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [27]),
        .Q(\u2/L5 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [28]),
        .Q(\u2/L5 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [29]),
        .Q(\u2/L5 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [2]),
        .Q(\u2/L5 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [30]),
        .Q(\u2/L5 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [31]),
        .Q(\u2/L5 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [32]),
        .Q(\u2/L5 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [3]),
        .Q(\u2/L5 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [4]),
        .Q(\u2/L5 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [5]),
        .Q(\u2/L5 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [6]),
        .Q(\u2/L5 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [7]),
        .Q(\u2/L5 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [8]),
        .Q(\u2/L5 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L5_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R4 [9]),
        .Q(\u2/L5 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [10]),
        .Q(\u2/L6 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [11]),
        .Q(\u2/L6 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [12]),
        .Q(\u2/L6 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [13]),
        .Q(\u2/L6 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [14]),
        .Q(\u2/L6 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [15]),
        .Q(\u2/L6 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [16]),
        .Q(\u2/L6 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [17]),
        .Q(\u2/L6 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [18]),
        .Q(\u2/L6 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [19]),
        .Q(\u2/L6 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [1]),
        .Q(\u2/L6 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [20]),
        .Q(\u2/L6 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [21]),
        .Q(\u2/L6 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [22]),
        .Q(\u2/L6 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [23]),
        .Q(\u2/L6 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [24]),
        .Q(\u2/L6 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [25]),
        .Q(\u2/L6 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [26]),
        .Q(\u2/L6 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [27]),
        .Q(\u2/L6 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [28]),
        .Q(\u2/L6 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [29]),
        .Q(\u2/L6 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [2]),
        .Q(\u2/L6 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [30]),
        .Q(\u2/L6 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [31]),
        .Q(\u2/L6 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [32]),
        .Q(\u2/L6 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [3]),
        .Q(\u2/L6 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [4]),
        .Q(\u2/L6 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [5]),
        .Q(\u2/L6 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [6]),
        .Q(\u2/L6 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [7]),
        .Q(\u2/L6 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [8]),
        .Q(\u2/L6 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L6_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R5 [9]),
        .Q(\u2/L6 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [10]),
        .Q(\u2/L7 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [11]),
        .Q(\u2/L7 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [12]),
        .Q(\u2/L7 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [13]),
        .Q(\u2/L7 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [14]),
        .Q(\u2/L7 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [15]),
        .Q(\u2/L7 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [16]),
        .Q(\u2/L7 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [17]),
        .Q(\u2/L7 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [18]),
        .Q(\u2/L7 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [19]),
        .Q(\u2/L7 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [1]),
        .Q(\u2/L7 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [20]),
        .Q(\u2/L7 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [21]),
        .Q(\u2/L7 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [22]),
        .Q(\u2/L7 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [23]),
        .Q(\u2/L7 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [24]),
        .Q(\u2/L7 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [25]),
        .Q(\u2/L7 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [26]),
        .Q(\u2/L7 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [27]),
        .Q(\u2/L7 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [28]),
        .Q(\u2/L7 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [29]),
        .Q(\u2/L7 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [2]),
        .Q(\u2/L7 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [30]),
        .Q(\u2/L7 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [31]),
        .Q(\u2/L7 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [32]),
        .Q(\u2/L7 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [3]),
        .Q(\u2/L7 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [4]),
        .Q(\u2/L7 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [5]),
        .Q(\u2/L7 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [6]),
        .Q(\u2/L7 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [7]),
        .Q(\u2/L7 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [8]),
        .Q(\u2/L7 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L7_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R6 [9]),
        .Q(\u2/L7 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [10]),
        .Q(\u2/L8 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [11]),
        .Q(\u2/L8 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [12]),
        .Q(\u2/L8 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [13]),
        .Q(\u2/L8 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [14]),
        .Q(\u2/L8 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [15]),
        .Q(\u2/L8 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [16]),
        .Q(\u2/L8 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [17]),
        .Q(\u2/L8 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [18]),
        .Q(\u2/L8 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [19]),
        .Q(\u2/L8 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [1]),
        .Q(\u2/L8 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [20]),
        .Q(\u2/L8 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [21]),
        .Q(\u2/L8 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [22]),
        .Q(\u2/L8 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [23]),
        .Q(\u2/L8 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [24]),
        .Q(\u2/L8 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [25]),
        .Q(\u2/L8 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [26]),
        .Q(\u2/L8 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [27]),
        .Q(\u2/L8 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [28]),
        .Q(\u2/L8 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [29]),
        .Q(\u2/L8 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [2]),
        .Q(\u2/L8 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [30]),
        .Q(\u2/L8 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [31]),
        .Q(\u2/L8 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [32]),
        .Q(\u2/L8 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [3]),
        .Q(\u2/L8 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [4]),
        .Q(\u2/L8 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [5]),
        .Q(\u2/L8 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [6]),
        .Q(\u2/L8 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [7]),
        .Q(\u2/L8 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [8]),
        .Q(\u2/L8 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L8_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R7 [9]),
        .Q(\u2/L8 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [10]),
        .Q(\u2/L9 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [11]),
        .Q(\u2/L9 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [12]),
        .Q(\u2/L9 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [13]),
        .Q(\u2/L9 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [14]),
        .Q(\u2/L9 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [15]),
        .Q(\u2/L9 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [16]),
        .Q(\u2/L9 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [17]),
        .Q(\u2/L9 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [18]),
        .Q(\u2/L9 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [19]),
        .Q(\u2/L9 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [1]),
        .Q(\u2/L9 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [20]),
        .Q(\u2/L9 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [21]),
        .Q(\u2/L9 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [22]),
        .Q(\u2/L9 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [23]),
        .Q(\u2/L9 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [24]),
        .Q(\u2/L9 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [25]),
        .Q(\u2/L9 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [26]),
        .Q(\u2/L9 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [27]),
        .Q(\u2/L9 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [28]),
        .Q(\u2/L9 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [29]),
        .Q(\u2/L9 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [2]),
        .Q(\u2/L9 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [30]),
        .Q(\u2/L9 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [31]),
        .Q(\u2/L9 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [32]),
        .Q(\u2/L9 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [3]),
        .Q(\u2/L9 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [4]),
        .Q(\u2/L9 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [5]),
        .Q(\u2/L9 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [6]),
        .Q(\u2/L9 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [7]),
        .Q(\u2/L9 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [8]),
        .Q(\u2/L9 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/L9_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R8 [9]),
        .Q(\u2/L9 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[10]_i_1 
       (.I0(\u2/IP [10]),
        .I1(\u2/out0 [10]),
        .O(\u2/R00 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[11]_i_1 
       (.I0(\u2/IP [11]),
        .I1(\u2/out0 [11]),
        .O(\u2/R00 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[12]_i_1 
       (.I0(\u2/IP [12]),
        .I1(\u2/out0 [12]),
        .O(\u2/R00 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[13]_i_1 
       (.I0(\u2/IP [13]),
        .I1(\u2/out0 [13]),
        .O(\u2/R00 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[14]_i_1 
       (.I0(\u2/IP [14]),
        .I1(\u2/out0 [14]),
        .O(\u2/R00 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[15]_i_1 
       (.I0(\u2/IP [15]),
        .I1(\u2/out0 [15]),
        .O(\u2/R00 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[16]_i_1 
       (.I0(\u2/IP [16]),
        .I1(\u2/out0 [16]),
        .O(\u2/R00 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[17]_i_1 
       (.I0(\u2/IP [17]),
        .I1(\u2/out0 [17]),
        .O(\u2/R00 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[18]_i_1 
       (.I0(\u2/IP [18]),
        .I1(\u2/out0 [18]),
        .O(\u2/R00 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[19]_i_1 
       (.I0(\u2/IP [19]),
        .I1(\u2/out0 [19]),
        .O(\u2/R00 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[1]_i_1 
       (.I0(\u2/IP [1]),
        .I1(\u2/out0 [1]),
        .O(\u2/R00 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[20]_i_1 
       (.I0(\u2/IP [20]),
        .I1(\u2/out0 [20]),
        .O(\u2/R00 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[21]_i_1 
       (.I0(\u2/IP [21]),
        .I1(\u2/out0 [21]),
        .O(\u2/R00 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[22]_i_1 
       (.I0(\u2/IP [22]),
        .I1(\u2/out0 [22]),
        .O(\u2/R00 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[23]_i_1 
       (.I0(\u2/IP [23]),
        .I1(\u2/out0 [23]),
        .O(\u2/R00 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[24]_i_1 
       (.I0(\u2/IP [24]),
        .I1(\u2/out0 [24]),
        .O(\u2/R00 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[25]_i_1 
       (.I0(\u2/IP [25]),
        .I1(\u2/out0 [25]),
        .O(\u2/R00 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[26]_i_1 
       (.I0(\u2/IP [26]),
        .I1(\u2/out0 [26]),
        .O(\u2/R00 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[27]_i_1 
       (.I0(\u2/IP [27]),
        .I1(\u2/out0 [27]),
        .O(\u2/R00 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[28]_i_1 
       (.I0(\u2/IP [28]),
        .I1(\u2/out0 [28]),
        .O(\u2/R00 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[29]_i_1 
       (.I0(\u2/IP [29]),
        .I1(\u2/out0 [29]),
        .O(\u2/R00 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[2]_i_1 
       (.I0(\u2/IP [2]),
        .I1(\u2/out0 [2]),
        .O(\u2/R00 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[30]_i_1 
       (.I0(\u2/IP [30]),
        .I1(\u2/out0 [30]),
        .O(\u2/R00 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[31]_i_1 
       (.I0(\u2/IP [31]),
        .I1(\u2/out0 [31]),
        .O(\u2/R00 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[32]_i_1 
       (.I0(\u2/IP [32]),
        .I1(\u2/out0 [32]),
        .O(\u2/R00 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[3]_i_1 
       (.I0(\u2/IP [3]),
        .I1(\u2/out0 [3]),
        .O(\u2/R00 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[4]_i_1 
       (.I0(\u2/IP [4]),
        .I1(\u2/out0 [4]),
        .O(\u2/R00 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[5]_i_1 
       (.I0(\u2/IP [5]),
        .I1(\u2/out0 [5]),
        .O(\u2/R00 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[6]_i_1 
       (.I0(\u2/IP [6]),
        .I1(\u2/out0 [6]),
        .O(\u2/R00 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[7]_i_1 
       (.I0(\u2/IP [7]),
        .I1(\u2/out0 [7]),
        .O(\u2/R00 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[8]_i_1 
       (.I0(\u2/IP [8]),
        .I1(\u2/out0 [8]),
        .O(\u2/R00 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R0[9]_i_1 
       (.I0(\u2/IP [9]),
        .I1(\u2/out0 [9]),
        .O(\u2/R00 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [22]),
        .Q(\u2/R0 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [21]),
        .Q(\u2/R0 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [20]),
        .Q(\u2/R0 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [19]),
        .Q(\u2/R0 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [18]),
        .Q(\u2/R0 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [17]),
        .Q(\u2/R0 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [16]),
        .Q(\u2/R0 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [15]),
        .Q(\u2/R0 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [14]),
        .Q(\u2/R0 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [13]),
        .Q(\u2/R0 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [31]),
        .Q(\u2/R0 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [12]),
        .Q(\u2/R0 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [11]),
        .Q(\u2/R0 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [10]),
        .Q(\u2/R0 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [9]),
        .Q(\u2/R0 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [8]),
        .Q(\u2/R0 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [7]),
        .Q(\u2/R0 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [6]),
        .Q(\u2/R0 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [5]),
        .Q(\u2/R0 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [4]),
        .Q(\u2/R0 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [3]),
        .Q(\u2/R0 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [30]),
        .Q(\u2/R0 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [2]),
        .Q(\u2/R0 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [1]),
        .Q(\u2/R0 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [0]),
        .Q(\u2/R0 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [29]),
        .Q(\u2/R0 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [28]),
        .Q(\u2/R0 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [27]),
        .Q(\u2/R0 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [26]),
        .Q(\u2/R0 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [25]),
        .Q(\u2/R0 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [24]),
        .Q(\u2/R0 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R0_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R00 [23]),
        .Q(\u2/R0 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[10]_i_1 
       (.I0(\u2/L9 [10]),
        .I1(\u2/out10 [10]),
        .O(\u2/R100 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[11]_i_1 
       (.I0(\u2/L9 [11]),
        .I1(\u2/out10 [11]),
        .O(\u2/R100 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[12]_i_1 
       (.I0(\u2/L9 [12]),
        .I1(\u2/out10 [12]),
        .O(\u2/R100 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[13]_i_1 
       (.I0(\u2/L9 [13]),
        .I1(\u2/out10 [13]),
        .O(\u2/R100 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[14]_i_1 
       (.I0(\u2/L9 [14]),
        .I1(\u2/out10 [14]),
        .O(\u2/R100 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[15]_i_1 
       (.I0(\u2/L9 [15]),
        .I1(\u2/out10 [15]),
        .O(\u2/R100 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[16]_i_1 
       (.I0(\u2/L9 [16]),
        .I1(\u2/out10 [16]),
        .O(\u2/R100 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[17]_i_1 
       (.I0(\u2/L9 [17]),
        .I1(\u2/out10 [17]),
        .O(\u2/R100 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[18]_i_1 
       (.I0(\u2/L9 [18]),
        .I1(\u2/out10 [18]),
        .O(\u2/R100 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[19]_i_1 
       (.I0(\u2/L9 [19]),
        .I1(\u2/out10 [19]),
        .O(\u2/R100 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[1]_i_1 
       (.I0(\u2/L9 [1]),
        .I1(\u2/out10 [1]),
        .O(\u2/R100 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[20]_i_1 
       (.I0(\u2/L9 [20]),
        .I1(\u2/out10 [20]),
        .O(\u2/R100 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[21]_i_1 
       (.I0(\u2/L9 [21]),
        .I1(\u2/out10 [21]),
        .O(\u2/R100 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[22]_i_1 
       (.I0(\u2/L9 [22]),
        .I1(\u2/out10 [22]),
        .O(\u2/R100 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[23]_i_1 
       (.I0(\u2/L9 [23]),
        .I1(\u2/out10 [23]),
        .O(\u2/R100 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[24]_i_1 
       (.I0(\u2/L9 [24]),
        .I1(\u2/out10 [24]),
        .O(\u2/R100 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[25]_i_1 
       (.I0(\u2/L9 [25]),
        .I1(\u2/out10 [25]),
        .O(\u2/R100 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[26]_i_1 
       (.I0(\u2/L9 [26]),
        .I1(\u2/out10 [26]),
        .O(\u2/R100 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[27]_i_1 
       (.I0(\u2/L9 [27]),
        .I1(\u2/out10 [27]),
        .O(\u2/R100 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[28]_i_1 
       (.I0(\u2/L9 [28]),
        .I1(\u2/out10 [28]),
        .O(\u2/R100 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[29]_i_1 
       (.I0(\u2/L9 [29]),
        .I1(\u2/out10 [29]),
        .O(\u2/R100 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[2]_i_1 
       (.I0(\u2/L9 [2]),
        .I1(\u2/out10 [2]),
        .O(\u2/R100 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[30]_i_1 
       (.I0(\u2/L9 [30]),
        .I1(\u2/out10 [30]),
        .O(\u2/R100 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[31]_i_1 
       (.I0(\u2/L9 [31]),
        .I1(\u2/out10 [31]),
        .O(\u2/R100 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[32]_i_1 
       (.I0(\u2/L9 [32]),
        .I1(\u2/out10 [32]),
        .O(\u2/R100 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[3]_i_1 
       (.I0(\u2/L9 [3]),
        .I1(\u2/out10 [3]),
        .O(\u2/R100 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[4]_i_1 
       (.I0(\u2/L9 [4]),
        .I1(\u2/out10 [4]),
        .O(\u2/R100 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[5]_i_1 
       (.I0(\u2/L9 [5]),
        .I1(\u2/out10 [5]),
        .O(\u2/R100 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[6]_i_1 
       (.I0(\u2/L9 [6]),
        .I1(\u2/out10 [6]),
        .O(\u2/R100 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[7]_i_1 
       (.I0(\u2/L9 [7]),
        .I1(\u2/out10 [7]),
        .O(\u2/R100 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[8]_i_1 
       (.I0(\u2/L9 [8]),
        .I1(\u2/out10 [8]),
        .O(\u2/R100 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R10[9]_i_1 
       (.I0(\u2/L9 [9]),
        .I1(\u2/out10 [9]),
        .O(\u2/R100 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [22]),
        .Q(\u2/R10_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [21]),
        .Q(\u2/R10_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [20]),
        .Q(\u2/R10_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [19]),
        .Q(\u2/R10_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [18]),
        .Q(\u2/R10_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [17]),
        .Q(\u2/R10_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [16]),
        .Q(\u2/R10_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [15]),
        .Q(\u2/R10_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [14]),
        .Q(\u2/R10_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [13]),
        .Q(\u2/R10_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [31]),
        .Q(\u2/R10_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [12]),
        .Q(\u2/R10_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [11]),
        .Q(\u2/R10_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [10]),
        .Q(\u2/R10_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [9]),
        .Q(\u2/R10_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [8]),
        .Q(\u2/R10_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [7]),
        .Q(\u2/R10_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [6]),
        .Q(\u2/R10_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [5]),
        .Q(\u2/R10_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [4]),
        .Q(\u2/R10_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [3]),
        .Q(\u2/R10_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [30]),
        .Q(\u2/R10_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [2]),
        .Q(\u2/R10_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [1]),
        .Q(\u2/R10_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [0]),
        .Q(\u2/R10_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [29]),
        .Q(\u2/R10_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [28]),
        .Q(\u2/R10_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [27]),
        .Q(\u2/R10_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [26]),
        .Q(\u2/R10_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [25]),
        .Q(\u2/R10_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [24]),
        .Q(\u2/R10_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R10_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R100 [23]),
        .Q(\u2/R10_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[10]_i_1 
       (.I0(\u2/L10 [10]),
        .I1(\u2/out11 [10]),
        .O(\u2/R110 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[11]_i_1 
       (.I0(\u2/L10 [11]),
        .I1(\u2/out11 [11]),
        .O(\u2/R110 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[12]_i_1 
       (.I0(\u2/L10 [12]),
        .I1(\u2/out11 [12]),
        .O(\u2/R110 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[13]_i_1 
       (.I0(\u2/L10 [13]),
        .I1(\u2/out11 [13]),
        .O(\u2/R110 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[14]_i_1 
       (.I0(\u2/L10 [14]),
        .I1(\u2/out11 [14]),
        .O(\u2/R110 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[15]_i_1 
       (.I0(\u2/L10 [15]),
        .I1(\u2/out11 [15]),
        .O(\u2/R110 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[16]_i_1 
       (.I0(\u2/L10 [16]),
        .I1(\u2/out11 [16]),
        .O(\u2/R110 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[17]_i_1 
       (.I0(\u2/L10 [17]),
        .I1(\u2/out11 [17]),
        .O(\u2/R110 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[18]_i_1 
       (.I0(\u2/L10 [18]),
        .I1(\u2/out11 [18]),
        .O(\u2/R110 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[19]_i_1 
       (.I0(\u2/L10 [19]),
        .I1(\u2/out11 [19]),
        .O(\u2/R110 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[1]_i_1 
       (.I0(\u2/L10 [1]),
        .I1(\u2/out11 [1]),
        .O(\u2/R110 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[20]_i_1 
       (.I0(\u2/L10 [20]),
        .I1(\u2/out11 [20]),
        .O(\u2/R110 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[21]_i_1 
       (.I0(\u2/L10 [21]),
        .I1(\u2/out11 [21]),
        .O(\u2/R110 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[22]_i_1 
       (.I0(\u2/L10 [22]),
        .I1(\u2/out11 [22]),
        .O(\u2/R110 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[23]_i_1 
       (.I0(\u2/L10 [23]),
        .I1(\u2/out11 [23]),
        .O(\u2/R110 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[24]_i_1 
       (.I0(\u2/L10 [24]),
        .I1(\u2/out11 [24]),
        .O(\u2/R110 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[25]_i_1 
       (.I0(\u2/L10 [25]),
        .I1(\u2/out11 [25]),
        .O(\u2/R110 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[26]_i_1 
       (.I0(\u2/L10 [26]),
        .I1(\u2/out11 [26]),
        .O(\u2/R110 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[27]_i_1 
       (.I0(\u2/L10 [27]),
        .I1(\u2/out11 [27]),
        .O(\u2/R110 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[28]_i_1 
       (.I0(\u2/L10 [28]),
        .I1(\u2/out11 [28]),
        .O(\u2/R110 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[29]_i_1 
       (.I0(\u2/L10 [29]),
        .I1(\u2/out11 [29]),
        .O(\u2/R110 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[2]_i_1 
       (.I0(\u2/L10 [2]),
        .I1(\u2/out11 [2]),
        .O(\u2/R110 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[30]_i_1 
       (.I0(\u2/L10 [30]),
        .I1(\u2/out11 [30]),
        .O(\u2/R110 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[31]_i_1 
       (.I0(\u2/L10 [31]),
        .I1(\u2/out11 [31]),
        .O(\u2/R110 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[32]_i_1 
       (.I0(\u2/L10 [32]),
        .I1(\u2/out11 [32]),
        .O(\u2/R110 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[3]_i_1 
       (.I0(\u2/L10 [3]),
        .I1(\u2/out11 [3]),
        .O(\u2/R110 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[4]_i_1 
       (.I0(\u2/L10 [4]),
        .I1(\u2/out11 [4]),
        .O(\u2/R110 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[5]_i_1 
       (.I0(\u2/L10 [5]),
        .I1(\u2/out11 [5]),
        .O(\u2/R110 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[6]_i_1 
       (.I0(\u2/L10 [6]),
        .I1(\u2/out11 [6]),
        .O(\u2/R110 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[7]_i_1 
       (.I0(\u2/L10 [7]),
        .I1(\u2/out11 [7]),
        .O(\u2/R110 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[8]_i_1 
       (.I0(\u2/L10 [8]),
        .I1(\u2/out11 [8]),
        .O(\u2/R110 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R11[9]_i_1 
       (.I0(\u2/L10 [9]),
        .I1(\u2/out11 [9]),
        .O(\u2/R110 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [22]),
        .Q(\u2/R11 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [21]),
        .Q(\u2/R11 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [20]),
        .Q(\u2/R11 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [19]),
        .Q(\u2/R11 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [18]),
        .Q(\u2/R11 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [17]),
        .Q(\u2/R11 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [16]),
        .Q(\u2/R11 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [15]),
        .Q(\u2/R11 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [14]),
        .Q(\u2/R11 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [13]),
        .Q(\u2/R11 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [31]),
        .Q(\u2/R11 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [12]),
        .Q(\u2/R11 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [11]),
        .Q(\u2/R11 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [10]),
        .Q(\u2/R11 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [9]),
        .Q(\u2/R11 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [8]),
        .Q(\u2/R11 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [7]),
        .Q(\u2/R11 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [6]),
        .Q(\u2/R11 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [5]),
        .Q(\u2/R11 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [4]),
        .Q(\u2/R11 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [3]),
        .Q(\u2/R11 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [30]),
        .Q(\u2/R11 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [2]),
        .Q(\u2/R11 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [1]),
        .Q(\u2/R11 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [0]),
        .Q(\u2/R11 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [29]),
        .Q(\u2/R11 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [28]),
        .Q(\u2/R11 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [27]),
        .Q(\u2/R11 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [26]),
        .Q(\u2/R11 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [25]),
        .Q(\u2/R11 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [24]),
        .Q(\u2/R11 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R11_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R110 [23]),
        .Q(\u2/R11 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[10]_i_1 
       (.I0(\u2/L11 [10]),
        .I1(\u2/out12 [10]),
        .O(\u2/R120 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[11]_i_1 
       (.I0(\u2/L11 [11]),
        .I1(\u2/out12 [11]),
        .O(\u2/R120 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[12]_i_1 
       (.I0(\u2/L11 [12]),
        .I1(\u2/out12 [12]),
        .O(\u2/R120 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[13]_i_1 
       (.I0(\u2/L11 [13]),
        .I1(\u2/out12 [13]),
        .O(\u2/R120 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[14]_i_1 
       (.I0(\u2/L11 [14]),
        .I1(\u2/out12 [14]),
        .O(\u2/R120 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[15]_i_1 
       (.I0(\u2/L11 [15]),
        .I1(\u2/out12 [15]),
        .O(\u2/R120 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[16]_i_1 
       (.I0(\u2/L11 [16]),
        .I1(\u2/out12 [16]),
        .O(\u2/R120 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[17]_i_1 
       (.I0(\u2/L11 [17]),
        .I1(\u2/out12 [17]),
        .O(\u2/R120 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[18]_i_1 
       (.I0(\u2/L11 [18]),
        .I1(\u2/out12 [18]),
        .O(\u2/R120 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[19]_i_1 
       (.I0(\u2/L11 [19]),
        .I1(\u2/out12 [19]),
        .O(\u2/R120 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[1]_i_1 
       (.I0(\u2/L11 [1]),
        .I1(\u2/out12 [1]),
        .O(\u2/R120 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[20]_i_1 
       (.I0(\u2/L11 [20]),
        .I1(\u2/out12 [20]),
        .O(\u2/R120 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[21]_i_1 
       (.I0(\u2/L11 [21]),
        .I1(\u2/out12 [21]),
        .O(\u2/R120 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[22]_i_1 
       (.I0(\u2/L11 [22]),
        .I1(\u2/out12 [22]),
        .O(\u2/R120 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[23]_i_1 
       (.I0(\u2/L11 [23]),
        .I1(\u2/out12 [23]),
        .O(\u2/R120 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[24]_i_1 
       (.I0(\u2/L11 [24]),
        .I1(\u2/out12 [24]),
        .O(\u2/R120 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[25]_i_1 
       (.I0(\u2/L11 [25]),
        .I1(\u2/out12 [25]),
        .O(\u2/R120 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[26]_i_1 
       (.I0(\u2/L11 [26]),
        .I1(\u2/out12 [26]),
        .O(\u2/R120 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[27]_i_1 
       (.I0(\u2/L11 [27]),
        .I1(\u2/out12 [27]),
        .O(\u2/R120 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[28]_i_1 
       (.I0(\u2/L11 [28]),
        .I1(\u2/out12 [28]),
        .O(\u2/R120 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[29]_i_1 
       (.I0(\u2/L11 [29]),
        .I1(\u2/out12 [29]),
        .O(\u2/R120 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[2]_i_1 
       (.I0(\u2/L11 [2]),
        .I1(\u2/out12 [2]),
        .O(\u2/R120 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[30]_i_1 
       (.I0(\u2/L11 [30]),
        .I1(\u2/out12 [30]),
        .O(\u2/R120 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[31]_i_1 
       (.I0(\u2/L11 [31]),
        .I1(\u2/out12 [31]),
        .O(\u2/R120 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[32]_i_1 
       (.I0(\u2/L11 [32]),
        .I1(\u2/out12 [32]),
        .O(\u2/R120 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[3]_i_1 
       (.I0(\u2/L11 [3]),
        .I1(\u2/out12 [3]),
        .O(\u2/R120 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[4]_i_1 
       (.I0(\u2/L11 [4]),
        .I1(\u2/out12 [4]),
        .O(\u2/R120 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[5]_i_1 
       (.I0(\u2/L11 [5]),
        .I1(\u2/out12 [5]),
        .O(\u2/R120 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[6]_i_1 
       (.I0(\u2/L11 [6]),
        .I1(\u2/out12 [6]),
        .O(\u2/R120 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[7]_i_1 
       (.I0(\u2/L11 [7]),
        .I1(\u2/out12 [7]),
        .O(\u2/R120 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[8]_i_1 
       (.I0(\u2/L11 [8]),
        .I1(\u2/out12 [8]),
        .O(\u2/R120 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R12[9]_i_1 
       (.I0(\u2/L11 [9]),
        .I1(\u2/out12 [9]),
        .O(\u2/R120 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [22]),
        .Q(\u2/R12 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [21]),
        .Q(\u2/R12 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [20]),
        .Q(\u2/R12 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [19]),
        .Q(\u2/R12 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [18]),
        .Q(\u2/R12 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [17]),
        .Q(\u2/R12 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [16]),
        .Q(\u2/R12 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [15]),
        .Q(\u2/R12 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [14]),
        .Q(\u2/R12 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [13]),
        .Q(\u2/R12 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [31]),
        .Q(\u2/R12 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [12]),
        .Q(\u2/R12 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [11]),
        .Q(\u2/R12 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [10]),
        .Q(\u2/R12 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [9]),
        .Q(\u2/R12 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [8]),
        .Q(\u2/R12 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [7]),
        .Q(\u2/R12 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [6]),
        .Q(\u2/R12 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [5]),
        .Q(\u2/R12 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [4]),
        .Q(\u2/R12 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [3]),
        .Q(\u2/R12 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [30]),
        .Q(\u2/R12 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [2]),
        .Q(\u2/R12 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [1]),
        .Q(\u2/R12 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [0]),
        .Q(\u2/R12 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [29]),
        .Q(\u2/R12 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [28]),
        .Q(\u2/R12 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [27]),
        .Q(\u2/R12 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [26]),
        .Q(\u2/R12 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [25]),
        .Q(\u2/R12 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [24]),
        .Q(\u2/R12 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R12_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R120 [23]),
        .Q(\u2/R12 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[10]_i_1 
       (.I0(\u2/L12 [10]),
        .I1(\u2/out13 [10]),
        .O(\u2/R130 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[11]_i_1 
       (.I0(\u2/L12 [11]),
        .I1(\u2/out13 [11]),
        .O(\u2/R130 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[12]_i_1 
       (.I0(\u2/L12 [12]),
        .I1(\u2/out13 [12]),
        .O(\u2/R130 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[13]_i_1 
       (.I0(\u2/L12 [13]),
        .I1(\u2/out13 [13]),
        .O(\u2/R130 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[14]_i_1 
       (.I0(\u2/L12 [14]),
        .I1(\u2/out13 [14]),
        .O(\u2/R130 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[15]_i_1 
       (.I0(\u2/L12 [15]),
        .I1(\u2/out13 [15]),
        .O(\u2/R130 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[16]_i_1 
       (.I0(\u2/L12 [16]),
        .I1(\u2/out13 [16]),
        .O(\u2/R130 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[17]_i_1 
       (.I0(\u2/L12 [17]),
        .I1(\u2/out13 [17]),
        .O(\u2/R130 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[18]_i_1 
       (.I0(\u2/L12 [18]),
        .I1(\u2/out13 [18]),
        .O(\u2/R130 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[19]_i_1 
       (.I0(\u2/L12 [19]),
        .I1(\u2/out13 [19]),
        .O(\u2/R130 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[1]_i_1 
       (.I0(\u2/L12 [1]),
        .I1(\u2/out13 [1]),
        .O(\u2/R130 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[20]_i_1 
       (.I0(\u2/L12 [20]),
        .I1(\u2/out13 [20]),
        .O(\u2/R130 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[21]_i_1 
       (.I0(\u2/L12 [21]),
        .I1(\u2/out13 [21]),
        .O(\u2/R130 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[22]_i_1 
       (.I0(\u2/L12 [22]),
        .I1(\u2/out13 [22]),
        .O(\u2/R130 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[23]_i_1 
       (.I0(\u2/L12 [23]),
        .I1(\u2/out13 [23]),
        .O(\u2/R130 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[24]_i_1 
       (.I0(\u2/L12 [24]),
        .I1(\u2/out13 [24]),
        .O(\u2/R130 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[25]_i_1 
       (.I0(\u2/L12 [25]),
        .I1(\u2/out13 [25]),
        .O(\u2/R130 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[26]_i_1 
       (.I0(\u2/L12 [26]),
        .I1(\u2/out13 [26]),
        .O(\u2/R130 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[27]_i_1 
       (.I0(\u2/L12 [27]),
        .I1(\u2/out13 [27]),
        .O(\u2/R130 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[28]_i_1 
       (.I0(\u2/L12 [28]),
        .I1(\u2/out13 [28]),
        .O(\u2/R130 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[29]_i_1 
       (.I0(\u2/L12 [29]),
        .I1(\u2/out13 [29]),
        .O(\u2/R130 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[2]_i_1 
       (.I0(\u2/L12 [2]),
        .I1(\u2/out13 [2]),
        .O(\u2/R130 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[30]_i_1 
       (.I0(\u2/L12 [30]),
        .I1(\u2/out13 [30]),
        .O(\u2/R130 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[31]_i_1 
       (.I0(\u2/L12 [31]),
        .I1(\u2/out13 [31]),
        .O(\u2/R130 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[32]_i_1 
       (.I0(\u2/L12 [32]),
        .I1(\u2/out13 [32]),
        .O(\u2/R130 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[3]_i_1 
       (.I0(\u2/L12 [3]),
        .I1(\u2/out13 [3]),
        .O(\u2/R130 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[4]_i_1 
       (.I0(\u2/L12 [4]),
        .I1(\u2/out13 [4]),
        .O(\u2/R130 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[5]_i_1 
       (.I0(\u2/L12 [5]),
        .I1(\u2/out13 [5]),
        .O(\u2/R130 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[6]_i_1 
       (.I0(\u2/L12 [6]),
        .I1(\u2/out13 [6]),
        .O(\u2/R130 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[7]_i_1 
       (.I0(\u2/L12 [7]),
        .I1(\u2/out13 [7]),
        .O(\u2/R130 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[8]_i_1 
       (.I0(\u2/L12 [8]),
        .I1(\u2/out13 [8]),
        .O(\u2/R130 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R13[9]_i_1 
       (.I0(\u2/L12 [9]),
        .I1(\u2/out13 [9]),
        .O(\u2/R130 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [22]),
        .Q(\u2/R13 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [21]),
        .Q(\u2/R13 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [20]),
        .Q(\u2/R13 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [19]),
        .Q(\u2/R13 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [18]),
        .Q(\u2/R13 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [17]),
        .Q(\u2/R13 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [16]),
        .Q(\u2/R13 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [15]),
        .Q(\u2/R13 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [14]),
        .Q(\u2/R13 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [13]),
        .Q(\u2/R13 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [31]),
        .Q(\u2/R13 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [12]),
        .Q(\u2/R13 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [11]),
        .Q(\u2/R13 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [10]),
        .Q(\u2/R13 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [9]),
        .Q(\u2/R13 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [8]),
        .Q(\u2/R13 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [7]),
        .Q(\u2/R13 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [6]),
        .Q(\u2/R13 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [5]),
        .Q(\u2/R13 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [4]),
        .Q(\u2/R13 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [3]),
        .Q(\u2/R13 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [30]),
        .Q(\u2/R13 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [2]),
        .Q(\u2/R13 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [1]),
        .Q(\u2/R13 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [0]),
        .Q(\u2/R13 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [29]),
        .Q(\u2/R13 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [28]),
        .Q(\u2/R13 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [27]),
        .Q(\u2/R13 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [26]),
        .Q(\u2/R13 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [25]),
        .Q(\u2/R13 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [24]),
        .Q(\u2/R13 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R13_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R130 [23]),
        .Q(\u2/R13 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[10]_i_1 
       (.I0(\u2/L13 [10]),
        .I1(\u2/out14 [10]),
        .O(\u2/R140 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[11]_i_1 
       (.I0(\u2/L13 [11]),
        .I1(\u2/out14 [11]),
        .O(\u2/R140 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[12]_i_1 
       (.I0(\u2/L13 [12]),
        .I1(\u2/out14 [12]),
        .O(\u2/R140 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[13]_i_1 
       (.I0(\u2/L13 [13]),
        .I1(\u2/out14 [13]),
        .O(\u2/R140 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[14]_i_1 
       (.I0(\u2/L13 [14]),
        .I1(\u2/out14 [14]),
        .O(\u2/R140 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[15]_i_1 
       (.I0(\u2/L13 [15]),
        .I1(\u2/out14 [15]),
        .O(\u2/R140 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[16]_i_1 
       (.I0(\u2/L13 [16]),
        .I1(\u2/out14 [16]),
        .O(\u2/R140 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[17]_i_1 
       (.I0(\u2/L13 [17]),
        .I1(\u2/out14 [17]),
        .O(\u2/R140 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[18]_i_1 
       (.I0(\u2/L13 [18]),
        .I1(\u2/out14 [18]),
        .O(\u2/R140 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[19]_i_1 
       (.I0(\u2/L13 [19]),
        .I1(\u2/out14 [19]),
        .O(\u2/R140 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[1]_i_1 
       (.I0(\u2/L13 [1]),
        .I1(\u2/out14 [1]),
        .O(\u2/R140 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[20]_i_1 
       (.I0(\u2/L13 [20]),
        .I1(\u2/out14 [20]),
        .O(\u2/R140 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[21]_i_1 
       (.I0(\u2/L13 [21]),
        .I1(\u2/out14 [21]),
        .O(\u2/R140 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[22]_i_1 
       (.I0(\u2/L13 [22]),
        .I1(\u2/out14 [22]),
        .O(\u2/R140 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[23]_i_1 
       (.I0(\u2/L13 [23]),
        .I1(\u2/out14 [23]),
        .O(\u2/R140 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[24]_i_1 
       (.I0(\u2/L13 [24]),
        .I1(\u2/out14 [24]),
        .O(\u2/R140 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[25]_i_1 
       (.I0(\u2/L13 [25]),
        .I1(\u2/out14 [25]),
        .O(\u2/R140 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[26]_i_1 
       (.I0(\u2/L13 [26]),
        .I1(\u2/out14 [26]),
        .O(\u2/R140 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[27]_i_1 
       (.I0(\u2/L13 [27]),
        .I1(\u2/out14 [27]),
        .O(\u2/R140 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[28]_i_1 
       (.I0(\u2/L13 [28]),
        .I1(\u2/out14 [28]),
        .O(\u2/R140 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[29]_i_1 
       (.I0(\u2/L13 [29]),
        .I1(\u2/out14 [29]),
        .O(\u2/R140 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[2]_i_1 
       (.I0(\u2/L13 [2]),
        .I1(\u2/out14 [2]),
        .O(\u2/R140 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[30]_i_1 
       (.I0(\u2/L13 [30]),
        .I1(\u2/out14 [30]),
        .O(\u2/R140 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[31]_i_1 
       (.I0(\u2/L13 [31]),
        .I1(\u2/out14 [31]),
        .O(\u2/R140 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[32]_i_1 
       (.I0(\u2/L13 [32]),
        .I1(\u2/out14 [32]),
        .O(\u2/R140 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[3]_i_1 
       (.I0(\u2/L13 [3]),
        .I1(\u2/out14 [3]),
        .O(\u2/R140 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[4]_i_1 
       (.I0(\u2/L13 [4]),
        .I1(\u2/out14 [4]),
        .O(\u2/R140 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[5]_i_1 
       (.I0(\u2/L13 [5]),
        .I1(\u2/out14 [5]),
        .O(\u2/R140 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[6]_i_1 
       (.I0(\u2/L13 [6]),
        .I1(\u2/out14 [6]),
        .O(\u2/R140 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[7]_i_1 
       (.I0(\u2/L13 [7]),
        .I1(\u2/out14 [7]),
        .O(\u2/R140 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[8]_i_1 
       (.I0(\u2/L13 [8]),
        .I1(\u2/out14 [8]),
        .O(\u2/R140 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R14[9]_i_1 
       (.I0(\u2/L13 [9]),
        .I1(\u2/out14 [9]),
        .O(\u2/R140 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [22]),
        .Q(\u2/FP [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [21]),
        .Q(\u2/FP [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [20]),
        .Q(\u2/FP [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [19]),
        .Q(\u2/FP [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [18]),
        .Q(\u2/FP [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [17]),
        .Q(\u2/FP [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [16]),
        .Q(\u2/FP [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [15]),
        .Q(\u2/FP [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [14]),
        .Q(\u2/FP [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [13]),
        .Q(\u2/FP [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [31]),
        .Q(\u2/FP [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [12]),
        .Q(\u2/FP [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [11]),
        .Q(\u2/FP [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [10]),
        .Q(\u2/FP [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [9]),
        .Q(\u2/FP [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [8]),
        .Q(\u2/FP [56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [7]),
        .Q(\u2/FP [57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [6]),
        .Q(\u2/FP [58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [5]),
        .Q(\u2/FP [59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [4]),
        .Q(\u2/FP [60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [3]),
        .Q(\u2/FP [61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [30]),
        .Q(\u2/FP [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [2]),
        .Q(\u2/FP [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [1]),
        .Q(\u2/FP [63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [0]),
        .Q(\u2/FP [64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [29]),
        .Q(\u2/FP [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [28]),
        .Q(\u2/FP [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [27]),
        .Q(\u2/FP [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [26]),
        .Q(\u2/FP [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [25]),
        .Q(\u2/FP [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [24]),
        .Q(\u2/FP [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R14_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R140 [23]),
        .Q(\u2/FP [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[10]_i_1 
       (.I0(\u2/L0 [10]),
        .I1(\u2/out1 [10]),
        .O(\u2/R10 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[11]_i_1 
       (.I0(\u2/L0 [11]),
        .I1(\u2/out1 [11]),
        .O(\u2/R10 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[12]_i_1 
       (.I0(\u2/L0 [12]),
        .I1(\u2/out1 [12]),
        .O(\u2/R10 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[13]_i_1 
       (.I0(\u2/L0 [13]),
        .I1(\u2/out1 [13]),
        .O(\u2/R10 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[14]_i_1 
       (.I0(\u2/L0 [14]),
        .I1(\u2/out1 [14]),
        .O(\u2/R10 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[15]_i_1 
       (.I0(\u2/L0 [15]),
        .I1(\u2/out1 [15]),
        .O(\u2/R10 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[16]_i_1 
       (.I0(\u2/L0 [16]),
        .I1(\u2/out1 [16]),
        .O(\u2/R10 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[17]_i_1 
       (.I0(\u2/L0 [17]),
        .I1(\u2/out1 [17]),
        .O(\u2/R10 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[18]_i_1 
       (.I0(\u2/L0 [18]),
        .I1(\u2/out1 [18]),
        .O(\u2/R10 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[19]_i_1 
       (.I0(\u2/L0 [19]),
        .I1(\u2/out1 [19]),
        .O(\u2/R10 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[1]_i_1 
       (.I0(\u2/L0 [1]),
        .I1(\u2/out1 [1]),
        .O(\u2/R10 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[20]_i_1 
       (.I0(\u2/L0 [20]),
        .I1(\u2/out1 [20]),
        .O(\u2/R10 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[21]_i_1 
       (.I0(\u2/L0 [21]),
        .I1(\u2/out1 [21]),
        .O(\u2/R10 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[22]_i_1 
       (.I0(\u2/L0 [22]),
        .I1(\u2/out1 [22]),
        .O(\u2/R10 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[23]_i_1 
       (.I0(\u2/L0 [23]),
        .I1(\u2/out1 [23]),
        .O(\u2/R10 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[24]_i_1 
       (.I0(\u2/L0 [24]),
        .I1(\u2/out1 [24]),
        .O(\u2/R10 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[25]_i_1 
       (.I0(\u2/L0 [25]),
        .I1(\u2/out1 [25]),
        .O(\u2/R10 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[26]_i_1 
       (.I0(\u2/L0 [26]),
        .I1(\u2/out1 [26]),
        .O(\u2/R10 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[27]_i_1 
       (.I0(\u2/L0 [27]),
        .I1(\u2/out1 [27]),
        .O(\u2/R10 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[28]_i_1 
       (.I0(\u2/L0 [28]),
        .I1(\u2/out1 [28]),
        .O(\u2/R10 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[29]_i_1 
       (.I0(\u2/L0 [29]),
        .I1(\u2/out1 [29]),
        .O(\u2/R10 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[2]_i_1 
       (.I0(\u2/L0 [2]),
        .I1(\u2/out1 [2]),
        .O(\u2/R10 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[30]_i_1 
       (.I0(\u2/L0 [30]),
        .I1(\u2/out1 [30]),
        .O(\u2/R10 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[31]_i_1 
       (.I0(\u2/L0 [31]),
        .I1(\u2/out1 [31]),
        .O(\u2/R10 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[32]_i_1 
       (.I0(\u2/L0 [32]),
        .I1(\u2/out1 [32]),
        .O(\u2/R10 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[3]_i_1 
       (.I0(\u2/L0 [3]),
        .I1(\u2/out1 [3]),
        .O(\u2/R10 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[4]_i_1 
       (.I0(\u2/L0 [4]),
        .I1(\u2/out1 [4]),
        .O(\u2/R10 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[5]_i_1 
       (.I0(\u2/L0 [5]),
        .I1(\u2/out1 [5]),
        .O(\u2/R10 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[6]_i_1 
       (.I0(\u2/L0 [6]),
        .I1(\u2/out1 [6]),
        .O(\u2/R10 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[7]_i_1 
       (.I0(\u2/L0 [7]),
        .I1(\u2/out1 [7]),
        .O(\u2/R10 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[8]_i_1 
       (.I0(\u2/L0 [8]),
        .I1(\u2/out1 [8]),
        .O(\u2/R10 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R1[9]_i_1 
       (.I0(\u2/L0 [9]),
        .I1(\u2/out1 [9]),
        .O(\u2/R10 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [22]),
        .Q(\u2/R1 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [21]),
        .Q(\u2/R1 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [20]),
        .Q(\u2/R1 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [19]),
        .Q(\u2/R1 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [18]),
        .Q(\u2/R1 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [17]),
        .Q(\u2/R1 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [16]),
        .Q(\u2/R1 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [15]),
        .Q(\u2/R1 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [14]),
        .Q(\u2/R1 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [13]),
        .Q(\u2/R1 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [31]),
        .Q(\u2/R1 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [12]),
        .Q(\u2/R1 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [11]),
        .Q(\u2/R1 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [10]),
        .Q(\u2/R1 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [9]),
        .Q(\u2/R1 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [8]),
        .Q(\u2/R1 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [7]),
        .Q(\u2/R1 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [6]),
        .Q(\u2/R1 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [5]),
        .Q(\u2/R1 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [4]),
        .Q(\u2/R1 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [3]),
        .Q(\u2/R1 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [30]),
        .Q(\u2/R1 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [2]),
        .Q(\u2/R1 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [1]),
        .Q(\u2/R1 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [0]),
        .Q(\u2/R1 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [29]),
        .Q(\u2/R1 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [28]),
        .Q(\u2/R1 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [27]),
        .Q(\u2/R1 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [26]),
        .Q(\u2/R1 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [25]),
        .Q(\u2/R1 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [24]),
        .Q(\u2/R1 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R10 [23]),
        .Q(\u2/R1 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[10]_i_1 
       (.I0(\u2/L1 [10]),
        .I1(\u2/out2 [10]),
        .O(\u2/R20 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[11]_i_1 
       (.I0(\u2/L1 [11]),
        .I1(\u2/out2 [11]),
        .O(\u2/R20 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[12]_i_1 
       (.I0(\u2/L1 [12]),
        .I1(\u2/out2 [12]),
        .O(\u2/R20 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[13]_i_1 
       (.I0(\u2/L1 [13]),
        .I1(\u2/out2 [13]),
        .O(\u2/R20 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[14]_i_1 
       (.I0(\u2/L1 [14]),
        .I1(\u2/out2 [14]),
        .O(\u2/R20 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[15]_i_1 
       (.I0(\u2/L1 [15]),
        .I1(\u2/out2 [15]),
        .O(\u2/R20 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[16]_i_1 
       (.I0(\u2/L1 [16]),
        .I1(\u2/out2 [16]),
        .O(\u2/R20 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[17]_i_1 
       (.I0(\u2/L1 [17]),
        .I1(\u2/out2 [17]),
        .O(\u2/R20 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[18]_i_1 
       (.I0(\u2/L1 [18]),
        .I1(\u2/out2 [18]),
        .O(\u2/R20 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[19]_i_1 
       (.I0(\u2/L1 [19]),
        .I1(\u2/out2 [19]),
        .O(\u2/R20 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[1]_i_1 
       (.I0(\u2/L1 [1]),
        .I1(\u2/out2 [1]),
        .O(\u2/R20 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[20]_i_1 
       (.I0(\u2/L1 [20]),
        .I1(\u2/out2 [20]),
        .O(\u2/R20 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[21]_i_1 
       (.I0(\u2/L1 [21]),
        .I1(\u2/out2 [21]),
        .O(\u2/R20 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[22]_i_1 
       (.I0(\u2/L1 [22]),
        .I1(\u2/out2 [22]),
        .O(\u2/R20 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[23]_i_1 
       (.I0(\u2/L1 [23]),
        .I1(\u2/out2 [23]),
        .O(\u2/R20 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[24]_i_1 
       (.I0(\u2/L1 [24]),
        .I1(\u2/out2 [24]),
        .O(\u2/R20 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[25]_i_1 
       (.I0(\u2/L1 [25]),
        .I1(\u2/out2 [25]),
        .O(\u2/R20 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[26]_i_1 
       (.I0(\u2/L1 [26]),
        .I1(\u2/out2 [26]),
        .O(\u2/R20 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[27]_i_1 
       (.I0(\u2/L1 [27]),
        .I1(\u2/out2 [27]),
        .O(\u2/R20 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[28]_i_1 
       (.I0(\u2/L1 [28]),
        .I1(\u2/out2 [28]),
        .O(\u2/R20 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[29]_i_1 
       (.I0(\u2/L1 [29]),
        .I1(\u2/out2 [29]),
        .O(\u2/R20 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[2]_i_1 
       (.I0(\u2/L1 [2]),
        .I1(\u2/out2 [2]),
        .O(\u2/R20 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[30]_i_1 
       (.I0(\u2/L1 [30]),
        .I1(\u2/out2 [30]),
        .O(\u2/R20 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[31]_i_1 
       (.I0(\u2/L1 [31]),
        .I1(\u2/out2 [31]),
        .O(\u2/R20 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[32]_i_1 
       (.I0(\u2/L1 [32]),
        .I1(\u2/out2 [32]),
        .O(\u2/R20 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[3]_i_1 
       (.I0(\u2/L1 [3]),
        .I1(\u2/out2 [3]),
        .O(\u2/R20 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[4]_i_1 
       (.I0(\u2/L1 [4]),
        .I1(\u2/out2 [4]),
        .O(\u2/R20 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[5]_i_1 
       (.I0(\u2/L1 [5]),
        .I1(\u2/out2 [5]),
        .O(\u2/R20 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[6]_i_1 
       (.I0(\u2/L1 [6]),
        .I1(\u2/out2 [6]),
        .O(\u2/R20 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[7]_i_1 
       (.I0(\u2/L1 [7]),
        .I1(\u2/out2 [7]),
        .O(\u2/R20 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[8]_i_1 
       (.I0(\u2/L1 [8]),
        .I1(\u2/out2 [8]),
        .O(\u2/R20 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R2[9]_i_1 
       (.I0(\u2/L1 [9]),
        .I1(\u2/out2 [9]),
        .O(\u2/R20 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [22]),
        .Q(\u2/R2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [21]),
        .Q(\u2/R2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [20]),
        .Q(\u2/R2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [19]),
        .Q(\u2/R2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [18]),
        .Q(\u2/R2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [17]),
        .Q(\u2/R2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [16]),
        .Q(\u2/R2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [15]),
        .Q(\u2/R2 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [14]),
        .Q(\u2/R2 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [13]),
        .Q(\u2/R2 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [31]),
        .Q(\u2/R2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [12]),
        .Q(\u2/R2 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [11]),
        .Q(\u2/R2 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [10]),
        .Q(\u2/R2 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [9]),
        .Q(\u2/R2 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [8]),
        .Q(\u2/R2 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [7]),
        .Q(\u2/R2 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [6]),
        .Q(\u2/R2 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [5]),
        .Q(\u2/R2 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [4]),
        .Q(\u2/R2 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [3]),
        .Q(\u2/R2 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [30]),
        .Q(\u2/R2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [2]),
        .Q(\u2/R2 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [1]),
        .Q(\u2/R2 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [0]),
        .Q(\u2/R2 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [29]),
        .Q(\u2/R2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [28]),
        .Q(\u2/R2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [27]),
        .Q(\u2/R2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [26]),
        .Q(\u2/R2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [25]),
        .Q(\u2/R2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [24]),
        .Q(\u2/R2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R2_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R20 [23]),
        .Q(\u2/R2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[10]_i_1 
       (.I0(\u2/L2 [10]),
        .I1(\u2/out3 [10]),
        .O(\u2/R30 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[11]_i_1 
       (.I0(\u2/L2 [11]),
        .I1(\u2/out3 [11]),
        .O(\u2/R30 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[12]_i_1 
       (.I0(\u2/L2 [12]),
        .I1(\u2/out3 [12]),
        .O(\u2/R30 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[13]_i_1 
       (.I0(\u2/L2 [13]),
        .I1(\u2/out3 [13]),
        .O(\u2/R30 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[14]_i_1 
       (.I0(\u2/L2 [14]),
        .I1(\u2/out3 [14]),
        .O(\u2/R30 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[15]_i_1 
       (.I0(\u2/L2 [15]),
        .I1(\u2/out3 [15]),
        .O(\u2/R30 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[16]_i_1 
       (.I0(\u2/L2 [16]),
        .I1(\u2/out3 [16]),
        .O(\u2/R30 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[17]_i_1 
       (.I0(\u2/L2 [17]),
        .I1(\u2/out3 [17]),
        .O(\u2/R30 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[18]_i_1 
       (.I0(\u2/L2 [18]),
        .I1(\u2/out3 [18]),
        .O(\u2/R30 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[19]_i_1 
       (.I0(\u2/L2 [19]),
        .I1(\u2/out3 [19]),
        .O(\u2/R30 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[1]_i_1 
       (.I0(\u2/L2 [1]),
        .I1(\u2/out3 [1]),
        .O(\u2/R30 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[20]_i_1 
       (.I0(\u2/L2 [20]),
        .I1(\u2/out3 [20]),
        .O(\u2/R30 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[21]_i_1 
       (.I0(\u2/L2 [21]),
        .I1(\u2/out3 [21]),
        .O(\u2/R30 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[22]_i_1 
       (.I0(\u2/L2 [22]),
        .I1(\u2/out3 [22]),
        .O(\u2/R30 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[23]_i_1 
       (.I0(\u2/L2 [23]),
        .I1(\u2/out3 [23]),
        .O(\u2/R30 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[24]_i_1 
       (.I0(\u2/L2 [24]),
        .I1(\u2/out3 [24]),
        .O(\u2/R30 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[25]_i_1 
       (.I0(\u2/L2 [25]),
        .I1(\u2/out3 [25]),
        .O(\u2/R30 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[26]_i_1 
       (.I0(\u2/L2 [26]),
        .I1(\u2/out3 [26]),
        .O(\u2/R30 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[27]_i_1 
       (.I0(\u2/L2 [27]),
        .I1(\u2/out3 [27]),
        .O(\u2/R30 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[28]_i_1 
       (.I0(\u2/L2 [28]),
        .I1(\u2/out3 [28]),
        .O(\u2/R30 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[29]_i_1 
       (.I0(\u2/L2 [29]),
        .I1(\u2/out3 [29]),
        .O(\u2/R30 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[2]_i_1 
       (.I0(\u2/L2 [2]),
        .I1(\u2/out3 [2]),
        .O(\u2/R30 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[30]_i_1 
       (.I0(\u2/L2 [30]),
        .I1(\u2/out3 [30]),
        .O(\u2/R30 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[31]_i_1 
       (.I0(\u2/L2 [31]),
        .I1(\u2/out3 [31]),
        .O(\u2/R30 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[32]_i_1 
       (.I0(\u2/L2 [32]),
        .I1(\u2/out3 [32]),
        .O(\u2/R30 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[3]_i_1 
       (.I0(\u2/L2 [3]),
        .I1(\u2/out3 [3]),
        .O(\u2/R30 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[4]_i_1 
       (.I0(\u2/L2 [4]),
        .I1(\u2/out3 [4]),
        .O(\u2/R30 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[5]_i_1 
       (.I0(\u2/L2 [5]),
        .I1(\u2/out3 [5]),
        .O(\u2/R30 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[6]_i_1 
       (.I0(\u2/L2 [6]),
        .I1(\u2/out3 [6]),
        .O(\u2/R30 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[7]_i_1 
       (.I0(\u2/L2 [7]),
        .I1(\u2/out3 [7]),
        .O(\u2/R30 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[8]_i_1 
       (.I0(\u2/L2 [8]),
        .I1(\u2/out3 [8]),
        .O(\u2/R30 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R3[9]_i_1 
       (.I0(\u2/L2 [9]),
        .I1(\u2/out3 [9]),
        .O(\u2/R30 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [22]),
        .Q(\u2/R3 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [21]),
        .Q(\u2/R3 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [20]),
        .Q(\u2/R3 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [19]),
        .Q(\u2/R3 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [18]),
        .Q(\u2/R3 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [17]),
        .Q(\u2/R3 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [16]),
        .Q(\u2/R3 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [15]),
        .Q(\u2/R3 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [14]),
        .Q(\u2/R3 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [13]),
        .Q(\u2/R3 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [31]),
        .Q(\u2/R3 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [12]),
        .Q(\u2/R3 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [11]),
        .Q(\u2/R3 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [10]),
        .Q(\u2/R3 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [9]),
        .Q(\u2/R3 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [8]),
        .Q(\u2/R3 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [7]),
        .Q(\u2/R3 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [6]),
        .Q(\u2/R3 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [5]),
        .Q(\u2/R3 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [4]),
        .Q(\u2/R3 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [3]),
        .Q(\u2/R3 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [30]),
        .Q(\u2/R3 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [2]),
        .Q(\u2/R3 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [1]),
        .Q(\u2/R3 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [0]),
        .Q(\u2/R3 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [29]),
        .Q(\u2/R3 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [28]),
        .Q(\u2/R3 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [27]),
        .Q(\u2/R3 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [26]),
        .Q(\u2/R3 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [25]),
        .Q(\u2/R3 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [24]),
        .Q(\u2/R3 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R3_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R30 [23]),
        .Q(\u2/R3 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[10]_i_1 
       (.I0(\u2/L3 [10]),
        .I1(\u2/out4 [10]),
        .O(\u2/R40 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[11]_i_1 
       (.I0(\u2/L3 [11]),
        .I1(\u2/out4 [11]),
        .O(\u2/R40 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[12]_i_1 
       (.I0(\u2/L3 [12]),
        .I1(\u2/out4 [12]),
        .O(\u2/R40 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[13]_i_1 
       (.I0(\u2/L3 [13]),
        .I1(\u2/out4 [13]),
        .O(\u2/R40 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[14]_i_1 
       (.I0(\u2/L3 [14]),
        .I1(\u2/out4 [14]),
        .O(\u2/R40 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[15]_i_1 
       (.I0(\u2/L3 [15]),
        .I1(\u2/out4 [15]),
        .O(\u2/R40 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[16]_i_1 
       (.I0(\u2/L3 [16]),
        .I1(\u2/out4 [16]),
        .O(\u2/R40 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[17]_i_1 
       (.I0(\u2/L3 [17]),
        .I1(\u2/out4 [17]),
        .O(\u2/R40 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[18]_i_1 
       (.I0(\u2/L3 [18]),
        .I1(\u2/out4 [18]),
        .O(\u2/R40 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[19]_i_1 
       (.I0(\u2/L3 [19]),
        .I1(\u2/out4 [19]),
        .O(\u2/R40 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[1]_i_1 
       (.I0(\u2/L3 [1]),
        .I1(\u2/out4 [1]),
        .O(\u2/R40 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[20]_i_1 
       (.I0(\u2/L3 [20]),
        .I1(\u2/out4 [20]),
        .O(\u2/R40 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[21]_i_1 
       (.I0(\u2/L3 [21]),
        .I1(\u2/out4 [21]),
        .O(\u2/R40 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[22]_i_1 
       (.I0(\u2/L3 [22]),
        .I1(\u2/out4 [22]),
        .O(\u2/R40 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[23]_i_1 
       (.I0(\u2/L3 [23]),
        .I1(\u2/out4 [23]),
        .O(\u2/R40 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[24]_i_1 
       (.I0(\u2/L3 [24]),
        .I1(\u2/out4 [24]),
        .O(\u2/R40 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[25]_i_1 
       (.I0(\u2/L3 [25]),
        .I1(\u2/out4 [25]),
        .O(\u2/R40 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[26]_i_1 
       (.I0(\u2/L3 [26]),
        .I1(\u2/out4 [26]),
        .O(\u2/R40 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[27]_i_1 
       (.I0(\u2/L3 [27]),
        .I1(\u2/out4 [27]),
        .O(\u2/R40 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[28]_i_1 
       (.I0(\u2/L3 [28]),
        .I1(\u2/out4 [28]),
        .O(\u2/R40 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[29]_i_1 
       (.I0(\u2/L3 [29]),
        .I1(\u2/out4 [29]),
        .O(\u2/R40 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[2]_i_1 
       (.I0(\u2/L3 [2]),
        .I1(\u2/out4 [2]),
        .O(\u2/R40 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[30]_i_1 
       (.I0(\u2/L3 [30]),
        .I1(\u2/out4 [30]),
        .O(\u2/R40 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[31]_i_1 
       (.I0(\u2/L3 [31]),
        .I1(\u2/out4 [31]),
        .O(\u2/R40 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[32]_i_1 
       (.I0(\u2/L3 [32]),
        .I1(\u2/out4 [32]),
        .O(\u2/R40 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[3]_i_1 
       (.I0(\u2/L3 [3]),
        .I1(\u2/out4 [3]),
        .O(\u2/R40 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[4]_i_1 
       (.I0(\u2/L3 [4]),
        .I1(\u2/out4 [4]),
        .O(\u2/R40 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[5]_i_1 
       (.I0(\u2/L3 [5]),
        .I1(\u2/out4 [5]),
        .O(\u2/R40 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[6]_i_1 
       (.I0(\u2/L3 [6]),
        .I1(\u2/out4 [6]),
        .O(\u2/R40 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[7]_i_1 
       (.I0(\u2/L3 [7]),
        .I1(\u2/out4 [7]),
        .O(\u2/R40 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[8]_i_1 
       (.I0(\u2/L3 [8]),
        .I1(\u2/out4 [8]),
        .O(\u2/R40 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R4[9]_i_1 
       (.I0(\u2/L3 [9]),
        .I1(\u2/out4 [9]),
        .O(\u2/R40 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [22]),
        .Q(\u2/R4 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [21]),
        .Q(\u2/R4 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [20]),
        .Q(\u2/R4 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [19]),
        .Q(\u2/R4 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [18]),
        .Q(\u2/R4 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [17]),
        .Q(\u2/R4 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [16]),
        .Q(\u2/R4 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [15]),
        .Q(\u2/R4 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [14]),
        .Q(\u2/R4 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [13]),
        .Q(\u2/R4 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [31]),
        .Q(\u2/R4 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [12]),
        .Q(\u2/R4 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [11]),
        .Q(\u2/R4 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [10]),
        .Q(\u2/R4 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [9]),
        .Q(\u2/R4 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [8]),
        .Q(\u2/R4 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [7]),
        .Q(\u2/R4 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [6]),
        .Q(\u2/R4 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [5]),
        .Q(\u2/R4 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [4]),
        .Q(\u2/R4 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [3]),
        .Q(\u2/R4 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [30]),
        .Q(\u2/R4 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [2]),
        .Q(\u2/R4 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [1]),
        .Q(\u2/R4 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [0]),
        .Q(\u2/R4 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [29]),
        .Q(\u2/R4 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [28]),
        .Q(\u2/R4 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [27]),
        .Q(\u2/R4 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [26]),
        .Q(\u2/R4 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [25]),
        .Q(\u2/R4 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [24]),
        .Q(\u2/R4 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R4_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R40 [23]),
        .Q(\u2/R4 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[10]_i_1 
       (.I0(\u2/L4 [10]),
        .I1(\u2/out5 [10]),
        .O(\u2/R50 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[11]_i_1 
       (.I0(\u2/L4 [11]),
        .I1(\u2/out5 [11]),
        .O(\u2/R50 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[12]_i_1 
       (.I0(\u2/L4 [12]),
        .I1(\u2/out5 [12]),
        .O(\u2/R50 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[13]_i_1 
       (.I0(\u2/L4 [13]),
        .I1(\u2/out5 [13]),
        .O(\u2/R50 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[14]_i_1 
       (.I0(\u2/L4 [14]),
        .I1(\u2/out5 [14]),
        .O(\u2/R50 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[15]_i_1 
       (.I0(\u2/L4 [15]),
        .I1(\u2/out5 [15]),
        .O(\u2/R50 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[16]_i_1 
       (.I0(\u2/L4 [16]),
        .I1(\u2/out5 [16]),
        .O(\u2/R50 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[17]_i_1 
       (.I0(\u2/L4 [17]),
        .I1(\u2/out5 [17]),
        .O(\u2/R50 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[18]_i_1 
       (.I0(\u2/L4 [18]),
        .I1(\u2/out5 [18]),
        .O(\u2/R50 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[19]_i_1 
       (.I0(\u2/L4 [19]),
        .I1(\u2/out5 [19]),
        .O(\u2/R50 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[1]_i_1 
       (.I0(\u2/L4 [1]),
        .I1(\u2/out5 [1]),
        .O(\u2/R50 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[20]_i_1 
       (.I0(\u2/L4 [20]),
        .I1(\u2/out5 [20]),
        .O(\u2/R50 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[21]_i_1 
       (.I0(\u2/L4 [21]),
        .I1(\u2/out5 [21]),
        .O(\u2/R50 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[22]_i_1 
       (.I0(\u2/L4 [22]),
        .I1(\u2/out5 [22]),
        .O(\u2/R50 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[23]_i_1 
       (.I0(\u2/L4 [23]),
        .I1(\u2/out5 [23]),
        .O(\u2/R50 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[24]_i_1 
       (.I0(\u2/L4 [24]),
        .I1(\u2/out5 [24]),
        .O(\u2/R50 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[25]_i_1 
       (.I0(\u2/L4 [25]),
        .I1(\u2/out5 [25]),
        .O(\u2/R50 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[26]_i_1 
       (.I0(\u2/L4 [26]),
        .I1(\u2/out5 [26]),
        .O(\u2/R50 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[27]_i_1 
       (.I0(\u2/L4 [27]),
        .I1(\u2/out5 [27]),
        .O(\u2/R50 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[28]_i_1 
       (.I0(\u2/L4 [28]),
        .I1(\u2/out5 [28]),
        .O(\u2/R50 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[29]_i_1 
       (.I0(\u2/L4 [29]),
        .I1(\u2/out5 [29]),
        .O(\u2/R50 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[2]_i_1 
       (.I0(\u2/L4 [2]),
        .I1(\u2/out5 [2]),
        .O(\u2/R50 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[30]_i_1 
       (.I0(\u2/L4 [30]),
        .I1(\u2/out5 [30]),
        .O(\u2/R50 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[31]_i_1 
       (.I0(\u2/L4 [31]),
        .I1(\u2/out5 [31]),
        .O(\u2/R50 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[32]_i_1 
       (.I0(\u2/L4 [32]),
        .I1(\u2/out5 [32]),
        .O(\u2/R50 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[3]_i_1 
       (.I0(\u2/L4 [3]),
        .I1(\u2/out5 [3]),
        .O(\u2/R50 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[4]_i_1 
       (.I0(\u2/L4 [4]),
        .I1(\u2/out5 [4]),
        .O(\u2/R50 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[5]_i_1 
       (.I0(\u2/L4 [5]),
        .I1(\u2/out5 [5]),
        .O(\u2/R50 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[6]_i_1 
       (.I0(\u2/L4 [6]),
        .I1(\u2/out5 [6]),
        .O(\u2/R50 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[7]_i_1 
       (.I0(\u2/L4 [7]),
        .I1(\u2/out5 [7]),
        .O(\u2/R50 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[8]_i_1 
       (.I0(\u2/L4 [8]),
        .I1(\u2/out5 [8]),
        .O(\u2/R50 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R5[9]_i_1 
       (.I0(\u2/L4 [9]),
        .I1(\u2/out5 [9]),
        .O(\u2/R50 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [22]),
        .Q(\u2/R5 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [21]),
        .Q(\u2/R5 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [20]),
        .Q(\u2/R5 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [19]),
        .Q(\u2/R5 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [18]),
        .Q(\u2/R5 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [17]),
        .Q(\u2/R5 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [16]),
        .Q(\u2/R5 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [15]),
        .Q(\u2/R5 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [14]),
        .Q(\u2/R5 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [13]),
        .Q(\u2/R5 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [31]),
        .Q(\u2/R5 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [12]),
        .Q(\u2/R5 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [11]),
        .Q(\u2/R5 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [10]),
        .Q(\u2/R5 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [9]),
        .Q(\u2/R5 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [8]),
        .Q(\u2/R5 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [7]),
        .Q(\u2/R5 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [6]),
        .Q(\u2/R5 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [5]),
        .Q(\u2/R5 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [4]),
        .Q(\u2/R5 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [3]),
        .Q(\u2/R5 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [30]),
        .Q(\u2/R5 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [2]),
        .Q(\u2/R5 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [1]),
        .Q(\u2/R5 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [0]),
        .Q(\u2/R5 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [29]),
        .Q(\u2/R5 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [28]),
        .Q(\u2/R5 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [27]),
        .Q(\u2/R5 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [26]),
        .Q(\u2/R5 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [25]),
        .Q(\u2/R5 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [24]),
        .Q(\u2/R5 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R5_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R50 [23]),
        .Q(\u2/R5 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[10]_i_1 
       (.I0(\u2/L5 [10]),
        .I1(\u2/out6 [10]),
        .O(\u2/R60 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[11]_i_1 
       (.I0(\u2/L5 [11]),
        .I1(\u2/out6 [11]),
        .O(\u2/R60 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[12]_i_1 
       (.I0(\u2/L5 [12]),
        .I1(\u2/out6 [12]),
        .O(\u2/R60 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[13]_i_1 
       (.I0(\u2/L5 [13]),
        .I1(\u2/out6 [13]),
        .O(\u2/R60 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[14]_i_1 
       (.I0(\u2/L5 [14]),
        .I1(\u2/out6 [14]),
        .O(\u2/R60 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[15]_i_1 
       (.I0(\u2/L5 [15]),
        .I1(\u2/out6 [15]),
        .O(\u2/R60 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[16]_i_1 
       (.I0(\u2/L5 [16]),
        .I1(\u2/out6 [16]),
        .O(\u2/R60 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[17]_i_1 
       (.I0(\u2/L5 [17]),
        .I1(\u2/out6 [17]),
        .O(\u2/R60 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[18]_i_1 
       (.I0(\u2/L5 [18]),
        .I1(\u2/out6 [18]),
        .O(\u2/R60 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[19]_i_1 
       (.I0(\u2/L5 [19]),
        .I1(\u2/out6 [19]),
        .O(\u2/R60 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[1]_i_1 
       (.I0(\u2/L5 [1]),
        .I1(\u2/out6 [1]),
        .O(\u2/R60 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[20]_i_1 
       (.I0(\u2/L5 [20]),
        .I1(\u2/out6 [20]),
        .O(\u2/R60 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[21]_i_1 
       (.I0(\u2/L5 [21]),
        .I1(\u2/out6 [21]),
        .O(\u2/R60 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[22]_i_1 
       (.I0(\u2/L5 [22]),
        .I1(\u2/out6 [22]),
        .O(\u2/R60 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[23]_i_1 
       (.I0(\u2/L5 [23]),
        .I1(\u2/out6 [23]),
        .O(\u2/R60 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[24]_i_1 
       (.I0(\u2/L5 [24]),
        .I1(\u2/out6 [24]),
        .O(\u2/R60 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[25]_i_1 
       (.I0(\u2/L5 [25]),
        .I1(\u2/out6 [25]),
        .O(\u2/R60 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[26]_i_1 
       (.I0(\u2/L5 [26]),
        .I1(\u2/out6 [26]),
        .O(\u2/R60 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[27]_i_1 
       (.I0(\u2/L5 [27]),
        .I1(\u2/out6 [27]),
        .O(\u2/R60 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[28]_i_1 
       (.I0(\u2/L5 [28]),
        .I1(\u2/out6 [28]),
        .O(\u2/R60 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[29]_i_1 
       (.I0(\u2/L5 [29]),
        .I1(\u2/out6 [29]),
        .O(\u2/R60 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[2]_i_1 
       (.I0(\u2/L5 [2]),
        .I1(\u2/out6 [2]),
        .O(\u2/R60 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[30]_i_1 
       (.I0(\u2/L5 [30]),
        .I1(\u2/out6 [30]),
        .O(\u2/R60 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[31]_i_1 
       (.I0(\u2/L5 [31]),
        .I1(\u2/out6 [31]),
        .O(\u2/R60 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[32]_i_1 
       (.I0(\u2/L5 [32]),
        .I1(\u2/out6 [32]),
        .O(\u2/R60 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[3]_i_1 
       (.I0(\u2/L5 [3]),
        .I1(\u2/out6 [3]),
        .O(\u2/R60 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[4]_i_1 
       (.I0(\u2/L5 [4]),
        .I1(\u2/out6 [4]),
        .O(\u2/R60 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[5]_i_1 
       (.I0(\u2/L5 [5]),
        .I1(\u2/out6 [5]),
        .O(\u2/R60 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[6]_i_1 
       (.I0(\u2/L5 [6]),
        .I1(\u2/out6 [6]),
        .O(\u2/R60 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[7]_i_1 
       (.I0(\u2/L5 [7]),
        .I1(\u2/out6 [7]),
        .O(\u2/R60 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[8]_i_1 
       (.I0(\u2/L5 [8]),
        .I1(\u2/out6 [8]),
        .O(\u2/R60 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R6[9]_i_1 
       (.I0(\u2/L5 [9]),
        .I1(\u2/out6 [9]),
        .O(\u2/R60 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [22]),
        .Q(\u2/R6 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [21]),
        .Q(\u2/R6 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [20]),
        .Q(\u2/R6 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [19]),
        .Q(\u2/R6 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [18]),
        .Q(\u2/R6 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [17]),
        .Q(\u2/R6 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [16]),
        .Q(\u2/R6 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [15]),
        .Q(\u2/R6 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [14]),
        .Q(\u2/R6 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [13]),
        .Q(\u2/R6 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [31]),
        .Q(\u2/R6 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [12]),
        .Q(\u2/R6 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [11]),
        .Q(\u2/R6 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [10]),
        .Q(\u2/R6 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [9]),
        .Q(\u2/R6 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [8]),
        .Q(\u2/R6 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [7]),
        .Q(\u2/R6 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [6]),
        .Q(\u2/R6 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [5]),
        .Q(\u2/R6 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [4]),
        .Q(\u2/R6 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [3]),
        .Q(\u2/R6 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [30]),
        .Q(\u2/R6 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [2]),
        .Q(\u2/R6 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [1]),
        .Q(\u2/R6 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [0]),
        .Q(\u2/R6 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [29]),
        .Q(\u2/R6 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [28]),
        .Q(\u2/R6 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [27]),
        .Q(\u2/R6 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [26]),
        .Q(\u2/R6 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [25]),
        .Q(\u2/R6 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [24]),
        .Q(\u2/R6 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R6_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R60 [23]),
        .Q(\u2/R6 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[10]_i_1 
       (.I0(\u2/L6 [10]),
        .I1(\u2/out7 [10]),
        .O(\u2/R70 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[11]_i_1 
       (.I0(\u2/L6 [11]),
        .I1(\u2/out7 [11]),
        .O(\u2/R70 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[12]_i_1 
       (.I0(\u2/L6 [12]),
        .I1(\u2/out7 [12]),
        .O(\u2/R70 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[13]_i_1 
       (.I0(\u2/L6 [13]),
        .I1(\u2/out7 [13]),
        .O(\u2/R70 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[14]_i_1 
       (.I0(\u2/L6 [14]),
        .I1(\u2/out7 [14]),
        .O(\u2/R70 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[15]_i_1 
       (.I0(\u2/L6 [15]),
        .I1(\u2/out7 [15]),
        .O(\u2/R70 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[16]_i_1 
       (.I0(\u2/L6 [16]),
        .I1(\u2/out7 [16]),
        .O(\u2/R70 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[17]_i_1 
       (.I0(\u2/L6 [17]),
        .I1(\u2/out7 [17]),
        .O(\u2/R70 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[18]_i_1 
       (.I0(\u2/L6 [18]),
        .I1(\u2/out7 [18]),
        .O(\u2/R70 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[19]_i_1 
       (.I0(\u2/L6 [19]),
        .I1(\u2/out7 [19]),
        .O(\u2/R70 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[1]_i_1 
       (.I0(\u2/L6 [1]),
        .I1(\u2/out7 [1]),
        .O(\u2/R70 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[20]_i_1 
       (.I0(\u2/L6 [20]),
        .I1(\u2/out7 [20]),
        .O(\u2/R70 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[21]_i_1 
       (.I0(\u2/L6 [21]),
        .I1(\u2/out7 [21]),
        .O(\u2/R70 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[22]_i_1 
       (.I0(\u2/L6 [22]),
        .I1(\u2/out7 [22]),
        .O(\u2/R70 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[23]_i_1 
       (.I0(\u2/L6 [23]),
        .I1(\u2/out7 [23]),
        .O(\u2/R70 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[24]_i_1 
       (.I0(\u2/L6 [24]),
        .I1(\u2/out7 [24]),
        .O(\u2/R70 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[25]_i_1 
       (.I0(\u2/L6 [25]),
        .I1(\u2/out7 [25]),
        .O(\u2/R70 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[26]_i_1 
       (.I0(\u2/L6 [26]),
        .I1(\u2/out7 [26]),
        .O(\u2/R70 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[27]_i_1 
       (.I0(\u2/L6 [27]),
        .I1(\u2/out7 [27]),
        .O(\u2/R70 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[28]_i_1 
       (.I0(\u2/L6 [28]),
        .I1(\u2/out7 [28]),
        .O(\u2/R70 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[29]_i_1 
       (.I0(\u2/L6 [29]),
        .I1(\u2/out7 [29]),
        .O(\u2/R70 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[2]_i_1 
       (.I0(\u2/L6 [2]),
        .I1(\u2/out7 [2]),
        .O(\u2/R70 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[30]_i_1 
       (.I0(\u2/L6 [30]),
        .I1(\u2/out7 [30]),
        .O(\u2/R70 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[31]_i_1 
       (.I0(\u2/L6 [31]),
        .I1(\u2/out7 [31]),
        .O(\u2/R70 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[32]_i_1 
       (.I0(\u2/L6 [32]),
        .I1(\u2/out7 [32]),
        .O(\u2/R70 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[3]_i_1 
       (.I0(\u2/L6 [3]),
        .I1(\u2/out7 [3]),
        .O(\u2/R70 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[4]_i_1 
       (.I0(\u2/L6 [4]),
        .I1(\u2/out7 [4]),
        .O(\u2/R70 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[5]_i_1 
       (.I0(\u2/L6 [5]),
        .I1(\u2/out7 [5]),
        .O(\u2/R70 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[6]_i_1 
       (.I0(\u2/L6 [6]),
        .I1(\u2/out7 [6]),
        .O(\u2/R70 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[7]_i_1 
       (.I0(\u2/L6 [7]),
        .I1(\u2/out7 [7]),
        .O(\u2/R70 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[8]_i_1 
       (.I0(\u2/L6 [8]),
        .I1(\u2/out7 [8]),
        .O(\u2/R70 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R7[9]_i_1 
       (.I0(\u2/L6 [9]),
        .I1(\u2/out7 [9]),
        .O(\u2/R70 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [22]),
        .Q(\u2/R7 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [21]),
        .Q(\u2/R7 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [20]),
        .Q(\u2/R7 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [19]),
        .Q(\u2/R7 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [18]),
        .Q(\u2/R7 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [17]),
        .Q(\u2/R7 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [16]),
        .Q(\u2/R7 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [15]),
        .Q(\u2/R7 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [14]),
        .Q(\u2/R7 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [13]),
        .Q(\u2/R7 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [31]),
        .Q(\u2/R7 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [12]),
        .Q(\u2/R7 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [11]),
        .Q(\u2/R7 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [10]),
        .Q(\u2/R7 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [9]),
        .Q(\u2/R7 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [8]),
        .Q(\u2/R7 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [7]),
        .Q(\u2/R7 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [6]),
        .Q(\u2/R7 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [5]),
        .Q(\u2/R7 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [4]),
        .Q(\u2/R7 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [3]),
        .Q(\u2/R7 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [30]),
        .Q(\u2/R7 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [2]),
        .Q(\u2/R7 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [1]),
        .Q(\u2/R7 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [0]),
        .Q(\u2/R7 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [29]),
        .Q(\u2/R7 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [28]),
        .Q(\u2/R7 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [27]),
        .Q(\u2/R7 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [26]),
        .Q(\u2/R7 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [25]),
        .Q(\u2/R7 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [24]),
        .Q(\u2/R7 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R7_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R70 [23]),
        .Q(\u2/R7 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[10]_i_1 
       (.I0(\u2/L7 [10]),
        .I1(\u2/out8 [10]),
        .O(\u2/R80 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[11]_i_1 
       (.I0(\u2/L7 [11]),
        .I1(\u2/out8 [11]),
        .O(\u2/R80 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[12]_i_1 
       (.I0(\u2/L7 [12]),
        .I1(\u2/out8 [12]),
        .O(\u2/R80 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[13]_i_1 
       (.I0(\u2/L7 [13]),
        .I1(\u2/out8 [13]),
        .O(\u2/R80 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[14]_i_1 
       (.I0(\u2/L7 [14]),
        .I1(\u2/out8 [14]),
        .O(\u2/R80 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[15]_i_1 
       (.I0(\u2/L7 [15]),
        .I1(\u2/out8 [15]),
        .O(\u2/R80 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[16]_i_1 
       (.I0(\u2/L7 [16]),
        .I1(\u2/out8 [16]),
        .O(\u2/R80 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[17]_i_1 
       (.I0(\u2/L7 [17]),
        .I1(\u2/out8 [17]),
        .O(\u2/R80 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[18]_i_1 
       (.I0(\u2/L7 [18]),
        .I1(\u2/out8 [18]),
        .O(\u2/R80 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[19]_i_1 
       (.I0(\u2/L7 [19]),
        .I1(\u2/out8 [19]),
        .O(\u2/R80 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[1]_i_1 
       (.I0(\u2/L7 [1]),
        .I1(\u2/out8 [1]),
        .O(\u2/R80 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[20]_i_1 
       (.I0(\u2/L7 [20]),
        .I1(\u2/out8 [20]),
        .O(\u2/R80 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[21]_i_1 
       (.I0(\u2/L7 [21]),
        .I1(\u2/out8 [21]),
        .O(\u2/R80 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[22]_i_1 
       (.I0(\u2/L7 [22]),
        .I1(\u2/out8 [22]),
        .O(\u2/R80 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[23]_i_1 
       (.I0(\u2/L7 [23]),
        .I1(\u2/out8 [23]),
        .O(\u2/R80 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[24]_i_1 
       (.I0(\u2/L7 [24]),
        .I1(\u2/out8 [24]),
        .O(\u2/R80 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[25]_i_1 
       (.I0(\u2/L7 [25]),
        .I1(\u2/out8 [25]),
        .O(\u2/R80 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[26]_i_1 
       (.I0(\u2/L7 [26]),
        .I1(\u2/out8 [26]),
        .O(\u2/R80 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[27]_i_1 
       (.I0(\u2/L7 [27]),
        .I1(\u2/out8 [27]),
        .O(\u2/R80 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[28]_i_1 
       (.I0(\u2/L7 [28]),
        .I1(\u2/out8 [28]),
        .O(\u2/R80 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[29]_i_1 
       (.I0(\u2/L7 [29]),
        .I1(\u2/out8 [29]),
        .O(\u2/R80 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[2]_i_1 
       (.I0(\u2/L7 [2]),
        .I1(\u2/out8 [2]),
        .O(\u2/R80 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[30]_i_1 
       (.I0(\u2/L7 [30]),
        .I1(\u2/out8 [30]),
        .O(\u2/R80 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[31]_i_1 
       (.I0(\u2/L7 [31]),
        .I1(\u2/out8 [31]),
        .O(\u2/R80 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[32]_i_1 
       (.I0(\u2/L7 [32]),
        .I1(\u2/out8 [32]),
        .O(\u2/R80 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[3]_i_1 
       (.I0(\u2/L7 [3]),
        .I1(\u2/out8 [3]),
        .O(\u2/R80 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[4]_i_1 
       (.I0(\u2/L7 [4]),
        .I1(\u2/out8 [4]),
        .O(\u2/R80 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[5]_i_1 
       (.I0(\u2/L7 [5]),
        .I1(\u2/out8 [5]),
        .O(\u2/R80 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[6]_i_1 
       (.I0(\u2/L7 [6]),
        .I1(\u2/out8 [6]),
        .O(\u2/R80 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[7]_i_1 
       (.I0(\u2/L7 [7]),
        .I1(\u2/out8 [7]),
        .O(\u2/R80 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[8]_i_1 
       (.I0(\u2/L7 [8]),
        .I1(\u2/out8 [8]),
        .O(\u2/R80 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R8[9]_i_1 
       (.I0(\u2/L7 [9]),
        .I1(\u2/out8 [9]),
        .O(\u2/R80 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [22]),
        .Q(\u2/R8 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [21]),
        .Q(\u2/R8 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [20]),
        .Q(\u2/R8 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [19]),
        .Q(\u2/R8 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [18]),
        .Q(\u2/R8 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [17]),
        .Q(\u2/R8 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [16]),
        .Q(\u2/R8 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [15]),
        .Q(\u2/R8 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [14]),
        .Q(\u2/R8 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [13]),
        .Q(\u2/R8 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [31]),
        .Q(\u2/R8 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [12]),
        .Q(\u2/R8 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [11]),
        .Q(\u2/R8 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [10]),
        .Q(\u2/R8 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [9]),
        .Q(\u2/R8 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [8]),
        .Q(\u2/R8 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [7]),
        .Q(\u2/R8 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [6]),
        .Q(\u2/R8 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [5]),
        .Q(\u2/R8 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [4]),
        .Q(\u2/R8 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [3]),
        .Q(\u2/R8 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [30]),
        .Q(\u2/R8 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [2]),
        .Q(\u2/R8 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [1]),
        .Q(\u2/R8 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [0]),
        .Q(\u2/R8 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [29]),
        .Q(\u2/R8 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [28]),
        .Q(\u2/R8 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [27]),
        .Q(\u2/R8 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [26]),
        .Q(\u2/R8 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [25]),
        .Q(\u2/R8 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [24]),
        .Q(\u2/R8 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R8_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R80 [23]),
        .Q(\u2/R8 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[10]_i_1 
       (.I0(\u2/L8 [10]),
        .I1(\u2/out9 [10]),
        .O(\u2/R90 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[11]_i_1 
       (.I0(\u2/L8 [11]),
        .I1(\u2/out9 [11]),
        .O(\u2/R90 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[12]_i_1 
       (.I0(\u2/L8 [12]),
        .I1(\u2/out9 [12]),
        .O(\u2/R90 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[13]_i_1 
       (.I0(\u2/L8 [13]),
        .I1(\u2/out9 [13]),
        .O(\u2/R90 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[14]_i_1 
       (.I0(\u2/L8 [14]),
        .I1(\u2/out9 [14]),
        .O(\u2/R90 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[15]_i_1 
       (.I0(\u2/L8 [15]),
        .I1(\u2/out9 [15]),
        .O(\u2/R90 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[16]_i_1 
       (.I0(\u2/L8 [16]),
        .I1(\u2/out9 [16]),
        .O(\u2/R90 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[17]_i_1 
       (.I0(\u2/L8 [17]),
        .I1(\u2/out9 [17]),
        .O(\u2/R90 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[18]_i_1 
       (.I0(\u2/L8 [18]),
        .I1(\u2/out9 [18]),
        .O(\u2/R90 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[19]_i_1 
       (.I0(\u2/L8 [19]),
        .I1(\u2/out9 [19]),
        .O(\u2/R90 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[1]_i_1 
       (.I0(\u2/L8 [1]),
        .I1(\u2/out9 [1]),
        .O(\u2/R90 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[20]_i_1 
       (.I0(\u2/L8 [20]),
        .I1(\u2/out9 [20]),
        .O(\u2/R90 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[21]_i_1 
       (.I0(\u2/L8 [21]),
        .I1(\u2/out9 [21]),
        .O(\u2/R90 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[22]_i_1 
       (.I0(\u2/L8 [22]),
        .I1(\u2/out9 [22]),
        .O(\u2/R90 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[23]_i_1 
       (.I0(\u2/L8 [23]),
        .I1(\u2/out9 [23]),
        .O(\u2/R90 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[24]_i_1 
       (.I0(\u2/L8 [24]),
        .I1(\u2/out9 [24]),
        .O(\u2/R90 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[25]_i_1 
       (.I0(\u2/L8 [25]),
        .I1(\u2/out9 [25]),
        .O(\u2/R90 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[26]_i_1 
       (.I0(\u2/L8 [26]),
        .I1(\u2/out9 [26]),
        .O(\u2/R90 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[27]_i_1 
       (.I0(\u2/L8 [27]),
        .I1(\u2/out9 [27]),
        .O(\u2/R90 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[28]_i_1 
       (.I0(\u2/L8 [28]),
        .I1(\u2/out9 [28]),
        .O(\u2/R90 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[29]_i_1 
       (.I0(\u2/L8 [29]),
        .I1(\u2/out9 [29]),
        .O(\u2/R90 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[2]_i_1 
       (.I0(\u2/L8 [2]),
        .I1(\u2/out9 [2]),
        .O(\u2/R90 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[30]_i_1 
       (.I0(\u2/L8 [30]),
        .I1(\u2/out9 [30]),
        .O(\u2/R90 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[31]_i_1 
       (.I0(\u2/L8 [31]),
        .I1(\u2/out9 [31]),
        .O(\u2/R90 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[32]_i_1 
       (.I0(\u2/L8 [32]),
        .I1(\u2/out9 [32]),
        .O(\u2/R90 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[3]_i_1 
       (.I0(\u2/L8 [3]),
        .I1(\u2/out9 [3]),
        .O(\u2/R90 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[4]_i_1 
       (.I0(\u2/L8 [4]),
        .I1(\u2/out9 [4]),
        .O(\u2/R90 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[5]_i_1 
       (.I0(\u2/L8 [5]),
        .I1(\u2/out9 [5]),
        .O(\u2/R90 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[6]_i_1 
       (.I0(\u2/L8 [6]),
        .I1(\u2/out9 [6]),
        .O(\u2/R90 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[7]_i_1 
       (.I0(\u2/L8 [7]),
        .I1(\u2/out9 [7]),
        .O(\u2/R90 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[8]_i_1 
       (.I0(\u2/L8 [8]),
        .I1(\u2/out9 [8]),
        .O(\u2/R90 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/R9[9]_i_1 
       (.I0(\u2/L8 [9]),
        .I1(\u2/out9 [9]),
        .O(\u2/R90 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [22]),
        .Q(\u2/R9 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [21]),
        .Q(\u2/R9 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [20]),
        .Q(\u2/R9 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [19]),
        .Q(\u2/R9 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [18]),
        .Q(\u2/R9 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [17]),
        .Q(\u2/R9 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [16]),
        .Q(\u2/R9 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [15]),
        .Q(\u2/R9 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [14]),
        .Q(\u2/R9 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [13]),
        .Q(\u2/R9 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [31]),
        .Q(\u2/R9 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [12]),
        .Q(\u2/R9 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [11]),
        .Q(\u2/R9 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [10]),
        .Q(\u2/R9 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [9]),
        .Q(\u2/R9 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [8]),
        .Q(\u2/R9 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [7]),
        .Q(\u2/R9 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [6]),
        .Q(\u2/R9 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [5]),
        .Q(\u2/R9 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [4]),
        .Q(\u2/R9 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [3]),
        .Q(\u2/R9 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [30]),
        .Q(\u2/R9 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [2]),
        .Q(\u2/R9 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [1]),
        .Q(\u2/R9 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [0]),
        .Q(\u2/R9 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [29]),
        .Q(\u2/R9 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [28]),
        .Q(\u2/R9 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [27]),
        .Q(\u2/R9 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [26]),
        .Q(\u2/R9 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [25]),
        .Q(\u2/R9 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [24]),
        .Q(\u2/R9 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/R9_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/R90 [23]),
        .Q(\u2/R9 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[0]),
        .Q(\u2/IP [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[10]),
        .Q(\u2/IP [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[11]),
        .Q(\u2/IP [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[12]),
        .Q(\u2/IP [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[13]),
        .Q(\u2/IP [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[14]),
        .Q(\u2/IP [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[15]),
        .Q(\u2/IP [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[16]),
        .Q(\u2/IP [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[17]),
        .Q(\u2/IP [59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[18]),
        .Q(\u2/IP [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[19]),
        .Q(\u2/IP [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[1]),
        .Q(\u2/IP [57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[20]),
        .Q(\u2/IP [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[21]),
        .Q(\u2/IP [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[22]),
        .Q(\u2/IP [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[23]),
        .Q(\u2/IP [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[24]),
        .Q(\u2/IP [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[25]),
        .Q(\u2/IP [60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[26]),
        .Q(\u2/IP [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[27]),
        .Q(\u2/IP [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[28]),
        .Q(\u2/IP [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[29]),
        .Q(\u2/IP [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[2]),
        .Q(\u2/IP [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[30]),
        .Q(\u2/IP [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[31]),
        .Q(\u2/IP [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[32]),
        .Q(\u2/IP [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[33]),
        .Q(\u2/IP [61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[34]),
        .Q(\u2/IP [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[35]),
        .Q(\u2/IP [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[36]),
        .Q(\u2/IP [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[37]),
        .Q(\u2/IP [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[38]),
        .Q(\u2/IP [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[39]),
        .Q(\u2/IP [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[3]),
        .Q(\u2/IP [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[40]),
        .Q(\u2/IP [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[41]),
        .Q(\u2/IP [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[42]),
        .Q(\u2/IP [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[43]),
        .Q(\u2/IP [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[44]),
        .Q(\u2/IP [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[45]),
        .Q(\u2/IP [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[46]),
        .Q(\u2/IP [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[47]),
        .Q(\u2/IP [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[48]),
        .Q(\u2/IP [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[49]),
        .Q(\u2/IP [63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[4]),
        .Q(\u2/IP [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[50]),
        .Q(\u2/IP [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[51]),
        .Q(\u2/IP [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[52]),
        .Q(\u2/IP [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[53]),
        .Q(\u2/IP [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[54]),
        .Q(\u2/IP [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[55]),
        .Q(\u2/IP [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[56]),
        .Q(\u2/IP [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[57]),
        .Q(\u2/IP [64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[58]),
        .Q(\u2/IP [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[59]),
        .Q(\u2/IP [56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[5]),
        .Q(\u2/IP [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[60]),
        .Q(\u2/IP [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[61]),
        .Q(\u2/IP [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[62]),
        .Q(\u2/IP [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[63]),
        .Q(\u2/IP [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[6]),
        .Q(\u2/IP [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[7]),
        .Q(\u2/IP [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[8]),
        .Q(\u2/IP [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desIn_r_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(stage2_out[9]),
        .Q(\u2/IP [58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[0]_i_1 
       (.I0(\u2/out15 [25]),
        .I1(\u2/L14 [25]),
        .O(\u2/FP [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[10]_i_1 
       (.I0(\u2/out15 [18]),
        .I1(\u2/L14 [18]),
        .O(\u2/FP [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[12]_i_1 
       (.I0(\u2/out15 [10]),
        .I1(\u2/L14 [10]),
        .O(\u2/FP [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[14]_i_1 
       (.I0(\u2/out15 [2]),
        .I1(\u2/L14 [2]),
        .O(\u2/FP [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[16]_i_1 
       (.I0(\u2/out15 [27]),
        .I1(\u2/L14 [27]),
        .O(\u2/FP [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[18]_i_1 
       (.I0(\u2/out15 [19]),
        .I1(\u2/L14 [19]),
        .O(\u2/FP [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[20]_i_1 
       (.I0(\u2/out15 [11]),
        .I1(\u2/L14 [11]),
        .O(\u2/FP [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[22]_i_1 
       (.I0(\u2/out15 [3]),
        .I1(\u2/L14 [3]),
        .O(\u2/FP [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[24]_i_1 
       (.I0(\u2/out15 [28]),
        .I1(\u2/L14 [28]),
        .O(\u2/FP [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[26]_i_1 
       (.I0(\u2/out15 [20]),
        .I1(\u2/L14 [20]),
        .O(\u2/FP [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[28]_i_1 
       (.I0(\u2/out15 [12]),
        .I1(\u2/L14 [12]),
        .O(\u2/FP [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[2]_i_1 
       (.I0(\u2/out15 [17]),
        .I1(\u2/L14 [17]),
        .O(\u2/FP [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[30]_i_1 
       (.I0(\u2/out15 [4]),
        .I1(\u2/L14 [4]),
        .O(\u2/FP [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[32]_i_1 
       (.I0(\u2/out15 [29]),
        .I1(\u2/L14 [29]),
        .O(\u2/FP [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[34]_i_1 
       (.I0(\u2/out15 [21]),
        .I1(\u2/L14 [21]),
        .O(\u2/FP [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[36]_i_1 
       (.I0(\u2/out15 [13]),
        .I1(\u2/L14 [13]),
        .O(\u2/FP [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[38]_i_1 
       (.I0(\u2/out15 [5]),
        .I1(\u2/L14 [5]),
        .O(\u2/FP [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[40]_i_1 
       (.I0(\u2/out15 [30]),
        .I1(\u2/L14 [30]),
        .O(\u2/FP [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[42]_i_1 
       (.I0(\u2/out15 [22]),
        .I1(\u2/L14 [22]),
        .O(\u2/FP [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[44]_i_1 
       (.I0(\u2/out15 [14]),
        .I1(\u2/L14 [14]),
        .O(\u2/FP [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[46]_i_1 
       (.I0(\u2/out15 [6]),
        .I1(\u2/L14 [6]),
        .O(\u2/FP [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[48]_i_1 
       (.I0(\u2/out15 [31]),
        .I1(\u2/L14 [31]),
        .O(\u2/FP [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[4]_i_1 
       (.I0(\u2/out15 [9]),
        .I1(\u2/L14 [9]),
        .O(\u2/FP [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[50]_i_1 
       (.I0(\u2/out15 [23]),
        .I1(\u2/L14 [23]),
        .O(\u2/FP [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[52]_i_1 
       (.I0(\u2/out15 [15]),
        .I1(\u2/L14 [15]),
        .O(\u2/FP [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[54]_i_1 
       (.I0(\u2/out15 [7]),
        .I1(\u2/L14 [7]),
        .O(\u2/FP [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[56]_i_1 
       (.I0(\u2/out15 [32]),
        .I1(\u2/L14 [32]),
        .O(\u2/FP [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[58]_i_1 
       (.I0(\u2/out15 [24]),
        .I1(\u2/L14 [24]),
        .O(\u2/FP [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[60]_i_1 
       (.I0(\u2/out15 [16]),
        .I1(\u2/L14 [16]),
        .O(\u2/FP [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[62]_i_1 
       (.I0(\u2/out15 [8]),
        .I1(\u2/L14 [8]),
        .O(\u2/FP [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[6]_i_1 
       (.I0(\u2/out15 [1]),
        .I1(\u2/L14 [1]),
        .O(\u2/FP [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \u2/desOut[8]_i_1 
       (.I0(\u2/out15 [26]),
        .I1(\u2/L14 [26]),
        .O(\u2/FP [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [25]),
        .Q(desOut[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [18]),
        .Q(desOut[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [50]),
        .Q(desOut[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [10]),
        .Q(desOut[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [42]),
        .Q(desOut[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [2]),
        .Q(desOut[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [34]),
        .Q(desOut[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [27]),
        .Q(desOut[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [59]),
        .Q(desOut[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [19]),
        .Q(desOut[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [51]),
        .Q(desOut[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [57]),
        .Q(desOut[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [11]),
        .Q(desOut[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [43]),
        .Q(desOut[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [3]),
        .Q(desOut[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [35]),
        .Q(desOut[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [28]),
        .Q(desOut[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [60]),
        .Q(desOut[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [20]),
        .Q(desOut[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [52]),
        .Q(desOut[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [12]),
        .Q(desOut[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [44]),
        .Q(desOut[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [17]),
        .Q(desOut[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [4]),
        .Q(desOut[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [36]),
        .Q(desOut[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [29]),
        .Q(desOut[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [61]),
        .Q(desOut[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [21]),
        .Q(desOut[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [53]),
        .Q(desOut[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [13]),
        .Q(desOut[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [45]),
        .Q(desOut[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [5]),
        .Q(desOut[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [37]),
        .Q(desOut[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [49]),
        .Q(desOut[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [30]),
        .Q(desOut[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [62]),
        .Q(desOut[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [22]),
        .Q(desOut[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [54]),
        .Q(desOut[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [14]),
        .Q(desOut[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [46]),
        .Q(desOut[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [6]),
        .Q(desOut[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [38]),
        .Q(desOut[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [31]),
        .Q(desOut[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [63]),
        .Q(desOut[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [9]),
        .Q(desOut[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [23]),
        .Q(desOut[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [55]),
        .Q(desOut[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [15]),
        .Q(desOut[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [47]),
        .Q(desOut[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [7]),
        .Q(desOut[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [39]),
        .Q(desOut[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [32]),
        .Q(desOut[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [64]),
        .Q(desOut[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [24]),
        .Q(desOut[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [56]),
        .Q(desOut[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [41]),
        .Q(desOut[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [16]),
        .Q(desOut[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [48]),
        .Q(desOut[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [8]),
        .Q(desOut[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [40]),
        .Q(desOut[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [1]),
        .Q(desOut[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [33]),
        .Q(desOut[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [26]),
        .Q(desOut[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/desOut_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/FP [58]),
        .Q(desOut[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][0]_srl2_n_0 ),
        .Q(\u2/key_r [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][10]_srl2_n_0 ),
        .Q(\u2/key_r [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][11]_srl2_n_0 ),
        .Q(\u2/key_r [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][12]_srl2_n_0 ),
        .Q(\u2/key_r [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][13]_srl2_n_0 ),
        .Q(\u2/key_r [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][14]_srl2_n_0 ),
        .Q(\u2/key_r [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][15]_srl2_n_0 ),
        .Q(\u2/key_r [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][16]_srl2_n_0 ),
        .Q(\u2/key_r [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][17]_srl2_n_0 ),
        .Q(\u2/key_r [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][18]_srl2_n_0 ),
        .Q(\u2/key_r [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][19]_srl2_n_0 ),
        .Q(\u2/key_r [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][1]_srl2_n_0 ),
        .Q(\u2/key_r [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][20]_srl2_n_0 ),
        .Q(\u2/key_r [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][21]_srl2_n_0 ),
        .Q(\u2/key_r [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][22]_srl2_n_0 ),
        .Q(\u2/key_r [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][23]_srl2_n_0 ),
        .Q(\u2/key_r [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][24]_srl2_n_0 ),
        .Q(\u2/key_r [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][25]_srl2_n_0 ),
        .Q(\u2/key_r [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][26]_srl2_n_0 ),
        .Q(\u2/key_r [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][27]_srl2_n_0 ),
        .Q(\u2/key_r [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][28]_srl2_n_0 ),
        .Q(\u2/key_r [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][29]_srl2_n_0 ),
        .Q(\u2/key_r [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][2]_srl2_n_0 ),
        .Q(\u2/key_r [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][30]_srl2_n_0 ),
        .Q(\u2/key_r [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][31]_srl2_n_0 ),
        .Q(\u2/key_r [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][32]_srl2_n_0 ),
        .Q(\u2/key_r [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][33]_srl2_n_0 ),
        .Q(\u2/key_r [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][34]_srl2_n_0 ),
        .Q(\u2/key_r [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][35]_srl2_n_0 ),
        .Q(\u2/key_r [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][36]_srl2_n_0 ),
        .Q(\u2/key_r [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][37]_srl2_n_0 ),
        .Q(\u2/key_r [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][38]_srl2_n_0 ),
        .Q(\u2/key_r [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][39]_srl2_n_0 ),
        .Q(\u2/key_r [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][3]_srl2_n_0 ),
        .Q(\u2/key_r [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][40]_srl2_n_0 ),
        .Q(\u2/key_r [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][41]_srl2_n_0 ),
        .Q(\u2/key_r [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][42]_srl2_n_0 ),
        .Q(\u2/key_r [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][43]_srl2_n_0 ),
        .Q(\u2/key_r [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][44]_srl2_n_0 ),
        .Q(\u2/key_r [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][45]_srl2_n_0 ),
        .Q(\u2/key_r [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][46]_srl2_n_0 ),
        .Q(\u2/key_r [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][47]_srl2_n_0 ),
        .Q(\u2/key_r [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][48]_srl2_n_0 ),
        .Q(\u2/key_r [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][49]_srl2_n_0 ),
        .Q(\u2/key_r [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][4]_srl2_n_0 ),
        .Q(\u2/key_r [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][50]_srl2_n_0 ),
        .Q(\u2/key_r [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][51]_srl2_n_0 ),
        .Q(\u2/key_r [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][52]_srl2_n_0 ),
        .Q(\u2/key_r [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][53]_srl2_n_0 ),
        .Q(\u2/key_r [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][54]_srl2_n_0 ),
        .Q(\u2/key_r [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][55]_srl2_n_0 ),
        .Q(\u2/key_r [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][5]_srl2_n_0 ),
        .Q(\u2/key_r [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][6]_srl2_n_0 ),
        .Q(\u2/key_r [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][7]_srl2_n_0 ),
        .Q(\u2/key_r [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][8]_srl2_n_0 ),
        .Q(\u2/key_r [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/key_r_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\key_c_r_reg[33][9]_srl2_n_0 ),
        .Q(\u2/key_r [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [0]),
        .Q(\u2/uk/K_r0_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [10]),
        .Q(\u2/uk/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [11]),
        .Q(\u2/uk/p_14_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [12]),
        .Q(\u2/uk/p_38_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [13]),
        .Q(\u2/uk/p_7_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [14]),
        .Q(\u2/uk/p_36_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [15]),
        .Q(\u2/uk/p_25_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [16]),
        .Q(\u2/uk/p_27_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [17]),
        .Q(\u2/uk/K_r0_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [18]),
        .Q(\u2/uk/p_37_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [19]),
        .Q(\u2/uk/K_r0_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [1]),
        .Q(\u2/uk/K_r0_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [20]),
        .Q(\u2/uk/p_2_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [21]),
        .Q(\u2/uk/p_24_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [22]),
        .Q(\u2/uk/K_r0_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [23]),
        .Q(\u2/uk/p_30_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [24]),
        .Q(\u2/uk/p_3_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [25]),
        .Q(\u2/uk/K_r0_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [26]),
        .Q(\u2/uk/p_9_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [27]),
        .Q(\u2/uk/p_5_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [28]),
        .Q(\u2/uk/p_20_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [29]),
        .Q(\u2/uk/p_31_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [2]),
        .Q(\u2/uk/K_r0_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [30]),
        .Q(\u2/uk/p_22_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [31]),
        .Q(\u2/uk/K_r0_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [32]),
        .Q(\u2/uk/K_r0_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [33]),
        .Q(\u2/uk/p_39_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [34]),
        .Q(\u2/uk/p_6_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [35]),
        .Q(\u2/uk/K_r0_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [36]),
        .Q(\u2/uk/K_r0_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [37]),
        .Q(\u2/uk/p_26_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [38]),
        .Q(\u2/uk/p_18_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [39]),
        .Q(\u2/uk/p_12_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [3]),
        .Q(\u2/uk/p_11_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [40]),
        .Q(\u2/uk/p_8_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [41]),
        .Q(\u2/uk/p_13_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [42]),
        .Q(\u2/uk/p_29_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [43]),
        .Q(\u2/uk/p_17_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [44]),
        .Q(\u2/uk/p_19_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [45]),
        .Q(\u2/uk/p_33_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [46]),
        .Q(\u2/uk/p_1_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [47]),
        .Q(\u2/uk/p_15_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [48]),
        .Q(\u2/uk/p_4_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [49]),
        .Q(\u2/uk/p_34_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [4]),
        .Q(\u2/uk/K_r0_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [50]),
        .Q(\u2/uk/p_28_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [51]),
        .Q(\u2/uk/p_35_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [52]),
        .Q(\u2/uk/K_r0_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [53]),
        .Q(\u2/uk/K_r0_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [54]),
        .Q(\u2/uk/p_40_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [55]),
        .Q(\u2/uk/K_r0_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [5]),
        .Q(\u2/uk/p_10_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [6]),
        .Q(\u2/uk/p_16_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [7]),
        .Q(\u2/uk/p_21_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [8]),
        .Q(\u2/uk/p_32_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r0_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/key_r [9]),
        .Q(\u2/uk/p_23_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [0]),
        .Q(\u2/uk/K_r10 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [10]),
        .Q(\u2/uk/K_r10 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [11]),
        .Q(\u2/uk/K_r10 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [12]),
        .Q(\u2/uk/K_r10 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [13]),
        .Q(\u2/uk/K_r10 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [14]),
        .Q(\u2/uk/K_r10 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [15]),
        .Q(\u2/uk/K_r10 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [16]),
        .Q(\u2/uk/K_r10 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [17]),
        .Q(\u2/uk/K_r10 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [18]),
        .Q(\u2/uk/K_r10 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [19]),
        .Q(\u2/uk/K_r10 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [1]),
        .Q(\u2/uk/K_r10 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [20]),
        .Q(\u2/uk/K_r10 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [21]),
        .Q(\u2/uk/K_r10 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [22]),
        .Q(\u2/uk/K_r10 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [23]),
        .Q(\u2/uk/K_r10 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [24]),
        .Q(\u2/uk/K_r10 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [25]),
        .Q(\u2/uk/K_r10 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [26]),
        .Q(\u2/uk/K_r10 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [27]),
        .Q(\u2/uk/K_r10 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [28]),
        .Q(\u2/uk/K_r10 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [29]),
        .Q(\u2/uk/K_r10 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [2]),
        .Q(\u2/uk/K_r10 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [30]),
        .Q(\u2/uk/K_r10 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [31]),
        .Q(\u2/uk/K_r10 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [32]),
        .Q(\u2/uk/K_r10 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [33]),
        .Q(\u2/uk/K_r10 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [34]),
        .Q(\u2/uk/K_r10 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [35]),
        .Q(\u2/uk/K_r10 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [36]),
        .Q(\u2/uk/K_r10 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [37]),
        .Q(\u2/uk/K_r10 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [38]),
        .Q(\u2/uk/K_r10 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [39]),
        .Q(\u2/uk/K_r10 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [3]),
        .Q(\u2/uk/K_r10 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [40]),
        .Q(\u2/uk/K_r10 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [41]),
        .Q(\u2/uk/K_r10 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [42]),
        .Q(\u2/uk/K_r10 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [43]),
        .Q(\u2/uk/K_r10 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [44]),
        .Q(\u2/uk/K_r10 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [45]),
        .Q(\u2/uk/K_r10 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [46]),
        .Q(\u2/uk/K_r10 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [47]),
        .Q(\u2/uk/K_r10 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [48]),
        .Q(\u2/uk/K_r10 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [49]),
        .Q(\u2/uk/K_r10 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [4]),
        .Q(\u2/uk/K_r10 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [50]),
        .Q(\u2/uk/K_r10 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [51]),
        .Q(\u2/uk/K_r10 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [52]),
        .Q(\u2/uk/K_r10 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [53]),
        .Q(\u2/uk/K_r10 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [54]),
        .Q(\u2/uk/K_r10 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [55]),
        .Q(\u2/uk/K_r10 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [5]),
        .Q(\u2/uk/K_r10 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [6]),
        .Q(\u2/uk/K_r10 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [7]),
        .Q(\u2/uk/K_r10 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [8]),
        .Q(\u2/uk/K_r10 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r10_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r9 [9]),
        .Q(\u2/uk/K_r10 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [0]),
        .Q(\u2/uk/K_r11 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [10]),
        .Q(\u2/uk/K_r11 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [11]),
        .Q(\u2/uk/K_r11 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [12]),
        .Q(\u2/uk/K_r11 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [13]),
        .Q(\u2/uk/K_r11 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [14]),
        .Q(\u2/uk/K_r11 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [15]),
        .Q(\u2/uk/K_r11 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [16]),
        .Q(\u2/uk/K_r11 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [17]),
        .Q(\u2/uk/K_r11 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [18]),
        .Q(\u2/uk/K_r11 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [19]),
        .Q(\u2/uk/K_r11 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [1]),
        .Q(\u2/uk/K_r11 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [20]),
        .Q(\u2/uk/K_r11 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [21]),
        .Q(\u2/uk/K_r11 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [22]),
        .Q(\u2/uk/K_r11 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [23]),
        .Q(\u2/uk/K_r11 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [24]),
        .Q(\u2/uk/K_r11 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [25]),
        .Q(\u2/uk/K_r11 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [26]),
        .Q(\u2/uk/K_r11 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [27]),
        .Q(\u2/uk/K_r11 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [28]),
        .Q(\u2/uk/K_r11 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [29]),
        .Q(\u2/uk/K_r11 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [2]),
        .Q(\u2/uk/K_r11 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [30]),
        .Q(\u2/uk/K_r11 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [31]),
        .Q(\u2/uk/K_r11 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [32]),
        .Q(\u2/uk/K_r11 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [33]),
        .Q(\u2/uk/K_r11 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [34]),
        .Q(\u2/uk/K_r11 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [35]),
        .Q(\u2/uk/K_r11 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [36]),
        .Q(\u2/uk/K_r11 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [37]),
        .Q(\u2/uk/K_r11 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [38]),
        .Q(\u2/uk/K_r11 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [39]),
        .Q(\u2/uk/K_r11 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [3]),
        .Q(\u2/uk/K_r11 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [40]),
        .Q(\u2/uk/K_r11 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [41]),
        .Q(\u2/uk/K_r11 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [42]),
        .Q(\u2/uk/K_r11 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [43]),
        .Q(\u2/uk/K_r11 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [44]),
        .Q(\u2/uk/K_r11 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [45]),
        .Q(\u2/uk/K_r11 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [46]),
        .Q(\u2/uk/K_r11 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [47]),
        .Q(\u2/uk/K_r11 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [48]),
        .Q(\u2/uk/K_r11 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [49]),
        .Q(\u2/uk/K_r11 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [4]),
        .Q(\u2/uk/K_r11 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [50]),
        .Q(\u2/uk/K_r11 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [51]),
        .Q(\u2/uk/K_r11 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [52]),
        .Q(\u2/uk/K_r11 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [53]),
        .Q(\u2/uk/K_r11 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [54]),
        .Q(\u2/uk/K_r11 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [55]),
        .Q(\u2/uk/K_r11 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [5]),
        .Q(\u2/uk/K_r11 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [6]),
        .Q(\u2/uk/K_r11 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [7]),
        .Q(\u2/uk/K_r11 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [8]),
        .Q(\u2/uk/K_r11 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r11_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r10 [9]),
        .Q(\u2/uk/K_r11 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [0]),
        .Q(\u2/uk/K_r12 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [10]),
        .Q(\u2/uk/K_r12 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [11]),
        .Q(\u2/uk/K_r12 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [12]),
        .Q(\u2/uk/K_r12 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [13]),
        .Q(\u2/uk/K_r12 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [14]),
        .Q(\u2/uk/K_r12 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [15]),
        .Q(\u2/uk/K_r12 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [16]),
        .Q(\u2/uk/K_r12 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [17]),
        .Q(\u2/uk/K_r12 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [18]),
        .Q(\u2/uk/K_r12 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [19]),
        .Q(\u2/uk/K_r12 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [1]),
        .Q(\u2/uk/K_r12 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [20]),
        .Q(\u2/uk/K_r12 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [21]),
        .Q(\u2/uk/K_r12 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [22]),
        .Q(\u2/uk/K_r12 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [23]),
        .Q(\u2/uk/K_r12 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [24]),
        .Q(\u2/uk/K_r12 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [25]),
        .Q(\u2/uk/K_r12 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [26]),
        .Q(\u2/uk/K_r12 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [27]),
        .Q(\u2/uk/K_r12 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [28]),
        .Q(\u2/uk/K_r12 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [29]),
        .Q(\u2/uk/K_r12 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [2]),
        .Q(\u2/uk/K_r12 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [30]),
        .Q(\u2/uk/K_r12 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [31]),
        .Q(\u2/uk/K_r12 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [32]),
        .Q(\u2/uk/K_r12 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [33]),
        .Q(\u2/uk/K_r12 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [34]),
        .Q(\u2/uk/K_r12 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [35]),
        .Q(\u2/uk/K_r12 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [36]),
        .Q(\u2/uk/K_r12 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [37]),
        .Q(\u2/uk/K_r12 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [38]),
        .Q(\u2/uk/K_r12 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [39]),
        .Q(\u2/uk/K_r12 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [3]),
        .Q(\u2/uk/K_r12 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [40]),
        .Q(\u2/uk/K_r12 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [41]),
        .Q(\u2/uk/K_r12 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [42]),
        .Q(\u2/uk/K_r12 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [43]),
        .Q(\u2/uk/K_r12 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [44]),
        .Q(\u2/uk/K_r12 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [45]),
        .Q(\u2/uk/K_r12 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [46]),
        .Q(\u2/uk/K_r12 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [47]),
        .Q(\u2/uk/K_r12 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [48]),
        .Q(\u2/uk/K_r12 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [49]),
        .Q(\u2/uk/K_r12 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [4]),
        .Q(\u2/uk/K_r12 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [50]),
        .Q(\u2/uk/K_r12 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [51]),
        .Q(\u2/uk/K_r12 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [52]),
        .Q(\u2/uk/K_r12 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [53]),
        .Q(\u2/uk/K_r12 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [54]),
        .Q(\u2/uk/K_r12 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [55]),
        .Q(\u2/uk/K_r12 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [5]),
        .Q(\u2/uk/K_r12 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [6]),
        .Q(\u2/uk/K_r12 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [7]),
        .Q(\u2/uk/K_r12 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [8]),
        .Q(\u2/uk/K_r12 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r12_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r11 [9]),
        .Q(\u2/uk/K_r12 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [0]),
        .Q(\u2/uk/K_r13 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [10]),
        .Q(\u2/uk/K_r13 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [11]),
        .Q(\u2/uk/K_r13 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [12]),
        .Q(\u2/uk/K_r13 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [13]),
        .Q(\u2/uk/K_r13 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [14]),
        .Q(\u2/uk/K_r13 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [15]),
        .Q(\u2/uk/K_r13 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [16]),
        .Q(\u2/uk/K_r13 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [17]),
        .Q(\u2/uk/K_r13 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [18]),
        .Q(\u2/uk/K_r13 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [19]),
        .Q(\u2/uk/K_r13 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [1]),
        .Q(\u2/uk/K_r13 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [20]),
        .Q(\u2/uk/K_r13 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [21]),
        .Q(\u2/uk/K_r13 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [22]),
        .Q(\u2/uk/K_r13 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [23]),
        .Q(\u2/uk/K_r13 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [24]),
        .Q(\u2/uk/K_r13 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [25]),
        .Q(\u2/uk/K_r13 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [26]),
        .Q(\u2/uk/K_r13 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [27]),
        .Q(\u2/uk/K_r13 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [28]),
        .Q(\u2/uk/K_r13 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [29]),
        .Q(\u2/uk/K_r13 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [2]),
        .Q(\u2/uk/K_r13 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [30]),
        .Q(\u2/uk/K_r13 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [31]),
        .Q(\u2/uk/K_r13 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [32]),
        .Q(\u2/uk/K_r13 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [33]),
        .Q(\u2/uk/K_r13 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [34]),
        .Q(\u2/uk/K_r13 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [35]),
        .Q(\u2/uk/K_r13 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [36]),
        .Q(\u2/uk/K_r13 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [37]),
        .Q(\u2/uk/K_r13 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [38]),
        .Q(\u2/uk/K_r13 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [39]),
        .Q(\u2/uk/K_r13 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [3]),
        .Q(\u2/uk/K_r13 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [40]),
        .Q(\u2/uk/K_r13 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [41]),
        .Q(\u2/uk/K_r13 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [42]),
        .Q(\u2/uk/K_r13 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [43]),
        .Q(\u2/uk/K_r13 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [44]),
        .Q(\u2/uk/K_r13 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [45]),
        .Q(\u2/uk/K_r13 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [46]),
        .Q(\u2/uk/K_r13 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [47]),
        .Q(\u2/uk/K_r13 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [48]),
        .Q(\u2/uk/K_r13 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [49]),
        .Q(\u2/uk/K_r13 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [4]),
        .Q(\u2/uk/K_r13 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [50]),
        .Q(\u2/uk/K_r13 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [51]),
        .Q(\u2/uk/K_r13 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [52]),
        .Q(\u2/uk/K_r13 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [53]),
        .Q(\u2/uk/K_r13 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [54]),
        .Q(\u2/uk/K_r13 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [55]),
        .Q(\u2/uk/K_r13 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [5]),
        .Q(\u2/uk/K_r13 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [6]),
        .Q(\u2/uk/K_r13 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [7]),
        .Q(\u2/uk/K_r13 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [8]),
        .Q(\u2/uk/K_r13 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r13_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r12 [9]),
        .Q(\u2/uk/K_r13 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [0]),
        .Q(\u2/uk/K_r14_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [10]),
        .Q(\u2/uk/K_r14_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [11]),
        .Q(\u2/uk/K_r14_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [12]),
        .Q(\u2/uk/K_r14_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [13]),
        .Q(\u2/uk/K_r14_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [14]),
        .Q(\u2/uk/K_r14_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [15]),
        .Q(\u2/uk/K_r14_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [16]),
        .Q(\u2/uk/K_r14_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [17]),
        .Q(\u2/uk/K_r14_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [18]),
        .Q(\u2/uk/K_r14_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [19]),
        .Q(\u2/uk/K_r14_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [1]),
        .Q(\u2/uk/K_r14_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [20]),
        .Q(\u2/uk/K_r14_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [21]),
        .Q(\u2/uk/K_r14_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [22]),
        .Q(\u2/uk/K_r14_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [23]),
        .Q(\u2/uk/K_r14_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [24]),
        .Q(\u2/uk/K_r14_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [25]),
        .Q(\u2/uk/K_r14_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [26]),
        .Q(\u2/uk/K_r14_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [27]),
        .Q(\u2/uk/K_r14_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [28]),
        .Q(\u2/uk/K_r14_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [29]),
        .Q(\u2/uk/K_r14_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [2]),
        .Q(\u2/uk/K_r14_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [30]),
        .Q(\u2/uk/K_r14_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [31]),
        .Q(\u2/uk/K_r14_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [32]),
        .Q(\u2/uk/K_r14_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [33]),
        .Q(\u2/uk/K_r14_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [34]),
        .Q(\u2/uk/K_r14_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [35]),
        .Q(\u2/uk/K_r14_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [36]),
        .Q(\u2/uk/K_r14_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [37]),
        .Q(\u2/uk/K_r14_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [38]),
        .Q(\u2/uk/K_r14_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [39]),
        .Q(\u2/uk/K_r14_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [3]),
        .Q(\u2/uk/K_r14_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [40]),
        .Q(\u2/uk/K_r14_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [41]),
        .Q(\u2/uk/K_r14_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [42]),
        .Q(\u2/uk/K_r14_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [43]),
        .Q(\u2/uk/K_r14_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [44]),
        .Q(\u2/uk/K_r14_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [45]),
        .Q(\u2/uk/K_r14_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [46]),
        .Q(\u2/uk/K_r14_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [47]),
        .Q(\u2/uk/K_r14_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [48]),
        .Q(\u2/uk/K_r14_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [49]),
        .Q(\u2/uk/K_r14_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [4]),
        .Q(\u2/uk/K_r14_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [50]),
        .Q(\u2/uk/K_r14_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [51]),
        .Q(\u2/uk/K_r14_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [52]),
        .Q(\u2/uk/K_r14_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [53]),
        .Q(\u2/uk/K_r14_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [54]),
        .Q(\u2/uk/K_r14_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [55]),
        .Q(\u2/uk/K_r14_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [5]),
        .Q(\u2/uk/K_r14_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [6]),
        .Q(\u2/uk/K_r14_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [7]),
        .Q(\u2/uk/K_r14_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [8]),
        .Q(\u2/uk/K_r14_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r14_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r13 [9]),
        .Q(\u2/uk/K_r14_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_ ),
        .Q(\u2/uk/K_r1 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_0_in ),
        .Q(\u2/uk/K_r1 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_14_in ),
        .Q(\u2/uk/K_r1 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_38_in ),
        .Q(\u2/uk/K_r1 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_7_in ),
        .Q(\u2/uk/K_r1 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_36_in ),
        .Q(\u2/uk/K_r1 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_25_in ),
        .Q(\u2/uk/K_r1 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_27_in ),
        .Q(\u2/uk/K_r1 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[17] ),
        .Q(\u2/uk/K_r1 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_37_in ),
        .Q(\u2/uk/K_r1 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[19] ),
        .Q(\u2/uk/K_r1 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[1] ),
        .Q(\u2/uk/K_r1 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_2_in ),
        .Q(\u2/uk/K_r1 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_24_in ),
        .Q(\u2/uk/K_r1 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[22] ),
        .Q(\u2/uk/K_r1 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_30_in ),
        .Q(\u2/uk/K_r1 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_3_in ),
        .Q(\u2/uk/K_r1 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[25] ),
        .Q(\u2/uk/K_r1 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_9_in ),
        .Q(\u2/uk/K_r1 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_5_in ),
        .Q(\u2/uk/K_r1 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_20_in ),
        .Q(\u2/uk/K_r1 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_31_in ),
        .Q(\u2/uk/K_r1 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[2] ),
        .Q(\u2/uk/K_r1 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_22_in ),
        .Q(\u2/uk/K_r1 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[31] ),
        .Q(\u2/uk/K_r1 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[32] ),
        .Q(\u2/uk/K_r1 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_39_in ),
        .Q(\u2/uk/K_r1 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_6_in ),
        .Q(\u2/uk/K_r1 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[35] ),
        .Q(\u2/uk/K_r1 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[36] ),
        .Q(\u2/uk/K_r1 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_26_in ),
        .Q(\u2/uk/K_r1 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_18_in ),
        .Q(\u2/uk/K_r1 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_12_in ),
        .Q(\u2/uk/K_r1 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_11_in ),
        .Q(\u2/uk/K_r1 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_8_in ),
        .Q(\u2/uk/K_r1 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_13_in ),
        .Q(\u2/uk/K_r1 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_29_in ),
        .Q(\u2/uk/K_r1 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_17_in ),
        .Q(\u2/uk/K_r1 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_19_in ),
        .Q(\u2/uk/K_r1 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_33_in ),
        .Q(\u2/uk/K_r1 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_1_in ),
        .Q(\u2/uk/K_r1 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_15_in ),
        .Q(\u2/uk/K_r1 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_4_in ),
        .Q(\u2/uk/K_r1 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_34_in ),
        .Q(\u2/uk/K_r1 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[4] ),
        .Q(\u2/uk/K_r1 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_28_in ),
        .Q(\u2/uk/K_r1 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_35_in ),
        .Q(\u2/uk/K_r1 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[52] ),
        .Q(\u2/uk/K_r1 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[53] ),
        .Q(\u2/uk/K_r1 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_40_in ),
        .Q(\u2/uk/K_r1 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r0_reg_n_0_[55] ),
        .Q(\u2/uk/K_r1 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_10_in ),
        .Q(\u2/uk/K_r1 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_16_in ),
        .Q(\u2/uk/K_r1 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_21_in ),
        .Q(\u2/uk/K_r1 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_32_in ),
        .Q(\u2/uk/K_r1 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r1_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_23_in ),
        .Q(\u2/uk/K_r1 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [0]),
        .Q(\u2/uk/K_r2 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [10]),
        .Q(\u2/uk/K_r2 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [11]),
        .Q(\u2/uk/K_r2 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [12]),
        .Q(\u2/uk/K_r2 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [13]),
        .Q(\u2/uk/K_r2 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [14]),
        .Q(\u2/uk/K_r2 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [15]),
        .Q(\u2/uk/K_r2 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [16]),
        .Q(\u2/uk/K_r2 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [17]),
        .Q(\u2/uk/K_r2 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [18]),
        .Q(\u2/uk/K_r2 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [19]),
        .Q(\u2/uk/K_r2 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [1]),
        .Q(\u2/uk/K_r2 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [20]),
        .Q(\u2/uk/K_r2 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [21]),
        .Q(\u2/uk/K_r2 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [22]),
        .Q(\u2/uk/K_r2 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [23]),
        .Q(\u2/uk/K_r2 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [24]),
        .Q(\u2/uk/K_r2 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [25]),
        .Q(\u2/uk/K_r2 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [26]),
        .Q(\u2/uk/K_r2 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [27]),
        .Q(\u2/uk/K_r2 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [28]),
        .Q(\u2/uk/K_r2 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [29]),
        .Q(\u2/uk/K_r2 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [2]),
        .Q(\u2/uk/K_r2 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [30]),
        .Q(\u2/uk/K_r2 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [31]),
        .Q(\u2/uk/K_r2 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [32]),
        .Q(\u2/uk/K_r2 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [33]),
        .Q(\u2/uk/K_r2 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [34]),
        .Q(\u2/uk/K_r2 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [35]),
        .Q(\u2/uk/K_r2 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [36]),
        .Q(\u2/uk/K_r2 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [37]),
        .Q(\u2/uk/K_r2 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [38]),
        .Q(\u2/uk/K_r2 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [39]),
        .Q(\u2/uk/K_r2 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [3]),
        .Q(\u2/uk/K_r2 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [40]),
        .Q(\u2/uk/K_r2 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [41]),
        .Q(\u2/uk/K_r2 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [42]),
        .Q(\u2/uk/K_r2 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [43]),
        .Q(\u2/uk/K_r2 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [44]),
        .Q(\u2/uk/K_r2 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [45]),
        .Q(\u2/uk/K_r2 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [46]),
        .Q(\u2/uk/K_r2 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [47]),
        .Q(\u2/uk/K_r2 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [48]),
        .Q(\u2/uk/K_r2 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [49]),
        .Q(\u2/uk/K_r2 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [4]),
        .Q(\u2/uk/K_r2 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [50]),
        .Q(\u2/uk/K_r2 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [51]),
        .Q(\u2/uk/K_r2 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [52]),
        .Q(\u2/uk/K_r2 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [53]),
        .Q(\u2/uk/K_r2 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [54]),
        .Q(\u2/uk/K_r2 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [55]),
        .Q(\u2/uk/K_r2 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [5]),
        .Q(\u2/uk/K_r2 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [6]),
        .Q(\u2/uk/K_r2 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [7]),
        .Q(\u2/uk/K_r2 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [8]),
        .Q(\u2/uk/K_r2 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r2_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r1 [9]),
        .Q(\u2/uk/K_r2 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [0]),
        .Q(\u2/uk/K_r3 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [10]),
        .Q(\u2/uk/K_r3 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [11]),
        .Q(\u2/uk/K_r3 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [12]),
        .Q(\u2/uk/K_r3 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [13]),
        .Q(\u2/uk/K_r3 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [14]),
        .Q(\u2/uk/K_r3 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [15]),
        .Q(\u2/uk/K_r3 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [16]),
        .Q(\u2/uk/K_r3 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [17]),
        .Q(\u2/uk/K_r3 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [18]),
        .Q(\u2/uk/K_r3 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [19]),
        .Q(\u2/uk/K_r3 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [1]),
        .Q(\u2/uk/K_r3 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [20]),
        .Q(\u2/uk/K_r3 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [21]),
        .Q(\u2/uk/K_r3 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [22]),
        .Q(\u2/uk/K_r3 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [23]),
        .Q(\u2/uk/K_r3 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [24]),
        .Q(\u2/uk/K_r3 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [25]),
        .Q(\u2/uk/K_r3 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [26]),
        .Q(\u2/uk/K_r3 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [27]),
        .Q(\u2/uk/K_r3 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [28]),
        .Q(\u2/uk/K_r3 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [29]),
        .Q(\u2/uk/K_r3 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [2]),
        .Q(\u2/uk/K_r3 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [30]),
        .Q(\u2/uk/K_r3 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [31]),
        .Q(\u2/uk/K_r3 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [32]),
        .Q(\u2/uk/K_r3 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [33]),
        .Q(\u2/uk/K_r3 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [34]),
        .Q(\u2/uk/K_r3 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [35]),
        .Q(\u2/uk/K_r3 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [36]),
        .Q(\u2/uk/K_r3 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [37]),
        .Q(\u2/uk/K_r3 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [38]),
        .Q(\u2/uk/K_r3 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [39]),
        .Q(\u2/uk/K_r3 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [3]),
        .Q(\u2/uk/K_r3 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [40]),
        .Q(\u2/uk/K_r3 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [41]),
        .Q(\u2/uk/K_r3 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [42]),
        .Q(\u2/uk/K_r3 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [43]),
        .Q(\u2/uk/K_r3 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [44]),
        .Q(\u2/uk/K_r3 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [45]),
        .Q(\u2/uk/K_r3 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [46]),
        .Q(\u2/uk/K_r3 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [47]),
        .Q(\u2/uk/K_r3 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [48]),
        .Q(\u2/uk/K_r3 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [49]),
        .Q(\u2/uk/K_r3 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [4]),
        .Q(\u2/uk/K_r3 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [50]),
        .Q(\u2/uk/K_r3 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [51]),
        .Q(\u2/uk/K_r3 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [52]),
        .Q(\u2/uk/K_r3 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [53]),
        .Q(\u2/uk/K_r3 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [54]),
        .Q(\u2/uk/K_r3 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [55]),
        .Q(\u2/uk/K_r3 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [5]),
        .Q(\u2/uk/K_r3 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [6]),
        .Q(\u2/uk/K_r3 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [7]),
        .Q(\u2/uk/K_r3 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [8]),
        .Q(\u2/uk/K_r3 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r3_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r2 [9]),
        .Q(\u2/uk/K_r3 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [0]),
        .Q(\u2/uk/K_r4_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [10]),
        .Q(\u2/uk/K_r4_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [11]),
        .Q(\u2/uk/K_r4_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [12]),
        .Q(\u2/uk/K_r4_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [13]),
        .Q(\u2/uk/K_r4_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [14]),
        .Q(\u2/uk/K_r4_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [15]),
        .Q(\u2/uk/K_r4_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [16]),
        .Q(\u2/uk/K_r4_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [17]),
        .Q(\u2/uk/K_r4_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [18]),
        .Q(\u2/uk/K_r4_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [19]),
        .Q(\u2/uk/K_r4_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [1]),
        .Q(\u2/uk/K_r4_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [20]),
        .Q(\u2/uk/K_r4_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [21]),
        .Q(\u2/uk/K_r4_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [22]),
        .Q(\u2/uk/K_r4_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [23]),
        .Q(\u2/uk/K_r4_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [24]),
        .Q(\u2/uk/K_r4_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [25]),
        .Q(\u2/uk/K_r4_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [26]),
        .Q(\u2/uk/K_r4_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [27]),
        .Q(\u2/uk/K_r4_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [28]),
        .Q(\u2/uk/K_r4_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [29]),
        .Q(\u2/uk/K_r4_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [2]),
        .Q(\u2/uk/K_r4_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [30]),
        .Q(\u2/uk/K_r4_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [31]),
        .Q(\u2/uk/K_r4_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [32]),
        .Q(\u2/uk/K_r4_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [33]),
        .Q(\u2/uk/K_r4_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [34]),
        .Q(\u2/uk/p_50_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [35]),
        .Q(\u2/uk/K_r4_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [36]),
        .Q(\u2/uk/K_r4_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [37]),
        .Q(\u2/uk/K_r4_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [38]),
        .Q(\u2/uk/K_r4_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [39]),
        .Q(\u2/uk/K_r4_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [3]),
        .Q(\u2/uk/K_r4_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [40]),
        .Q(\u2/uk/p_49_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [41]),
        .Q(\u2/uk/K_r4_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [42]),
        .Q(\u2/uk/K_r4_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [43]),
        .Q(\u2/uk/p_44_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [44]),
        .Q(\u2/uk/K_r4_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [45]),
        .Q(\u2/uk/K_r4_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [46]),
        .Q(\u2/uk/p_47_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [47]),
        .Q(\u2/uk/K_r4_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [48]),
        .Q(\u2/uk/K_r4_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [49]),
        .Q(\u2/uk/K_r4_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [4]),
        .Q(\u2/uk/K_r4_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [50]),
        .Q(\u2/uk/K_r4_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [51]),
        .Q(\u2/uk/K_r4_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [52]),
        .Q(\u2/uk/K_r4_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [53]),
        .Q(\u2/uk/p_51_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [54]),
        .Q(\u2/uk/K_r4_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [55]),
        .Q(\u2/uk/K_r4_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [5]),
        .Q(\u2/uk/K_r4_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [6]),
        .Q(\u2/uk/K_r4_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [7]),
        .Q(\u2/uk/K_r4_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [8]),
        .Q(\u2/uk/p_42_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r4_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r3 [9]),
        .Q(\u2/uk/K_r4_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_ ),
        .Q(\u2/uk/K_r5 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[10] ),
        .Q(\u2/uk/K_r5 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[11] ),
        .Q(\u2/uk/K_r5 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[12] ),
        .Q(\u2/uk/K_r5 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[13] ),
        .Q(\u2/uk/K_r5 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[14] ),
        .Q(\u2/uk/K_r5 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[15] ),
        .Q(\u2/uk/K_r5 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[16] ),
        .Q(\u2/uk/K_r5 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[17] ),
        .Q(\u2/uk/K_r5 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[18] ),
        .Q(\u2/uk/K_r5 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[19] ),
        .Q(\u2/uk/K_r5 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[1] ),
        .Q(\u2/uk/K_r5 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[20] ),
        .Q(\u2/uk/K_r5 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[21] ),
        .Q(\u2/uk/K_r5 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[22] ),
        .Q(\u2/uk/K_r5 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[23] ),
        .Q(\u2/uk/K_r5 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[24] ),
        .Q(\u2/uk/K_r5 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[25] ),
        .Q(\u2/uk/K_r5 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[26] ),
        .Q(\u2/uk/K_r5 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[27] ),
        .Q(\u2/uk/K_r5 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[28] ),
        .Q(\u2/uk/K_r5 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[29] ),
        .Q(\u2/uk/K_r5 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[2] ),
        .Q(\u2/uk/K_r5 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[30] ),
        .Q(\u2/uk/K_r5 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[31] ),
        .Q(\u2/uk/K_r5 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[32] ),
        .Q(\u2/uk/K_r5 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[33] ),
        .Q(\u2/uk/K_r5 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_50_in ),
        .Q(\u2/uk/K_r5 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[35] ),
        .Q(\u2/uk/K_r5 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[36] ),
        .Q(\u2/uk/K_r5 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[37] ),
        .Q(\u2/uk/K_r5 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[38] ),
        .Q(\u2/uk/K_r5 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[39] ),
        .Q(\u2/uk/K_r5 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[3] ),
        .Q(\u2/uk/K_r5 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_49_in ),
        .Q(\u2/uk/K_r5 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[41] ),
        .Q(\u2/uk/K_r5 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[42] ),
        .Q(\u2/uk/K_r5 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_44_in ),
        .Q(\u2/uk/K_r5 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[44] ),
        .Q(\u2/uk/K_r5 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[45] ),
        .Q(\u2/uk/K_r5 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_47_in ),
        .Q(\u2/uk/K_r5 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[47] ),
        .Q(\u2/uk/K_r5 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[48] ),
        .Q(\u2/uk/K_r5 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[49] ),
        .Q(\u2/uk/K_r5 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[4] ),
        .Q(\u2/uk/K_r5 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[50] ),
        .Q(\u2/uk/K_r5 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[51] ),
        .Q(\u2/uk/K_r5 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[52] ),
        .Q(\u2/uk/K_r5 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_51_in ),
        .Q(\u2/uk/K_r5 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[54] ),
        .Q(\u2/uk/K_r5 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[55] ),
        .Q(\u2/uk/K_r5 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[5] ),
        .Q(\u2/uk/K_r5 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[6] ),
        .Q(\u2/uk/K_r5 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[7] ),
        .Q(\u2/uk/K_r5 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_42_in ),
        .Q(\u2/uk/K_r5 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r5_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r4_reg_n_0_[9] ),
        .Q(\u2/uk/K_r5 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [0]),
        .Q(\u2/uk/K_r6_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [10]),
        .Q(\u2/uk/K_r6_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [11]),
        .Q(\u2/uk/K_r6_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [12]),
        .Q(\u2/uk/K_r6_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [13]),
        .Q(\u2/uk/p_52_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [14]),
        .Q(\u2/uk/K_r6_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [15]),
        .Q(\u2/uk/K_r6_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [16]),
        .Q(\u2/uk/K_r6_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [17]),
        .Q(\u2/uk/K_r6_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [18]),
        .Q(\u2/uk/K_r6_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [19]),
        .Q(\u2/uk/K_r6_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [1]),
        .Q(\u2/uk/K_r6_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [20]),
        .Q(\u2/uk/K_r6_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [21]),
        .Q(\u2/uk/K_r6_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [22]),
        .Q(\u2/uk/K_r6_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [23]),
        .Q(\u2/uk/K_r6_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [24]),
        .Q(\u2/uk/K_r6_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [25]),
        .Q(\u2/uk/K_r6_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [26]),
        .Q(\u2/uk/K_r6_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [27]),
        .Q(\u2/uk/K_r6_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [28]),
        .Q(\u2/uk/K_r6_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [29]),
        .Q(\u2/uk/K_r6_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [2]),
        .Q(\u2/uk/K_r6_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [30]),
        .Q(\u2/uk/K_r6_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [31]),
        .Q(\u2/uk/K_r6_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [32]),
        .Q(\u2/uk/K_r6_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [33]),
        .Q(\u2/uk/K_r6_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [34]),
        .Q(\u2/uk/K_r6_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [35]),
        .Q(\u2/uk/K_r6_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [36]),
        .Q(\u2/uk/K_r6_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [37]),
        .Q(\u2/uk/K_r6_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [38]),
        .Q(\u2/uk/K_r6_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [39]),
        .Q(\u2/uk/K_r6_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [3]),
        .Q(\u2/uk/K_r6_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [40]),
        .Q(\u2/uk/K_r6_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [41]),
        .Q(\u2/uk/K_r6_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [42]),
        .Q(\u2/uk/p_41_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [43]),
        .Q(\u2/uk/p_45_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [44]),
        .Q(\u2/uk/K_r6_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [45]),
        .Q(\u2/uk/K_r6_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [46]),
        .Q(\u2/uk/K_r6_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [47]),
        .Q(\u2/uk/K_r6_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [48]),
        .Q(\u2/uk/K_r6_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [49]),
        .Q(\u2/uk/p_43_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [4]),
        .Q(\u2/uk/K_r6_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [50]),
        .Q(\u2/uk/K_r6_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [51]),
        .Q(\u2/uk/K_r6_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [52]),
        .Q(\u2/uk/K_r6_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [53]),
        .Q(\u2/uk/K_r6_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [54]),
        .Q(\u2/uk/K_r6_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [55]),
        .Q(\u2/uk/K_r6_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [5]),
        .Q(\u2/uk/K_r6_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [6]),
        .Q(\u2/uk/p_53_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [7]),
        .Q(\u2/uk/K_r6_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [8]),
        .Q(\u2/uk/K_r6_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r6_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r5 [9]),
        .Q(\u2/uk/K_r6_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_ ),
        .Q(\u2/uk/K_r7_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[10] ),
        .Q(\u2/uk/K_r7_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[11] ),
        .Q(\u2/uk/K_r7_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[12] ),
        .Q(\u2/uk/K_r7_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_52_in ),
        .Q(\u2/uk/K_r7_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[14] ),
        .Q(\u2/uk/K_r7_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[15] ),
        .Q(\u2/uk/K_r7_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[16] ),
        .Q(\u2/uk/K_r7_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[17] ),
        .Q(\u2/uk/K_r7_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[18] ),
        .Q(\u2/uk/K_r7_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[19] ),
        .Q(\u2/uk/K_r7_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[1] ),
        .Q(\u2/uk/K_r7_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[20] ),
        .Q(\u2/uk/K_r7_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[21] ),
        .Q(\u2/uk/K_r7_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[22] ),
        .Q(\u2/uk/K_r7_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[23] ),
        .Q(\u2/uk/K_r7_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[24] ),
        .Q(\u2/uk/K_r7_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[25] ),
        .Q(\u2/uk/K_r7_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[26] ),
        .Q(\u2/uk/K_r7_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[27] ),
        .Q(\u2/uk/K_r7_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[28] ),
        .Q(\u2/uk/K_r7_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[29] ),
        .Q(\u2/uk/K_r7_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[2] ),
        .Q(\u2/uk/K_r7_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[30] ),
        .Q(\u2/uk/K_r7_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[31] ),
        .Q(\u2/uk/K_r7_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[32] ),
        .Q(\u2/uk/K_r7_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[33] ),
        .Q(\u2/uk/K_r7_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[34] ),
        .Q(\u2/uk/K_r7_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[35] ),
        .Q(\u2/uk/K_r7_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[36] ),
        .Q(\u2/uk/K_r7_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[37] ),
        .Q(\u2/uk/K_r7_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[38] ),
        .Q(\u2/uk/K_r7_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[39] ),
        .Q(\u2/uk/K_r7_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[3] ),
        .Q(\u2/uk/K_r7_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[40] ),
        .Q(\u2/uk/K_r7_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[41] ),
        .Q(\u2/uk/K_r7_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_41_in ),
        .Q(\u2/uk/K_r7_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_45_in ),
        .Q(\u2/uk/K_r7_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[44] ),
        .Q(\u2/uk/p_48_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[45] ),
        .Q(\u2/uk/K_r7_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[46] ),
        .Q(\u2/uk/K_r7_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[47] ),
        .Q(\u2/uk/K_r7_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[48] ),
        .Q(\u2/uk/K_r7_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_43_in ),
        .Q(\u2/uk/K_r7_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[4] ),
        .Q(\u2/uk/K_r7_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[50] ),
        .Q(\u2/uk/K_r7_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[51] ),
        .Q(\u2/uk/K_r7_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[52] ),
        .Q(\u2/uk/K_r7_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[53] ),
        .Q(\u2/uk/K_r7_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[54] ),
        .Q(\u2/uk/K_r7_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[55] ),
        .Q(\u2/uk/K_r7_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[5] ),
        .Q(\u2/uk/K_r7_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_53_in ),
        .Q(\u2/uk/K_r7_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[7] ),
        .Q(\u2/uk/K_r7_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[8] ),
        .Q(\u2/uk/K_r7_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r7_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r6_reg_n_0_[9] ),
        .Q(\u2/uk/K_r7_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_ ),
        .Q(\u2/uk/K_r8 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[10] ),
        .Q(\u2/uk/K_r8 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[11] ),
        .Q(\u2/uk/K_r8 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[12] ),
        .Q(\u2/uk/K_r8 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[13] ),
        .Q(\u2/uk/K_r8 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[14] ),
        .Q(\u2/uk/K_r8 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[15] ),
        .Q(\u2/uk/K_r8 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[16] ),
        .Q(\u2/uk/K_r8 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[17] ),
        .Q(\u2/uk/K_r8 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[18] ),
        .Q(\u2/uk/K_r8 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[19] ),
        .Q(\u2/uk/K_r8 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[1] ),
        .Q(\u2/uk/K_r8 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[20] ),
        .Q(\u2/uk/K_r8 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[21] ),
        .Q(\u2/uk/K_r8 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[22] ),
        .Q(\u2/uk/K_r8 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[23] ),
        .Q(\u2/uk/K_r8 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[24] ),
        .Q(\u2/uk/K_r8 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[25] ),
        .Q(\u2/uk/K_r8 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[26] ),
        .Q(\u2/uk/K_r8 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[27] ),
        .Q(\u2/uk/K_r8 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[28] ),
        .Q(\u2/uk/K_r8 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[29] ),
        .Q(\u2/uk/K_r8 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[2] ),
        .Q(\u2/uk/K_r8 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[30] ),
        .Q(\u2/uk/K_r8 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[31] ),
        .Q(\u2/uk/K_r8 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[32] ),
        .Q(\u2/uk/K_r8 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[33] ),
        .Q(\u2/uk/K_r8 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[34] ),
        .Q(\u2/uk/K_r8 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[35] ),
        .Q(\u2/uk/K_r8 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[36] ),
        .Q(\u2/uk/K_r8 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[37] ),
        .Q(\u2/uk/K_r8 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[38] ),
        .Q(\u2/uk/K_r8 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[39] ),
        .Q(\u2/uk/K_r8 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[3] ),
        .Q(\u2/uk/K_r8 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[40] ),
        .Q(\u2/uk/K_r8 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[41] ),
        .Q(\u2/uk/K_r8 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[42] ),
        .Q(\u2/uk/K_r8 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[43] ),
        .Q(\u2/uk/K_r8 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/p_48_in ),
        .Q(\u2/uk/K_r8 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[45] ),
        .Q(\u2/uk/K_r8 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[46] ),
        .Q(\u2/uk/K_r8 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[47] ),
        .Q(\u2/uk/K_r8 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[48] ),
        .Q(\u2/uk/K_r8 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[49] ),
        .Q(\u2/uk/K_r8 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[4] ),
        .Q(\u2/uk/K_r8 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[50] ),
        .Q(\u2/uk/K_r8 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[51] ),
        .Q(\u2/uk/K_r8 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[52] ),
        .Q(\u2/uk/K_r8 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[53] ),
        .Q(\u2/uk/K_r8 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[54] ),
        .Q(\u2/uk/K_r8 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[55] ),
        .Q(\u2/uk/K_r8 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[5] ),
        .Q(\u2/uk/K_r8 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[6] ),
        .Q(\u2/uk/K_r8 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[7] ),
        .Q(\u2/uk/K_r8 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[8] ),
        .Q(\u2/uk/K_r8 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r8_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r7_reg_n_0_[9] ),
        .Q(\u2/uk/K_r8 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [0]),
        .Q(\u2/uk/K_r9 [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [10]),
        .Q(\u2/uk/K_r9 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [11]),
        .Q(\u2/uk/K_r9 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [12]),
        .Q(\u2/uk/K_r9 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [13]),
        .Q(\u2/uk/K_r9 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [14]),
        .Q(\u2/uk/K_r9 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [15]),
        .Q(\u2/uk/K_r9 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [16]),
        .Q(\u2/uk/K_r9 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [17]),
        .Q(\u2/uk/K_r9 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [18]),
        .Q(\u2/uk/K_r9 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [19]),
        .Q(\u2/uk/K_r9 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [1]),
        .Q(\u2/uk/K_r9 [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [20]),
        .Q(\u2/uk/K_r9 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [21]),
        .Q(\u2/uk/K_r9 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [22]),
        .Q(\u2/uk/K_r9 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [23]),
        .Q(\u2/uk/K_r9 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [24]),
        .Q(\u2/uk/K_r9 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [25]),
        .Q(\u2/uk/K_r9 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [26]),
        .Q(\u2/uk/K_r9 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [27]),
        .Q(\u2/uk/K_r9 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [28]),
        .Q(\u2/uk/K_r9 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [29]),
        .Q(\u2/uk/K_r9 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [2]),
        .Q(\u2/uk/K_r9 [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [30]),
        .Q(\u2/uk/K_r9 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [31]),
        .Q(\u2/uk/K_r9 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [32]),
        .Q(\u2/uk/K_r9 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [33]),
        .Q(\u2/uk/K_r9 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [34]),
        .Q(\u2/uk/K_r9 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [35]),
        .Q(\u2/uk/K_r9 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [36]),
        .Q(\u2/uk/K_r9 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [37]),
        .Q(\u2/uk/K_r9 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [38]),
        .Q(\u2/uk/K_r9 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [39]),
        .Q(\u2/uk/K_r9 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [3]),
        .Q(\u2/uk/K_r9 [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [40]),
        .Q(\u2/uk/K_r9 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [41]),
        .Q(\u2/uk/K_r9 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [42]),
        .Q(\u2/uk/K_r9 [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [43]),
        .Q(\u2/uk/K_r9 [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [44]),
        .Q(\u2/uk/K_r9 [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [45]),
        .Q(\u2/uk/K_r9 [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [46]),
        .Q(\u2/uk/K_r9 [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [47]),
        .Q(\u2/uk/K_r9 [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [48]),
        .Q(\u2/uk/K_r9 [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [49]),
        .Q(\u2/uk/K_r9 [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [4]),
        .Q(\u2/uk/K_r9 [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [50]),
        .Q(\u2/uk/K_r9 [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [51]),
        .Q(\u2/uk/K_r9 [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [52]),
        .Q(\u2/uk/K_r9 [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [53]),
        .Q(\u2/uk/K_r9 [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [54]),
        .Q(\u2/uk/K_r9 [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [55]),
        .Q(\u2/uk/K_r9 [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [5]),
        .Q(\u2/uk/K_r9 [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [6]),
        .Q(\u2/uk/K_r9 [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [7]),
        .Q(\u2/uk/K_r9 [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [8]),
        .Q(\u2/uk/K_r9 [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \u2/uk/K_r9_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\u2/uk/K_r8 [9]),
        .Q(\u2/uk/K_r9 [9]),
        .R(\<const0>__0__0 ));
endmodule
