module msp430_vhdl
   (clk,
    rst,
    addr,
    din,
    dout,
    rd,
    wr,
    lbe,
    hbe,
    irq,
    iack,
    halt);
  input clk;
  input rst;
  output [15:1]addr;
  input [15:0]din;
  output [15:0]dout;
  output rd;
  output wr;
  output lbe;
  output hbe;
  input [14:0]irq;
  output [14:0]iack;
  input halt;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire FSM_sequential_state;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[0]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_state[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:8]L;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:1]addr;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_1_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[10]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_18_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_18_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_18_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_19_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_19_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_19_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_1_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_24_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_24_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_24_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_24_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_24_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_24_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_24_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_25_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_25_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_25_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[11]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[12]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[13]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[14]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_38_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_38_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_38_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_38_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[15]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[1]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[2]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_18_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_18_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_18_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_23_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_23_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_23_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_23_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_23_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_23_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_23_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_24_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_24_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_24_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[3]_INST_0_i_9_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_7_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[4]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[5]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[6]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_18_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_18_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_18_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_23_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_23_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_23_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_23_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_23_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_23_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_23_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_24_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_24_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_24_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[7]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[8]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \addr[9]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]as;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]bsaddr;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \bsaddr[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]bsaddr__0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire bw;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]data3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]data4;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]din;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]doc;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]dout;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[0]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[10]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_8_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_8_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_8_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_8_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[11]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[12]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[12]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[12]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[12]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[12]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[12]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[12]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[12]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[12]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[12]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[12]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[12]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_10_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_10_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_10_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_10_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_20_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[13]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_18_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_29_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[14]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_100_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_101_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_102_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_103_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_104_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_109_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_21_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_21_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_21_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_21_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_21_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_21_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_21_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_25_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_25_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_25_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_25_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_25_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_25_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_25_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_26_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_26_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_26_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_26_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_26_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_26_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_26_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_28_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_28_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_28_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_28_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_28_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_28_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_29_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_29_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_29_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_29_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_29_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_29_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_29_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_30_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_30_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_30_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_30_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_30_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_30_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_30_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_39_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_39_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_39_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_39_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_39_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_39_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_39_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_51_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_51_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_51_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_51_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_51_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_51_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_51_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_56_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_56_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_56_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_56_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_56_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_56_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_56_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_61_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_61_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_61_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_61_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_61_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_61_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_61_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_66_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_66_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_66_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_66_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_66_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_66_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_66_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_71_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_71_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_71_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_71_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_71_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_71_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_71_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_80_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_95_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_96_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_97_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_99_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[15]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[1]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[1]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[1]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[1]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[1]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[1]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[1]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[1]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[1]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[1]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_11_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_11_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_11_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_11_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_30_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_30_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_30_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_30_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_30_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_30_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_30_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_31_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_31_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_31_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_31_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_31_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_31_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_31_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_6_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_6_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_6_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_6_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_7_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_7_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_7_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_7_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[2]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_5_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[3]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_11_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_11_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_11_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_11_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_16_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_43_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_43_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_43_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_43_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_43_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_43_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_43_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_44_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_44_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_44_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_44_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_44_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_44_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_44_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_6_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_6_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_6_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_6_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_8_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_8_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_8_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_8_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[4]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_12_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[5]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_1_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_7_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[6]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_7_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[7]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[8]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[8]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[8]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[8]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[8]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[8]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[8]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[8]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[8]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[8]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[8]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[8]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_22_n_0_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \dout[9]_INST_0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire eqOp105_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire eqOp113_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire eqOp135_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire eqOp93_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire girq;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire halt;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hbe;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]iack;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[14]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[14]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[14]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \iack[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]irq;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:1]irqaddr;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire irqaddr0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqaddr[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqaddr[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqaddr[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqaddr[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqaddr[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqaddr[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqaddr[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqaddr[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lbe_INST_0_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]nstate;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire nstate1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in6_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_13_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_1_in108_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_1_in122_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_2_in88_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_4_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]pc;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]pc_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[11]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[11]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[11]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[11]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[15]_i_7_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[15]_i_7_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[15]_i_7_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[15]_i_7_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[3]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \pc_reg[7]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]plusOp;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]plusOp2_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]plusOp3_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]plusOp4_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[10][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[11][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[12][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[13][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[14][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[15][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[4][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[5][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[6][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[7][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[8][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[9][8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_a0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]r_code;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_code[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_code[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_code[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_code[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_code[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_code[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]r_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\r_reg[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[10][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\r_reg[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[11][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\r_reg[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[12][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\r_reg[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[13][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\r_reg[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[14][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\r_reg[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[15][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\r_reg[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[4][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\r_reg[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[5][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\r_reg[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[6][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\r_reg[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[7][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\r_reg[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[8][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\r_reg[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[9][8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_47_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_48_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_49_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_50_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_51_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_52_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_53_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_54_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_57_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_58_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_60_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_61_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_63_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_64_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_65_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_66_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_67_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_69_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_70_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rd_INST_0_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:1]\rrd[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rrs;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [13:0]\rrs[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rrs[0][4]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \rrs[0][7]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rst;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [2:0]soc;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sp;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sp19_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[0]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]sp_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[0]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[0]_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[0]_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[0]_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[4]_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[4]_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[4]_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[8]_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[8]_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sp_reg[8]_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sr;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sr1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[8]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[8]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[8]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[8]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]sr_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg[0]_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sr_reg_n_0_;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire src;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire src0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \src[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \src[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]src__0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]state;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \state[0]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \state[2]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \state[3]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \state[4]_repN ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]state_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire wr;

  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000AAAAAA2A)) 
    \FSM_sequential_state[0]_i_1 
       (.I0(\FSM_sequential_state[0]_i_2_n_0 ),
        .I1(state[0]),
        .I2(eqOp105_in),
        .I3(\FSM_sequential_state[0]_i_4_n_0 ),
        .I4(\FSM_sequential_state[0]_i_5_n_0 ),
        .I5(\FSM_sequential_state[0]_i_6_n_0 ),
        .O(\FSM_sequential_state[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAC0CC)) 
    \FSM_sequential_state[0]_i_10 
       (.I0(rd_INST_0_i_16_n_0),
        .I1(eqOp135_in),
        .I2(soc[1]),
        .I3(soc[2]),
        .I4(state[1]),
        .I5(state[2]),
        .O(FSM_sequential_state));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FF07FFFF)) 
    \FSM_sequential_state[0]_i_11 
       (.I0(nstate1),
        .I1(rd_INST_0_i_19_n_0),
        .I2(\FSM_sequential_state[3]_i_8_n_0 ),
        .I3(\FSM_sequential_state[0]_i_12_n_0 ),
        .I4(eqOp135_in),
        .I5(\FSM_sequential_state[0]_i_13_n_0 ),
        .O(\FSM_sequential_state[0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \FSM_sequential_state[0]_i_12 
       (.I0(state[1]),
        .I1(state[0]),
        .O(\FSM_sequential_state[0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000002F20202)) 
    \FSM_sequential_state[0]_i_13 
       (.I0(eqOp93_in),
        .I1(girq),
        .I2(eqOp135_in),
        .I3(eqOp113_in),
        .I4(rd_INST_0_i_19_n_0),
        .I5(state[1]),
        .O(\FSM_sequential_state[0]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF5455)) 
    \FSM_sequential_state[0]_i_2 
       (.I0(\sr_reg_n_0_[4] ),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\addr[15]_INST_0_i_11_n_0 ),
        .I4(\FSM_sequential_state[0]_i_7_n_0 ),
        .I5(girq),
        .O(\FSM_sequential_state[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000CCCCC4CC)) 
    \FSM_sequential_state[0]_i_3 
       (.I0(soc[1]),
        .I1(as[0]),
        .I2(\r_code[11]_i_1_n_0 ),
        .I3(soc[2]),
        .I4(\r_code[10]_i_1_n_0 ),
        .I5(as[1]),
        .O(eqOp105_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_state[0]_i_4 
       (.I0(rd_INST_0_i_16_n_0),
        .I1(rd_INST_0_i_21_n_0),
        .O(\FSM_sequential_state[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFB)) 
    \FSM_sequential_state[0]_i_5 
       (.I0(eqOp93_in),
        .I1(rd_INST_0_i_21_n_0),
        .I2(eqOp135_in),
        .I3(\dout[13]_INST_0_i_3_n_0 ),
        .I4(state[2]),
        .I5(state[1]),
        .O(\FSM_sequential_state[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFEFFFEFFFE0000)) 
    \FSM_sequential_state[0]_i_6 
       (.I0(state[2]),
        .I1(state[3]),
        .I2(state[0]),
        .I3(state[1]),
        .I4(\FSM_sequential_state[0]_i_8_n_0 ),
        .I5(state[4]),
        .O(\FSM_sequential_state[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h03AF030FFFAFFFAF)) 
    \FSM_sequential_state[0]_i_7 
       (.I0(\FSM_sequential_state[0]_i_9_n_0 ),
        .I1(state[2]),
        .I2(state[0]),
        .I3(state[1]),
        .I4(rd_INST_0_i_19_n_0),
        .I5(FSM_sequential_state),
        .O(\FSM_sequential_state[0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC4D40D70D4D47D7D)) 
    \FSM_sequential_state[0]_i_8 
       (.I0(girq),
        .I1(state[0]),
        .I2(state[1]),
        .I3(state[3]),
        .I4(state[2]),
        .I5(\FSM_sequential_state[0]_i_11_n_0 ),
        .O(\FSM_sequential_state[0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFEFF)) 
    \FSM_sequential_state[0]_i_9 
       (.I0(\dout[13]_INST_0_i_3_n_0 ),
        .I1(eqOp135_in),
        .I2(rd_INST_0_i_21_n_0),
        .I3(rd_INST_0_i_16_n_0),
        .O(\FSM_sequential_state[0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEFEEEEEEEEEEE)) 
    \FSM_sequential_state[1]_i_1 
       (.I0(\FSM_sequential_state[1]_i_2_n_0 ),
        .I1(\FSM_sequential_state[1]_i_3_n_0 ),
        .I2(\FSM_sequential_state[1]_i_4_n_0 ),
        .I3(\FSM_sequential_state[1]_i_5_n_0 ),
        .I4(state[4]),
        .I5(state[0]),
        .O(\FSM_sequential_state[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_state[1]_i_10 
       (.I0(state[3]),
        .I1(rd_INST_0_i_16_n_0),
        .O(\FSM_sequential_state[1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00AA00AE)) 
    \FSM_sequential_state[1]_i_11 
       (.I0(eqOp93_in),
        .I1(rd_INST_0_i_16_n_0),
        .I2(rd_INST_0_i_21_n_0),
        .I3(eqOp135_in),
        .I4(\dout[13]_INST_0_i_3_n_0 ),
        .O(\FSM_sequential_state[1]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_state[1]_i_12 
       (.I0(eqOp135_in),
        .I1(rd_INST_0_i_19_n_0),
        .O(\FSM_sequential_state[1]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_state[1]_i_13 
       (.I0(state[0]),
        .I1(state[4]),
        .O(\FSM_sequential_state[1]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF67660000)) 
    \FSM_sequential_state[1]_i_2 
       (.I0(state[4]),
        .I1(state[3]),
        .I2(\FSM_sequential_state[1]_i_6_n_0 ),
        .I3(\FSM_sequential_state[1]_i_7_n_0 ),
        .I4(\FSM_sequential_state[1]_i_8_n_0 ),
        .I5(\FSM_sequential_state[1]_i_9_n_0 ),
        .O(\FSM_sequential_state[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0101010000000200)) 
    \FSM_sequential_state[1]_i_3 
       (.I0(state[3]),
        .I1(state[1]),
        .I2(state[4]),
        .I3(\sr_reg_n_0_[4] ),
        .I4(girq),
        .I5(state[2]),
        .O(\FSM_sequential_state[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0303030347474744)) 
    \FSM_sequential_state[1]_i_4 
       (.I0(state[4]),
        .I1(state[2]),
        .I2(\FSM_sequential_state[1]_i_10_n_0 ),
        .I3(\FSM_sequential_state[1]_i_11_n_0 ),
        .I4(\FSM_sequential_state[1]_i_12_n_0 ),
        .I5(state[1]),
        .O(\FSM_sequential_state[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_state[1]_i_5 
       (.I0(\sr_reg_n_0_[4] ),
        .I1(girq),
        .O(\FSM_sequential_state[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0C0080CC8CCC80CC)) 
    \FSM_sequential_state[1]_i_6 
       (.I0(soc[0]),
        .I1(eqOp135_in),
        .I2(soc[1]),
        .I3(soc[2]),
        .I4(rd_INST_0_i_19_n_0),
        .I5(eqOp113_in),
        .O(\FSM_sequential_state[1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBAABAA)) 
    \FSM_sequential_state[1]_i_7 
       (.I0(eqOp135_in),
        .I1(eqOp93_in),
        .I2(\dout[13]_INST_0_i_3_n_0 ),
        .I3(rd_INST_0_i_21_n_0),
        .I4(state[1]),
        .O(\FSM_sequential_state[1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \FSM_sequential_state[1]_i_8 
       (.I0(state[2]),
        .I1(state[0]),
        .I2(state[1]),
        .O(\FSM_sequential_state[1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040004045400540)) 
    \FSM_sequential_state[1]_i_9 
       (.I0(\FSM_sequential_state[1]_i_13_n_0 ),
        .I1(state[1]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(\sr_reg_n_0_[4] ),
        .I5(girq),
        .O(\FSM_sequential_state[1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3111)) 
    \FSM_sequential_state[2]_i_1 
       (.I0(\FSM_sequential_state[2]_i_2_n_0 ),
        .I1(state[4]),
        .I2(state[0]),
        .I3(\FSM_sequential_state[2]_i_3_n_0 ),
        .O(\FSM_sequential_state[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8FA8F8F8FBF)) 
    \FSM_sequential_state[2]_i_2 
       (.I0(state[0]),
        .I1(state[2]),
        .I2(state[3]),
        .I3(girq),
        .I4(\sr_reg_n_0_[4] ),
        .I5(state[1]),
        .O(\FSM_sequential_state[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000F0FFF008C0FFF)) 
    \FSM_sequential_state[2]_i_3 
       (.I0(rd_INST_0_i_19_n_0),
        .I1(\FSM_sequential_state[2]_i_4_n_0 ),
        .I2(\FSM_sequential_state[2]_i_5_n_0 ),
        .I3(state[1]),
        .I4(\FSM_sequential_state[2]_i_6_n_0 ),
        .I5(state[2]),
        .O(\FSM_sequential_state[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8FFF8F8F88888888)) 
    \FSM_sequential_state[2]_i_4 
       (.I0(\FSM_sequential_state[2]_i_7_n_0 ),
        .I1(\FSM_sequential_state[3]_i_7_n_0 ),
        .I2(\FSM_sequential_state[2]_i_5_n_0 ),
        .I3(eqOp93_in),
        .I4(state[2]),
        .I5(\FSM_sequential_state[1]_i_11_n_0 ),
        .O(\FSM_sequential_state[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_state[2]_i_5 
       (.I0(girq),
        .I1(\sr_reg_n_0_[4] ),
        .O(\FSM_sequential_state[2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4FF)) 
    \FSM_sequential_state[2]_i_6 
       (.I0(rd_INST_0_i_16_n_0),
        .I1(state[1]),
        .I2(state[2]),
        .I3(state[3]),
        .O(\FSM_sequential_state[2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88AAA0AA)) 
    \FSM_sequential_state[2]_i_7 
       (.I0(eqOp135_in),
        .I1(soc[0]),
        .I2(rd_INST_0_i_19_n_0),
        .I3(soc[2]),
        .I4(soc[1]),
        .O(\FSM_sequential_state[2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000F000FDD)) 
    \FSM_sequential_state[3]_i_1 
       (.I0(\FSM_sequential_state[3]_i_2_n_0 ),
        .I1(\FSM_sequential_state[3]_i_3_n_0 ),
        .I2(\FSM_sequential_state[3]_i_4_n_0 ),
        .I3(state[2]),
        .I4(\FSM_sequential_state[3]_i_5_n_0 ),
        .I5(state[4]),
        .O(\FSM_sequential_state[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEAEE00FF)) 
    \FSM_sequential_state[3]_i_2 
       (.I0(state[2]),
        .I1(state[0]),
        .I2(rd_INST_0_i_16_n_0),
        .I3(state[3]),
        .I4(state[1]),
        .O(\FSM_sequential_state[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001000100015501)) 
    \FSM_sequential_state[3]_i_3 
       (.I0(state[1]),
        .I1(\FSM_sequential_state[3]_i_6_n_0 ),
        .I2(eqOp93_in),
        .I3(eqOp135_in),
        .I4(\FSM_sequential_state[3]_i_7_n_0 ),
        .I5(\FSM_sequential_state[3]_i_8_n_0 ),
        .O(\FSM_sequential_state[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFA1F)) 
    \FSM_sequential_state[3]_i_4 
       (.I0(state[1]),
        .I1(girq),
        .I2(state[0]),
        .I3(state[3]),
        .O(\FSM_sequential_state[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_state[3]_i_5 
       (.I0(state[0]),
        .I1(state[1]),
        .O(\FSM_sequential_state[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBA)) 
    \FSM_sequential_state[3]_i_6 
       (.I0(\dout[13]_INST_0_i_3_n_0 ),
        .I1(rd_INST_0_i_21_n_0),
        .I2(rd_INST_0_i_16_n_0),
        .O(\FSM_sequential_state[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFD5)) 
    \FSM_sequential_state[3]_i_7 
       (.I0(as[1]),
        .I1(\addr[15]_INST_0_i_11_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(nstate1),
        .O(\FSM_sequential_state[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000505030000000)) 
    \FSM_sequential_state[3]_i_8 
       (.I0(r_code[7]),
        .I1(din[7]),
        .I2(soc[1]),
        .I3(din[9]),
        .I4(p_2_in88_in),
        .I5(r_code[9]),
        .O(\FSM_sequential_state[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \FSM_sequential_state[4]_i_1 
       (.I0(halt),
        .O(\FSM_sequential_state[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h08100010)) 
    \FSM_sequential_state[4]_i_2 
       (.I0(state[3]),
        .I1(state[2]),
        .I2(state[4]),
        .I3(state[1]),
        .I4(state[0]),
        .O(\FSM_sequential_state[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \FSM_sequential_state[4]_i_3 
       (.I0(rst),
        .O(\FSM_sequential_state[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \FSM_sequential_state_reg[0] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .D(\FSM_sequential_state[0]_i_1_n_0 ),
        .PRE(\FSM_sequential_state[4]_i_3_n_0 ),
        .Q(state[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "FSM_sequential_state_reg[0]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \FSM_sequential_state_reg[0]_replica 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .D(\FSM_sequential_state[0]_i_1_n_0 ),
        .PRE(\FSM_sequential_state[4]_i_3_n_0 ),
        .Q(\state[0]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \FSM_sequential_state_reg[1] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\FSM_sequential_state[1]_i_1_n_0 ),
        .Q(state[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \FSM_sequential_state_reg[2] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\FSM_sequential_state[2]_i_1_n_0 ),
        .Q(state[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "FSM_sequential_state_reg[2]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \FSM_sequential_state_reg[2]_replica 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\FSM_sequential_state[2]_i_1_n_0 ),
        .Q(\state[2]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \FSM_sequential_state_reg[3] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\FSM_sequential_state[3]_i_1_n_0 ),
        .Q(state[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "FSM_sequential_state_reg[3]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \FSM_sequential_state_reg[3]_replica 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\FSM_sequential_state[3]_i_1_n_0 ),
        .Q(\state[3]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \FSM_sequential_state_reg[4] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .D(\FSM_sequential_state[4]_i_2_n_0 ),
        .PRE(\FSM_sequential_state[4]_i_3_n_0 ),
        .Q(state[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "FSM_sequential_state_reg[4]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \FSM_sequential_state_reg[4]_replica 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .D(\FSM_sequential_state[4]_i_2_n_0 ),
        .PRE(\FSM_sequential_state[4]_i_3_n_0 ),
        .Q(\state[4]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1F11)) 
    \addr[10]_INST_0 
       (.I0(\addr[15]_INST_0_i_1_n_0 ),
        .I1(\addr[10]_INST_0_i_1_n_0_repN ),
        .I2(\addr[15]_INST_0_i_3_n_0 ),
        .I3(sp_reg[10]),
        .I4(\addr[10]_INST_0_i_2_n_0 ),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(addr[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[10]_INST_0_i_10 
       (.I0(\r_reg[15] [10]),
        .I1(\r_reg[14] [10]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [10]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [10]),
        .O(\addr[10]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[10]_INST_0_i_11 
       (.I0(\r_reg[7] [10]),
        .I1(\r_reg[6] [10]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [10]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [10]),
        .O(\addr[10]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[10]_INST_0_i_12 
       (.I0(\addr[11]_INST_0_i_24_n_5 ),
        .I1(p_4_in),
        .I2(pc[10]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[10]),
        .O(\addr[10]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \addr[10]_INST_0_i_13 
       (.I0(\addr[10]_INST_0_i_15_n_0 ),
        .I1(\addr[10]_INST_0_i_16_n_0 ),
        .O(\addr[10]_INST_0_i_13_n_0 ),
        .S(\r_code[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \addr[10]_INST_0_i_14 
       (.I0(\addr[10]_INST_0_i_17_n_0 ),
        .I1(\addr[10]_INST_0_i_18_n_0 ),
        .O(\addr[10]_INST_0_i_14_n_0 ),
        .S(\r_code[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5F503F3F5F503030)) 
    \addr[10]_INST_0_i_15 
       (.I0(\addr[15]_INST_0_i_20_n_0 ),
        .I1(\addr[10]_INST_0_i_5_n_0 ),
        .I2(soc[2]),
        .I3(sp_reg[10]),
        .I4(soc[1]),
        .I5(pc[10]),
        .O(\addr[10]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[10]_INST_0_i_16 
       (.I0(\r_reg[7] [10]),
        .I1(\r_reg[6] [10]),
        .I2(soc[2]),
        .I3(\r_reg[5] [10]),
        .I4(soc[1]),
        .I5(\r_reg[4] [10]),
        .O(\addr[10]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[10]_INST_0_i_17 
       (.I0(\r_reg[11] [10]),
        .I1(\r_reg[10] [10]),
        .I2(soc[2]),
        .I3(\r_reg[9] [10]),
        .I4(soc[1]),
        .I5(\r_reg[8] [10]),
        .O(\addr[10]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[10]_INST_0_i_18 
       (.I0(\r_reg[15] [10]),
        .I1(\r_reg[14] [10]),
        .I2(soc[2]),
        .I3(\r_reg[13] [10]),
        .I4(soc[1]),
        .I5(\r_reg[12] [10]),
        .O(\addr[10]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "addr[10]_INST_0_i_1" *) 
  LUT6 #(
    .INIT(64'h0000000011101111)) 
    \addr[10]_INST_0_i_1_replica 
       (.I0(\addr[10]_INST_0_i_3_n_0 ),
        .I1(\addr[10]_INST_0_i_4_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\addr[10]_INST_0_i_5_n_0 ),
        .I4(\addr[14]_INST_0_i_5_n_0 ),
        .I5(\addr[10]_INST_0_i_6_n_0 ),
        .O(\addr[10]_INST_0_i_1_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00005455)) 
    \addr[10]_INST_0_i_1_rewire 
       (.I0(\addr[10]_INST_0_i_3_n_0 ),
        .I1(\r_code[3]_i_1_n_0 ),
        .I2(\addr[10]_INST_0_i_5_n_0 ),
        .I3(\addr[14]_INST_0_i_5_n_0 ),
        .I4(\addr[10]_INST_0_i_6_n_0 ),
        .O(\addr[10]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    \addr[10]_INST_0_i_2 
       (.I0(data3[10]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[10]_INST_0_i_7_n_0 ),
        .I3(\addr[15]_INST_0_i_17_n_0 ),
        .I4(\addr[10]_INST_0_i_8_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[10]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEA202A00000000)) 
    \addr[10]_INST_0_i_3 
       (.I0(\addr[10]_INST_0_i_9_n_0 ),
        .I1(din[2]),
        .I2(p_2_in88_in),
        .I3(r_code[2]),
        .I4(\addr[10]_INST_0_i_10_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\addr[10]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA0000A808)) 
    \addr[10]_INST_0_i_4 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(pc[10]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(sp_reg[10]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_9_n_0 ),
        .O(\addr[10]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFBBFCB8FFFFFFFF)) 
    \addr[10]_INST_0_i_5 
       (.I0(din[4]),
        .I1(p_2_in88_in),
        .I2(r_code[4]),
        .I3(din[5]),
        .I4(r_code[5]),
        .I5(\sr_reg_n_0_[10] ),
        .O(\addr[10]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000505030000000)) 
    \addr[10]_INST_0_i_6 
       (.I0(r_code[3]),
        .I1(din[3]),
        .I2(\addr[10]_INST_0_i_11_n_0 ),
        .I3(din[2]),
        .I4(p_2_in88_in),
        .I5(r_code[2]),
        .O(\addr[10]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[10]_INST_0_i_7 
       (.I0(\addr[10]_INST_0_i_12_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[10]),
        .I3(state[0]),
        .I4(plusOp4_out[10]),
        .O(\addr[10]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \addr[10]_INST_0_i_8 
       (.I0(\addr[10]_INST_0_i_13_n_0 ),
        .I1(\addr[10]_INST_0_i_14_n_0 ),
        .O(\addr[10]_INST_0_i_8_n_0 ),
        .S(\r_code[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[10]_INST_0_i_9 
       (.I0(\r_reg[11] [10]),
        .I1(\r_reg[10] [10]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [10]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [10]),
        .O(\addr[10]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1F11)) 
    \addr[11]_INST_0 
       (.I0(\addr[15]_INST_0_i_1_n_0 ),
        .I1(\addr[11]_INST_0_i_1_n_0_repN ),
        .I2(\addr[15]_INST_0_i_3_n_0 ),
        .I3(sp_reg[11]),
        .I4(\addr[11]_INST_0_i_2_n_0 ),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(addr[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[11]_INST_0_i_10 
       (.I0(\r_reg[11] [11]),
        .I1(\r_reg[10] [11]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [11]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [11]),
        .O(\addr[11]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[11]_INST_0_i_11 
       (.I0(\r_reg[15] [11]),
        .I1(\r_reg[14] [11]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [11]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [11]),
        .O(\addr[11]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[11]_INST_0_i_12 
       (.I0(\r_reg[7] [11]),
        .I1(\r_reg[6] [11]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [11]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [11]),
        .O(\addr[11]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h63)) 
    \addr[11]_INST_0_i_13_rewire 
       (.I0(\addr[11]_INST_0_i_4_n_0 ),
        .I1(din[11]),
        .I2(\addr[11]_INST_0_i_1_n_0 ),
        .O(\addr[11]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h63)) 
    \addr[11]_INST_0_i_14_rewire 
       (.I0(\addr[10]_INST_0_i_4_n_0 ),
        .I1(din[10]),
        .I2(\addr[10]_INST_0_i_1_n_0 ),
        .O(\addr[11]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[11]_INST_0_i_15 
       (.I0(din[9]),
        .I1(\rrs[0] [9]),
        .O(\addr[11]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[11]_INST_0_i_16 
       (.I0(din[8]),
        .I1(\rrs[0] [8]),
        .O(\addr[11]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[11]_INST_0_i_17 
       (.I0(\addr[11]_INST_0_i_24_n_4 ),
        .I1(p_4_in),
        .I2(pc[11]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[11]),
        .O(\addr[11]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[11]_INST_0_i_18 
       (.CI(\addr[7]_INST_0_i_17_n_0 ),
        .CO({\addr[11]_INST_0_i_18_n_0 ,\addr[11]_INST_0_i_18_n_1 ,\addr[11]_INST_0_i_18_n_2 ,\addr[11]_INST_0_i_18_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(din[11:8]),
        .O(plusOp3_out[11:8]),
        .S({\addr[11]_INST_0_i_26_n_0 ,\addr[11]_INST_0_i_27_n_0 ,\addr[11]_INST_0_i_28_n_0 ,\addr[11]_INST_0_i_29_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[11]_INST_0_i_19 
       (.CI(\addr[7]_INST_0_i_18_n_0 ),
        .CO({\addr[11]_INST_0_i_19_n_0 ,\addr[11]_INST_0_i_19_n_1 ,\addr[11]_INST_0_i_19_n_2 ,\addr[11]_INST_0_i_19_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(din[11:8]),
        .O(plusOp4_out[11:8]),
        .S({\addr[11]_INST_0_i_30_n_0 ,\addr[11]_INST_0_i_31_n_0 ,\addr[11]_INST_0_i_32_n_0 ,\addr[11]_INST_0_i_33_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "addr[11]_INST_0_i_1" *) 
  LUT6 #(
    .INIT(64'h0000000011101111)) 
    \addr[11]_INST_0_i_1_replica 
       (.I0(\addr[11]_INST_0_i_3_n_0 ),
        .I1(\addr[11]_INST_0_i_4_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\addr[11]_INST_0_i_5_n_0 ),
        .I4(\addr[14]_INST_0_i_5_n_0 ),
        .I5(\addr[11]_INST_0_i_6_n_0 ),
        .O(\addr[11]_INST_0_i_1_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00005455)) 
    \addr[11]_INST_0_i_1_rewire 
       (.I0(\addr[11]_INST_0_i_3_n_0 ),
        .I1(\r_code[3]_i_1_n_0 ),
        .I2(\addr[11]_INST_0_i_5_n_0 ),
        .I3(\addr[14]_INST_0_i_5_n_0 ),
        .I4(\addr[11]_INST_0_i_6_n_0 ),
        .O(\addr[11]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000FFB8B8)) 
    \addr[11]_INST_0_i_2 
       (.I0(data3[11]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[11]_INST_0_i_8_n_0 ),
        .I3(\addr[11]_INST_0_i_9_n_0 ),
        .I4(\addr[15]_INST_0_i_17_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[11]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000002022220020)) 
    \addr[11]_INST_0_i_20 
       (.I0(soc[2]),
        .I1(\r_code[10]_i_1_n_0 ),
        .I2(\sr_reg_n_0_[11] ),
        .I3(lbe_INST_0_i_8_n_0),
        .I4(soc[1]),
        .I5(\addr[15]_INST_0_i_20_n_0 ),
        .O(\addr[11]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA3A3A3A0A0A3A0A0)) 
    \addr[11]_INST_0_i_21 
       (.I0(\addr[11]_INST_0_i_34_n_0 ),
        .I1(soc[2]),
        .I2(\r_code[10]_i_1_n_0 ),
        .I3(soc[1]),
        .I4(pc[11]),
        .I5(sp_reg[11]),
        .O(\addr[11]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[11]_INST_0_i_22 
       (.I0(\r_reg[15] [11]),
        .I1(\r_reg[14] [11]),
        .I2(soc[2]),
        .I3(\r_reg[13] [11]),
        .I4(soc[1]),
        .I5(\r_reg[12] [11]),
        .O(\addr[11]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[11]_INST_0_i_23 
       (.I0(\r_reg[11] [11]),
        .I1(\r_reg[10] [11]),
        .I2(soc[2]),
        .I3(\r_reg[9] [11]),
        .I4(soc[1]),
        .I5(\r_reg[8] [11]),
        .O(\addr[11]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[11]_INST_0_i_24 
       (.CI(\addr[7]_INST_0_i_23_n_0 ),
        .CO({\addr[11]_INST_0_i_24_n_0 ,\addr[11]_INST_0_i_24_n_1 ,\addr[11]_INST_0_i_24_n_2 ,\addr[11]_INST_0_i_24_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(bsaddr__0[11:8]),
        .O({\addr[11]_INST_0_i_24_n_4 ,\addr[11]_INST_0_i_24_n_5 ,\addr[11]_INST_0_i_24_n_6 ,\addr[11]_INST_0_i_24_n_7 }),
        .S({\addr[11]_INST_0_i_35_n_0 ,\addr[11]_INST_0_i_36_n_0 ,\addr[11]_INST_0_i_37_n_0 ,\addr[11]_INST_0_i_38_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[11]_INST_0_i_25 
       (.CI(\addr[7]_INST_0_i_24_n_0 ),
        .CO({\addr[11]_INST_0_i_25_n_0 ,\addr[11]_INST_0_i_25_n_1 ,\addr[11]_INST_0_i_25_n_2 ,\addr[11]_INST_0_i_25_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(bsaddr__0[11:8]),
        .O(plusOp2_out[11:8]),
        .S({\addr[11]_INST_0_i_39_n_0 ,\addr[11]_INST_0_i_40_n_0 ,\addr[11]_INST_0_i_41_n_0 ,\addr[11]_INST_0_i_42_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[11]_INST_0_i_26 
       (.I0(din[11]),
        .I1(\rrd[0] [11]),
        .O(\addr[11]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[11]_INST_0_i_27 
       (.I0(din[10]),
        .I1(\rrd[0] [10]),
        .O(\addr[11]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[11]_INST_0_i_28 
       (.I0(din[9]),
        .I1(\rrd[0] [9]),
        .O(\addr[11]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[11]_INST_0_i_29 
       (.I0(din[8]),
        .I1(\rrd[0] [8]),
        .O(\addr[11]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEA202A00000000)) 
    \addr[11]_INST_0_i_3 
       (.I0(\addr[11]_INST_0_i_10_n_0 ),
        .I1(din[2]),
        .I2(p_2_in88_in),
        .I3(r_code[2]),
        .I4(\addr[11]_INST_0_i_11_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\addr[11]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[11]_INST_0_i_30 
       (.I0(din[11]),
        .I1(\addr[11]_INST_0_i_9_n_0 ),
        .O(\addr[11]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[11]_INST_0_i_31 
       (.I0(din[10]),
        .I1(\addr[10]_INST_0_i_8_n_0 ),
        .O(\addr[11]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[11]_INST_0_i_32 
       (.I0(din[9]),
        .I1(\addr[9]_INST_0_i_8_n_0 ),
        .O(\addr[11]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[11]_INST_0_i_33 
       (.I0(din[8]),
        .I1(\addr[8]_INST_0_i_8_n_0 ),
        .O(\addr[11]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[11]_INST_0_i_34 
       (.I0(\r_reg[7] [11]),
        .I1(\r_reg[6] [11]),
        .I2(soc[2]),
        .I3(\r_reg[5] [11]),
        .I4(soc[1]),
        .I5(\r_reg[4] [11]),
        .O(\addr[11]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[11]_INST_0_i_35 
       (.I0(bsaddr__0[11]),
        .I1(\addr[11]_INST_0_i_9_n_0 ),
        .O(\addr[11]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[11]_INST_0_i_36 
       (.I0(bsaddr__0[10]),
        .I1(\addr[10]_INST_0_i_8_n_0 ),
        .O(\addr[11]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[11]_INST_0_i_37 
       (.I0(bsaddr__0[9]),
        .I1(\addr[9]_INST_0_i_8_n_0 ),
        .O(\addr[11]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[11]_INST_0_i_38 
       (.I0(bsaddr__0[8]),
        .I1(\addr[8]_INST_0_i_8_n_0 ),
        .O(\addr[11]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h63)) 
    \addr[11]_INST_0_i_39_rewire 
       (.I0(\addr[11]_INST_0_i_4_n_0 ),
        .I1(bsaddr__0[11]),
        .I2(\addr[11]_INST_0_i_1_n_0 ),
        .O(\addr[11]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA0000A808)) 
    \addr[11]_INST_0_i_4 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(pc[11]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(sp_reg[11]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_9_n_0 ),
        .O(\addr[11]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h63)) 
    \addr[11]_INST_0_i_40_rewire 
       (.I0(\addr[10]_INST_0_i_4_n_0 ),
        .I1(bsaddr__0[10]),
        .I2(\addr[10]_INST_0_i_1_n_0 ),
        .O(\addr[11]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[11]_INST_0_i_41 
       (.I0(bsaddr__0[9]),
        .I1(\rrs[0] [9]),
        .O(\addr[11]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[11]_INST_0_i_42 
       (.I0(bsaddr__0[8]),
        .I1(\rrs[0] [8]),
        .O(\addr[11]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEEAAA)) 
    \addr[11]_INST_0_i_43 
       (.I0(\addr[11]_INST_0_i_3_n_0 ),
        .I1(\addr[15]_INST_0_i_11_n_0 ),
        .I2(\addr[3]_INST_0_i_47_n_0 ),
        .I3(\sr_reg_n_0_[11] ),
        .I4(\addr[11]_INST_0_i_47_n_0 ),
        .I5(\addr[11]_INST_0_i_6_n_0 ),
        .O(\rrd[0] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEEAAA)) 
    \addr[11]_INST_0_i_44 
       (.I0(\addr[10]_INST_0_i_3_n_0 ),
        .I1(\addr[15]_INST_0_i_11_n_0 ),
        .I2(\sr_reg_n_0_[10] ),
        .I3(\addr[3]_INST_0_i_47_n_0 ),
        .I4(\addr[11]_INST_0_i_48_n_0 ),
        .I5(\addr[10]_INST_0_i_6_n_0 ),
        .O(\rrd[0] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEAEAEAFF)) 
    \addr[11]_INST_0_i_45 
       (.I0(\addr[9]_INST_0_i_6_n_0 ),
        .I1(\addr[15]_INST_0_i_11_n_0 ),
        .I2(\addr[11]_INST_0_i_49_n_0 ),
        .I3(\r_code[3]_i_1_n_0 ),
        .I4(\addr[9]_INST_0_i_3_n_0 ),
        .O(\rrd[0] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEAEAEAFF)) 
    \addr[11]_INST_0_i_46 
       (.I0(\addr[8]_INST_0_i_6_n_0 ),
        .I1(\addr[15]_INST_0_i_11_n_0 ),
        .I2(\addr[11]_INST_0_i_50_n_0 ),
        .I3(\r_code[3]_i_1_n_0 ),
        .I4(\addr[8]_INST_0_i_3_n_0 ),
        .O(\rrd[0] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \addr[11]_INST_0_i_47 
       (.I0(pc[11]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(sp_reg[11]),
        .I3(\r_code[1]_i_1_n_0 ),
        .O(\addr[11]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \addr[11]_INST_0_i_48 
       (.I0(pc[10]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(sp_reg[10]),
        .I3(\r_code[1]_i_1_n_0 ),
        .O(\addr[11]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF454045404540)) 
    \addr[11]_INST_0_i_49 
       (.I0(\r_code[1]_i_1_n_0 ),
        .I1(sp_reg[9]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(pc[9]),
        .I4(\addr[3]_INST_0_i_47_n_0 ),
        .I5(\sr_reg_n_0_[9] ),
        .O(\addr[11]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFBBFCB8FFFFFFFF)) 
    \addr[11]_INST_0_i_5 
       (.I0(din[4]),
        .I1(p_2_in88_in),
        .I2(r_code[4]),
        .I3(din[5]),
        .I4(r_code[5]),
        .I5(\sr_reg_n_0_[11] ),
        .O(\addr[11]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF454045404540)) 
    \addr[11]_INST_0_i_50 
       (.I0(\r_code[1]_i_1_n_0 ),
        .I1(sp_reg[8]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(pc[8]),
        .I4(\addr[3]_INST_0_i_47_n_0 ),
        .I5(\sr_reg_n_0_[8] ),
        .O(\addr[11]_INST_0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000505030000000)) 
    \addr[11]_INST_0_i_6 
       (.I0(r_code[3]),
        .I1(din[3]),
        .I2(\addr[11]_INST_0_i_12_n_0 ),
        .I3(din[2]),
        .I4(p_2_in88_in),
        .I5(r_code[2]),
        .O(\addr[11]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[11]_INST_0_i_7 
       (.CI(\addr[7]_INST_0_i_6_n_0 ),
        .CO({\addr[11]_INST_0_i_7_n_0 ,\addr[11]_INST_0_i_7_n_1 ,\addr[11]_INST_0_i_7_n_2 ,\addr[11]_INST_0_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(din[11:8]),
        .O(data3[11:8]),
        .S({\addr[11]_INST_0_i_13_n_0 ,\addr[11]_INST_0_i_14_n_0 ,\addr[11]_INST_0_i_15_n_0 ,\addr[11]_INST_0_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[11]_INST_0_i_8 
       (.I0(\addr[11]_INST_0_i_17_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[11]),
        .I3(state[0]),
        .I4(plusOp4_out[11]),
        .O(\addr[11]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0FFF00011111111)) 
    \addr[11]_INST_0_i_9 
       (.I0(\addr[11]_INST_0_i_20_n_0 ),
        .I1(\addr[11]_INST_0_i_21_n_0 ),
        .I2(\addr[11]_INST_0_i_22_n_0 ),
        .I3(\r_code[10]_i_1_n_0 ),
        .I4(\addr[11]_INST_0_i_23_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\addr[11]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4F44)) 
    \addr[12]_INST_0 
       (.I0(\addr[15]_INST_0_i_1_n_0 ),
        .I1(rrs),
        .I2(\addr[15]_INST_0_i_3_n_0 ),
        .I3(sp_reg[12]),
        .I4(\addr[12]_INST_0_i_2_n_0 ),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(addr[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[12]_INST_0_i_10 
       (.I0(\r_reg[15] [12]),
        .I1(\r_reg[14] [12]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [12]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [12]),
        .O(\addr[12]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[12]_INST_0_i_11 
       (.I0(\r_reg[7] [12]),
        .I1(\r_reg[6] [12]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [12]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [12]),
        .O(\addr[12]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[12]_INST_0_i_12 
       (.I0(\addr[15]_INST_0_i_38_n_7 ),
        .I1(p_4_in),
        .I2(pc[12]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[12]),
        .O(\addr[12]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[12]_INST_0_i_13 
       (.I0(\r_reg[15] [12]),
        .I1(\r_reg[14] [12]),
        .I2(soc[2]),
        .I3(\r_reg[13] [12]),
        .I4(soc[1]),
        .I5(\r_reg[12] [12]),
        .O(\addr[12]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[12]_INST_0_i_14 
       (.I0(\r_reg[11] [12]),
        .I1(\r_reg[10] [12]),
        .I2(soc[2]),
        .I3(\r_reg[9] [12]),
        .I4(soc[1]),
        .I5(\r_reg[8] [12]),
        .O(\addr[12]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[12]_INST_0_i_15 
       (.I0(\r_reg[7] [12]),
        .I1(\r_reg[6] [12]),
        .I2(soc[2]),
        .I3(\r_reg[5] [12]),
        .I4(soc[1]),
        .I5(\r_reg[4] [12]),
        .O(\addr[12]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF000F0FF55335533)) 
    \addr[12]_INST_0_i_16 
       (.I0(sp_reg[12]),
        .I1(pc[12]),
        .I2(\addr[15]_INST_0_i_20_n_0 ),
        .I3(soc[1]),
        .I4(\addr[12]_INST_0_i_5_n_0 ),
        .I5(soc[2]),
        .O(\addr[12]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "addr[12]_INST_0_i_1" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEFEEEEEE)) 
    \addr[12]_INST_0_i_1_replica 
       (.I0(\addr[12]_INST_0_i_3_n_0 ),
        .I1(\addr[12]_INST_0_i_4_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\addr[12]_INST_0_i_5_n_0 ),
        .I4(\addr[14]_INST_0_i_5_n_0 ),
        .I5(\addr[12]_INST_0_i_6_n_0 ),
        .O(rrs));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFBAAA)) 
    \addr[12]_INST_0_i_1_rewire 
       (.I0(\addr[12]_INST_0_i_3_n_0 ),
        .I1(\r_code[3]_i_1_n_0 ),
        .I2(\addr[12]_INST_0_i_5_n_0 ),
        .I3(\addr[14]_INST_0_i_5_n_0 ),
        .I4(\addr[12]_INST_0_i_6_n_0 ),
        .O(\rrs[0] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000FFB8B8)) 
    \addr[12]_INST_0_i_2 
       (.I0(data3[12]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[12]_INST_0_i_7_n_0 ),
        .I3(\addr[12]_INST_0_i_8_n_0 ),
        .I4(\addr[15]_INST_0_i_17_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[12]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEA202A00000000)) 
    \addr[12]_INST_0_i_3 
       (.I0(\addr[12]_INST_0_i_9_n_0 ),
        .I1(din[2]),
        .I2(p_2_in88_in),
        .I3(r_code[2]),
        .I4(\addr[12]_INST_0_i_10_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\addr[12]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA0000A808)) 
    \addr[12]_INST_0_i_4 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(pc[12]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(sp_reg[12]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_9_n_0 ),
        .O(\addr[12]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00002020000A202A)) 
    \addr[12]_INST_0_i_5 
       (.I0(\sr_reg_n_0_[12] ),
        .I1(din[4]),
        .I2(p_2_in88_in),
        .I3(r_code[4]),
        .I4(din[5]),
        .I5(r_code[5]),
        .O(\addr[12]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000505030000000)) 
    \addr[12]_INST_0_i_6 
       (.I0(r_code[3]),
        .I1(din[3]),
        .I2(\addr[12]_INST_0_i_11_n_0 ),
        .I3(din[2]),
        .I4(p_2_in88_in),
        .I5(r_code[2]),
        .O(\addr[12]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[12]_INST_0_i_7 
       (.I0(\addr[12]_INST_0_i_12_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[12]),
        .I3(state[0]),
        .I4(plusOp4_out[12]),
        .O(\addr[12]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAACCAACCF0FFF000)) 
    \addr[12]_INST_0_i_8 
       (.I0(\addr[12]_INST_0_i_13_n_0 ),
        .I1(\addr[12]_INST_0_i_14_n_0 ),
        .I2(\addr[12]_INST_0_i_15_n_0 ),
        .I3(\r_code[10]_i_1_n_0 ),
        .I4(\addr[12]_INST_0_i_16_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\addr[12]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[12]_INST_0_i_9 
       (.I0(\r_reg[11] [12]),
        .I1(\r_reg[10] [12]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [12]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [12]),
        .O(\addr[12]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4F44)) 
    \addr[13]_INST_0 
       (.I0(\addr[15]_INST_0_i_1_n_0 ),
        .I1(\rrs[0] [13]),
        .I2(\addr[15]_INST_0_i_3_n_0 ),
        .I3(sp_reg[13]),
        .I4(\addr[13]_INST_0_i_2_n_0 ),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(addr[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEFEEEEEE)) 
    \addr[13]_INST_0_i_1 
       (.I0(\addr[13]_INST_0_i_3_n_0 ),
        .I1(\addr[13]_INST_0_i_4_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\addr[13]_INST_0_i_5_n_0 ),
        .I4(\addr[14]_INST_0_i_5_n_0 ),
        .I5(\addr[13]_INST_0_i_6_n_0 ),
        .O(\rrs[0] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[13]_INST_0_i_10 
       (.I0(\r_reg[15] [13]),
        .I1(\r_reg[14] [13]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [13]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [13]),
        .O(\addr[13]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[13]_INST_0_i_11 
       (.I0(\r_reg[7] [13]),
        .I1(\r_reg[6] [13]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [13]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [13]),
        .O(\addr[13]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[13]_INST_0_i_12 
       (.I0(\addr[15]_INST_0_i_38_n_6 ),
        .I1(p_4_in),
        .I2(pc[13]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[13]),
        .O(\addr[13]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[13]_INST_0_i_13 
       (.I0(\r_reg[15] [13]),
        .I1(\r_reg[14] [13]),
        .I2(soc[2]),
        .I3(\r_reg[13] [13]),
        .I4(soc[1]),
        .I5(\r_reg[12] [13]),
        .O(\addr[13]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[13]_INST_0_i_14 
       (.I0(\r_reg[11] [13]),
        .I1(\r_reg[10] [13]),
        .I2(soc[2]),
        .I3(\r_reg[9] [13]),
        .I4(soc[1]),
        .I5(\r_reg[8] [13]),
        .O(\addr[13]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5F50CFCF5F50C0C0)) 
    \addr[13]_INST_0_i_15 
       (.I0(\addr[15]_INST_0_i_20_n_0 ),
        .I1(\addr[13]_INST_0_i_5_n_0 ),
        .I2(soc[2]),
        .I3(sp_reg[13]),
        .I4(soc[1]),
        .I5(pc[13]),
        .O(\addr[13]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[13]_INST_0_i_16 
       (.I0(\r_reg[7] [13]),
        .I1(\r_reg[6] [13]),
        .I2(soc[2]),
        .I3(\r_reg[5] [13]),
        .I4(soc[1]),
        .I5(\r_reg[4] [13]),
        .O(\addr[13]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000FFB8B8)) 
    \addr[13]_INST_0_i_2 
       (.I0(data3[13]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[13]_INST_0_i_7_n_0 ),
        .I3(\addr[13]_INST_0_i_8_n_0 ),
        .I4(\addr[15]_INST_0_i_17_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[13]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEA202A00000000)) 
    \addr[13]_INST_0_i_3 
       (.I0(\addr[13]_INST_0_i_9_n_0 ),
        .I1(din[2]),
        .I2(p_2_in88_in),
        .I3(r_code[2]),
        .I4(\addr[13]_INST_0_i_10_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\addr[13]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA0000A808)) 
    \addr[13]_INST_0_i_4 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(pc[13]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(sp_reg[13]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_9_n_0 ),
        .O(\addr[13]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00002020000A202A)) 
    \addr[13]_INST_0_i_5 
       (.I0(\sr_reg_n_0_[13] ),
        .I1(din[4]),
        .I2(p_2_in88_in),
        .I3(r_code[4]),
        .I4(din[5]),
        .I5(r_code[5]),
        .O(\addr[13]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000505030000000)) 
    \addr[13]_INST_0_i_6 
       (.I0(r_code[3]),
        .I1(din[3]),
        .I2(\addr[13]_INST_0_i_11_n_0 ),
        .I3(din[2]),
        .I4(p_2_in88_in),
        .I5(r_code[2]),
        .O(\addr[13]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[13]_INST_0_i_7 
       (.I0(\addr[13]_INST_0_i_12_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[13]),
        .I3(state[0]),
        .I4(plusOp4_out[13]),
        .O(\addr[13]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAACCCCFF000F0F)) 
    \addr[13]_INST_0_i_8 
       (.I0(\addr[13]_INST_0_i_13_n_0 ),
        .I1(\addr[13]_INST_0_i_14_n_0 ),
        .I2(\addr[13]_INST_0_i_15_n_0 ),
        .I3(\addr[13]_INST_0_i_16_n_0 ),
        .I4(\r_code[10]_i_1_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\addr[13]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[13]_INST_0_i_9 
       (.I0(\r_reg[11] [13]),
        .I1(\r_reg[10] [13]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [13]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [13]),
        .O(\addr[13]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1F11)) 
    \addr[14]_INST_0 
       (.I0(\addr[15]_INST_0_i_1_n_0 ),
        .I1(\addr[14]_INST_0_i_1_n_0 ),
        .I2(\addr[15]_INST_0_i_3_n_0 ),
        .I3(sp_reg[14]),
        .I4(\addr[14]_INST_0_i_2_n_0 ),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(addr[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000FF8A)) 
    \addr[14]_INST_0_i_1 
       (.I0(\addr[14]_INST_0_i_3_n_0 ),
        .I1(\addr[14]_INST_0_i_4_n_0 ),
        .I2(\addr[14]_INST_0_i_5_n_0 ),
        .I3(\r_code[3]_i_1_n_0 ),
        .I4(\addr[14]_INST_0_i_6_n_0 ),
        .I5(\addr[14]_INST_0_i_7_n_0 ),
        .O(\addr[14]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[14]_INST_0_i_10 
       (.I0(\r_reg[7] [14]),
        .I1(\r_reg[6] [14]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [14]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [14]),
        .O(\addr[14]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[14]_INST_0_i_11 
       (.I0(\r_reg[11] [14]),
        .I1(\r_reg[10] [14]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [14]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [14]),
        .O(\addr[14]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[14]_INST_0_i_12 
       (.I0(\r_reg[15] [14]),
        .I1(\r_reg[14] [14]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [14]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [14]),
        .O(\addr[14]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[14]_INST_0_i_13 
       (.I0(\addr[15]_INST_0_i_38_n_5 ),
        .I1(p_4_in),
        .I2(pc[14]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[14]),
        .O(\addr[14]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \addr[14]_INST_0_i_14 
       (.I0(\addr[14]_INST_0_i_16_n_0 ),
        .I1(\addr[14]_INST_0_i_17_n_0 ),
        .O(\addr[14]_INST_0_i_14_n_0 ),
        .S(\r_code[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \addr[14]_INST_0_i_15 
       (.I0(\addr[14]_INST_0_i_18_n_0 ),
        .I1(\addr[14]_INST_0_i_19_n_0 ),
        .O(\addr[14]_INST_0_i_15_n_0 ),
        .S(\r_code[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5F503F3F5F503030)) 
    \addr[14]_INST_0_i_16 
       (.I0(\addr[15]_INST_0_i_20_n_0 ),
        .I1(\addr[14]_INST_0_i_4_n_0 ),
        .I2(soc[2]),
        .I3(sp_reg[14]),
        .I4(soc[1]),
        .I5(pc[14]),
        .O(\addr[14]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[14]_INST_0_i_17 
       (.I0(\r_reg[7] [14]),
        .I1(\r_reg[6] [14]),
        .I2(soc[2]),
        .I3(\r_reg[5] [14]),
        .I4(soc[1]),
        .I5(\r_reg[4] [14]),
        .O(\addr[14]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[14]_INST_0_i_18 
       (.I0(\r_reg[11] [14]),
        .I1(\r_reg[10] [14]),
        .I2(soc[2]),
        .I3(\r_reg[9] [14]),
        .I4(soc[1]),
        .I5(\r_reg[8] [14]),
        .O(\addr[14]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[14]_INST_0_i_19 
       (.I0(\r_reg[15] [14]),
        .I1(\r_reg[14] [14]),
        .I2(soc[2]),
        .I3(\r_reg[13] [14]),
        .I4(soc[1]),
        .I5(\r_reg[12] [14]),
        .O(\addr[14]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    \addr[14]_INST_0_i_2 
       (.I0(data3[14]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[14]_INST_0_i_8_n_0 ),
        .I3(\addr[15]_INST_0_i_17_n_0 ),
        .I4(\addr[14]_INST_0_i_9_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[14]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    \addr[14]_INST_0_i_3 
       (.I0(r_code[2]),
        .I1(p_2_in88_in),
        .I2(din[2]),
        .I3(\addr[14]_INST_0_i_10_n_0 ),
        .O(\addr[14]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFBBFCB8FFFFFFFF)) 
    \addr[14]_INST_0_i_4 
       (.I0(din[4]),
        .I1(p_2_in88_in),
        .I2(r_code[4]),
        .I3(din[5]),
        .I4(r_code[5]),
        .I5(\sr_reg_n_0_[14] ),
        .O(\addr[14]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000404005004540)) 
    \addr[14]_INST_0_i_5 
       (.I0(\r_code[0]_i_1_n_0 ),
        .I1(din[1]),
        .I2(p_2_in88_in),
        .I3(r_code[1]),
        .I4(din[2]),
        .I5(r_code[2]),
        .O(\addr[14]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA0000A808)) 
    \addr[14]_INST_0_i_6 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(pc[14]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(sp_reg[14]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_9_n_0 ),
        .O(\addr[14]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEA202A00000000)) 
    \addr[14]_INST_0_i_7 
       (.I0(\addr[14]_INST_0_i_11_n_0 ),
        .I1(din[2]),
        .I2(p_2_in88_in),
        .I3(r_code[2]),
        .I4(\addr[14]_INST_0_i_12_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\addr[14]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[14]_INST_0_i_8 
       (.I0(\addr[14]_INST_0_i_13_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[14]),
        .I3(state[0]),
        .I4(plusOp4_out[14]),
        .O(\addr[14]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \addr[14]_INST_0_i_9 
       (.I0(\addr[14]_INST_0_i_14_n_0 ),
        .I1(\addr[14]_INST_0_i_15_n_0 ),
        .O(\addr[14]_INST_0_i_9_n_0 ),
        .S(\r_code[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4F44)) 
    \addr[15]_INST_0 
       (.I0(\addr[15]_INST_0_i_1_n_0 ),
        .I1(\addr[15]_INST_0_i_2_n_0 ),
        .I2(\addr[15]_INST_0_i_3_n_0 ),
        .I3(sp_reg[15]),
        .I4(\addr[15]_INST_0_i_4_n_0 ),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(addr[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00019108FFFFFFFF)) 
    \addr[15]_INST_0_i_1 
       (.I0(state[2]),
        .I1(state[3]),
        .I2(state[0]),
        .I3(state[1]),
        .I4(state[4]),
        .I5(\addr[15]_INST_0_i_6_n_0 ),
        .O(\addr[15]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \addr[15]_INST_0_i_10 
       (.I0(pc[15]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(sp_reg[15]),
        .I3(\r_code[1]_i_1_n_0 ),
        .O(\addr[15]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00053305)) 
    \addr[15]_INST_0_i_11 
       (.I0(r_code[2]),
        .I1(din[2]),
        .I2(r_code[3]),
        .I3(p_2_in88_in),
        .I4(din[3]),
        .O(\addr[15]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFFF5D)) 
    \addr[15]_INST_0_i_12 
       (.I0(\r_code[3]_i_1_n_0 ),
        .I1(\r_reg[12] [15]),
        .I2(\addr[15]_INST_0_i_21_n_0 ),
        .I3(\addr[15]_INST_0_i_22_n_0 ),
        .I4(\addr[15]_INST_0_i_23_n_0 ),
        .I5(\addr[15]_INST_0_i_24_n_0 ),
        .O(\addr[15]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[15]_INST_0_i_13 
       (.CI(\addr[11]_INST_0_i_7_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,din[14:12]}),
        .O(data3[15:12]),
        .S({\addr[15]_INST_0_i_25_n_0 ,\addr[15]_INST_0_i_26_n_0 ,\addr[15]_INST_0_i_27_n_0 ,\addr[15]_INST_0_i_28_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000C200)) 
    \addr[15]_INST_0_i_14 
       (.I0(eqOp113_in),
        .I1(state[1]),
        .I2(state[0]),
        .I3(state[2]),
        .I4(state[4]),
        .I5(state[3]),
        .O(\addr[15]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[15]_INST_0_i_15 
       (.I0(\addr[15]_INST_0_i_30_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[15]),
        .I3(state[0]),
        .I4(plusOp4_out[15]),
        .O(\addr[15]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \addr[15]_INST_0_i_16 
       (.I0(\addr[15]_INST_0_i_34_n_0 ),
        .I1(\addr[15]_INST_0_i_35_n_0 ),
        .O(\addr[15]_INST_0_i_16_n_0 ),
        .S(\r_code[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FB0000000000)) 
    \addr[15]_INST_0_i_17 
       (.I0(\r_code[11]_i_1_n_0 ),
        .I1(soc[2]),
        .I2(\r_code[10]_i_1_n_0 ),
        .I3(as[1]),
        .I4(\dout[13]_INST_0_i_3_n_0 ),
        .I5(p_2_in88_in),
        .O(\addr[15]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABEBABAAEA)) 
    \addr[15]_INST_0_i_18 
       (.I0(\addr[15]_INST_0_i_6_n_0 ),
        .I1(state[2]),
        .I2(state[3]),
        .I3(state[0]),
        .I4(state[1]),
        .I5(state[4]),
        .O(\addr[15]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFED)) 
    \addr[15]_INST_0_i_19 
       (.I0(state[3]),
        .I1(state[4]),
        .I2(state[2]),
        .I3(state[0]),
        .I4(state[1]),
        .O(\addr[15]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF10000)) 
    \addr[15]_INST_0_i_2 
       (.I0(\addr[15]_INST_0_i_7_n_0 ),
        .I1(\addr[15]_INST_0_i_8_n_0 ),
        .I2(\addr[15]_INST_0_i_9_n_0 ),
        .I3(\addr[15]_INST_0_i_10_n_0 ),
        .I4(\addr[15]_INST_0_i_11_n_0 ),
        .I5(\addr[15]_INST_0_i_12_n_0 ),
        .O(\addr[15]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h335FFF5F)) 
    \addr[15]_INST_0_i_20 
       (.I0(r_code[5]),
        .I1(din[5]),
        .I2(r_code[4]),
        .I3(p_2_in88_in),
        .I4(din[4]),
        .O(\addr[15]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFBFBFFAFFBABF)) 
    \addr[15]_INST_0_i_21 
       (.I0(\r_code[0]_i_1_n_0 ),
        .I1(din[2]),
        .I2(p_2_in88_in),
        .I3(r_code[2]),
        .I4(din[1]),
        .I5(r_code[1]),
        .O(\addr[15]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AF00C000A000C0)) 
    \addr[15]_INST_0_i_22 
       (.I0(\r_reg[9] [15]),
        .I1(\r_reg[8] [15]),
        .I2(\addr[3]_INST_0_i_9_n_0 ),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[13] [15]),
        .O(\addr[15]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAF00AC00A000AC00)) 
    \addr[15]_INST_0_i_23 
       (.I0(\addr[15]_INST_0_i_36_n_0 ),
        .I1(\r_reg[14] [15]),
        .I2(\addr[3]_INST_0_i_9_n_0 ),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[15] [15]),
        .O(\addr[15]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000FFF7)) 
    \addr[15]_INST_0_i_24 
       (.I0(\r_reg[5] [15]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_9_n_0 ),
        .I4(\r_code[3]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_37_n_0 ),
        .O(\addr[15]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[15]_INST_0_i_25 
       (.I0(din[15]),
        .I1(\addr[15]_INST_0_i_2_n_0 ),
        .O(\addr[15]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[15]_INST_0_i_26 
       (.I0(din[14]),
        .I1(\addr[14]_INST_0_i_1_n_0 ),
        .O(\addr[15]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[15]_INST_0_i_27 
       (.I0(din[13]),
        .I1(\rrs[0] [13]),
        .O(\addr[15]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h36)) 
    \addr[15]_INST_0_i_28_rewire 
       (.I0(\addr[12]_INST_0_i_4_n_0 ),
        .I1(din[12]),
        .I2(\rrs[0] [12]),
        .O(\addr[15]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h040C0C0C)) 
    \addr[15]_INST_0_i_29 
       (.I0(\r_code[0]_i_1_n_0 ),
        .I1(as[0]),
        .I2(as[1]),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(\addr[15]_INST_0_i_11_n_0 ),
        .O(eqOp113_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBEFFFFB9)) 
    \addr[15]_INST_0_i_3 
       (.I0(state[4]),
        .I1(state[1]),
        .I2(state[0]),
        .I3(state[3]),
        .I4(state[2]),
        .O(\addr[15]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[15]_INST_0_i_30 
       (.I0(\addr[15]_INST_0_i_38_n_4 ),
        .I1(p_4_in),
        .I2(pc[15]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[15]),
        .O(\addr[15]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFDFDFF)) 
    \addr[15]_INST_0_i_31 
       (.I0(state[3]),
        .I1(state[4]),
        .I2(state[2]),
        .I3(state[1]),
        .I4(state[0]),
        .O(\addr[15]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[15]_INST_0_i_32 
       (.CI(\addr[11]_INST_0_i_18_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,din[14:12]}),
        .O(plusOp3_out[15:12]),
        .S({\addr[15]_INST_0_i_42_n_0 ,\addr[15]_INST_0_i_43_n_0 ,\addr[15]_INST_0_i_44_n_0 ,\addr[15]_INST_0_i_45_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[15]_INST_0_i_33 
       (.CI(\addr[11]_INST_0_i_19_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,din[14:12]}),
        .O(plusOp4_out[15:12]),
        .S({\addr[15]_INST_0_i_46_n_0 ,\addr[15]_INST_0_i_47_n_0 ,\addr[15]_INST_0_i_48_n_0 ,\addr[15]_INST_0_i_49_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \addr[15]_INST_0_i_34 
       (.I0(\addr[15]_INST_0_i_50_n_0 ),
        .I1(\addr[15]_INST_0_i_51_n_0 ),
        .O(\addr[15]_INST_0_i_34_n_0 ),
        .S(\r_code[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \addr[15]_INST_0_i_35 
       (.I0(\addr[15]_INST_0_i_52_n_0 ),
        .I1(\addr[15]_INST_0_i_53_n_0 ),
        .O(\addr[15]_INST_0_i_35_n_0 ),
        .S(\r_code[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \addr[15]_INST_0_i_36 
       (.I0(\r_reg[11] [15]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\r_reg[10] [15]),
        .O(\addr[15]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00A000FC00A0000C)) 
    \addr[15]_INST_0_i_37 
       (.I0(\r_reg[7] [15]),
        .I1(\r_reg[4] [15]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_9_n_0 ),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[6] [15]),
        .O(\addr[15]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[15]_INST_0_i_38 
       (.CI(\addr[11]_INST_0_i_24_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,bsaddr__0[14:12]}),
        .O({\addr[15]_INST_0_i_38_n_4 ,\addr[15]_INST_0_i_38_n_5 ,\addr[15]_INST_0_i_38_n_6 ,\addr[15]_INST_0_i_38_n_7 }),
        .S({\addr[15]_INST_0_i_54_n_0 ,\addr[15]_INST_0_i_55_n_0 ,\addr[15]_INST_0_i_56_n_0 ,\addr[15]_INST_0_i_57_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000080)) 
    \addr[15]_INST_0_i_39 
       (.I0(state[2]),
        .I1(state[1]),
        .I2(state[3]),
        .I3(state[4]),
        .I4(state[0]),
        .O(p_4_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000FFB8B8)) 
    \addr[15]_INST_0_i_4 
       (.I0(data3[15]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[15]_INST_0_i_15_n_0 ),
        .I3(\addr[15]_INST_0_i_16_n_0 ),
        .I4(\addr[15]_INST_0_i_17_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[15]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEFFFFFFFFF)) 
    \addr[15]_INST_0_i_40 
       (.I0(state[2]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[0]),
        .I4(state[1]),
        .I5(eqOp113_in),
        .O(\addr[15]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[15]_INST_0_i_41 
       (.CI(\addr[11]_INST_0_i_25_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,bsaddr__0[14:12]}),
        .O(plusOp2_out[15:12]),
        .S({\addr[15]_INST_0_i_58_n_0 ,\addr[15]_INST_0_i_59_n_0 ,\addr[15]_INST_0_i_60_n_0 ,\addr[15]_INST_0_i_61_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[15]_INST_0_i_42 
       (.I0(din[15]),
        .I1(\addr[15]_INST_0_i_62_n_0 ),
        .O(\addr[15]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[15]_INST_0_i_43 
       (.I0(din[14]),
        .I1(\rrd[0] [14]),
        .O(\addr[15]_INST_0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[15]_INST_0_i_44 
       (.I0(din[13]),
        .I1(\rrd[0] [13]),
        .O(\addr[15]_INST_0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[15]_INST_0_i_45 
       (.I0(din[12]),
        .I1(\rrd[0] [12]),
        .O(\addr[15]_INST_0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[15]_INST_0_i_46 
       (.I0(din[15]),
        .I1(\addr[15]_INST_0_i_16_n_0 ),
        .O(\addr[15]_INST_0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[15]_INST_0_i_47 
       (.I0(din[14]),
        .I1(\addr[14]_INST_0_i_9_n_0 ),
        .O(\addr[15]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[15]_INST_0_i_48 
       (.I0(din[13]),
        .I1(\addr[13]_INST_0_i_8_n_0 ),
        .O(\addr[15]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[15]_INST_0_i_49 
       (.I0(din[12]),
        .I1(\addr[12]_INST_0_i_8_n_0 ),
        .O(\addr[15]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00100000)) 
    \addr[15]_INST_0_i_5 
       (.I0(state[1]),
        .I1(state[3]),
        .I2(state[4]),
        .I3(state[2]),
        .I4(state[0]),
        .O(\addr[15]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A0C0CFAFAFC0CF)) 
    \addr[15]_INST_0_i_50 
       (.I0(\addr[15]_INST_0_i_20_n_0 ),
        .I1(\addr[15]_INST_0_i_7_n_0 ),
        .I2(soc[2]),
        .I3(pc[15]),
        .I4(soc[1]),
        .I5(sp_reg[15]),
        .O(\addr[15]_INST_0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[15]_INST_0_i_51 
       (.I0(\r_reg[7] [15]),
        .I1(\r_reg[6] [15]),
        .I2(soc[2]),
        .I3(\r_reg[5] [15]),
        .I4(soc[1]),
        .I5(\r_reg[4] [15]),
        .O(\addr[15]_INST_0_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[15]_INST_0_i_52 
       (.I0(\r_reg[11] [15]),
        .I1(\r_reg[10] [15]),
        .I2(soc[2]),
        .I3(\r_reg[9] [15]),
        .I4(soc[1]),
        .I5(\r_reg[8] [15]),
        .O(\addr[15]_INST_0_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[15]_INST_0_i_53 
       (.I0(\r_reg[15] [15]),
        .I1(\r_reg[14] [15]),
        .I2(soc[2]),
        .I3(\r_reg[13] [15]),
        .I4(soc[1]),
        .I5(\r_reg[12] [15]),
        .O(\addr[15]_INST_0_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[15]_INST_0_i_54 
       (.I0(bsaddr__0[15]),
        .I1(\addr[15]_INST_0_i_16_n_0 ),
        .O(\addr[15]_INST_0_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[15]_INST_0_i_55 
       (.I0(bsaddr__0[14]),
        .I1(\addr[14]_INST_0_i_9_n_0 ),
        .O(\addr[15]_INST_0_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[15]_INST_0_i_56 
       (.I0(bsaddr__0[13]),
        .I1(\addr[13]_INST_0_i_8_n_0 ),
        .O(\addr[15]_INST_0_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[15]_INST_0_i_57 
       (.I0(bsaddr__0[12]),
        .I1(\addr[12]_INST_0_i_8_n_0 ),
        .O(\addr[15]_INST_0_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[15]_INST_0_i_58 
       (.I0(bsaddr__0[15]),
        .I1(\addr[15]_INST_0_i_2_n_0 ),
        .O(\addr[15]_INST_0_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[15]_INST_0_i_59 
       (.I0(bsaddr__0[14]),
        .I1(\addr[14]_INST_0_i_1_n_0 ),
        .O(\addr[15]_INST_0_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7000000070707070)) 
    \addr[15]_INST_0_i_6 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(\r_code[1]_i_1_n_0 ),
        .I2(as[1]),
        .I3(eqOp135_in),
        .I4(p_2_in88_in),
        .I5(\addr[15]_INST_0_i_19_n_0 ),
        .O(\addr[15]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[15]_INST_0_i_60 
       (.I0(bsaddr__0[13]),
        .I1(\rrs[0] [13]),
        .O(\addr[15]_INST_0_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h36)) 
    \addr[15]_INST_0_i_61_rewire 
       (.I0(\addr[12]_INST_0_i_4_n_0 ),
        .I1(bsaddr__0[12]),
        .I2(\rrs[0] [12]),
        .O(\addr[15]_INST_0_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFEEEAAAA)) 
    \addr[15]_INST_0_i_62 
       (.I0(\addr[15]_INST_0_i_12_n_0 ),
        .I1(\addr[15]_INST_0_i_10_n_0 ),
        .I2(\addr[3]_INST_0_i_47_n_0 ),
        .I3(\sr_reg_n_0_[15] ),
        .I4(\addr[15]_INST_0_i_11_n_0 ),
        .O(\addr[15]_INST_0_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEEAAA)) 
    \addr[15]_INST_0_i_63 
       (.I0(\addr[13]_INST_0_i_3_n_0 ),
        .I1(\addr[15]_INST_0_i_11_n_0 ),
        .I2(\sr_reg_n_0_[13] ),
        .I3(\addr[3]_INST_0_i_47_n_0 ),
        .I4(\addr[15]_INST_0_i_65_n_0 ),
        .I5(\addr[13]_INST_0_i_6_n_0 ),
        .O(\rrd[0] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEEAAA)) 
    \addr[15]_INST_0_i_64 
       (.I0(\addr[12]_INST_0_i_3_n_0 ),
        .I1(\addr[15]_INST_0_i_11_n_0 ),
        .I2(\sr_reg_n_0_[12] ),
        .I3(\addr[3]_INST_0_i_47_n_0 ),
        .I4(\addr[15]_INST_0_i_66_n_0 ),
        .I5(\addr[12]_INST_0_i_6_n_0 ),
        .O(\rrd[0] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \addr[15]_INST_0_i_65 
       (.I0(pc[13]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(sp_reg[13]),
        .I3(\r_code[1]_i_1_n_0 ),
        .O(\addr[15]_INST_0_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \addr[15]_INST_0_i_66 
       (.I0(pc[12]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(sp_reg[12]),
        .I3(\r_code[1]_i_1_n_0 ),
        .O(\addr[15]_INST_0_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFBBFCB8FFFFFFFF)) 
    \addr[15]_INST_0_i_7 
       (.I0(din[4]),
        .I1(p_2_in88_in),
        .I2(r_code[4]),
        .I3(din[5]),
        .I4(r_code[5]),
        .I5(\sr_reg_n_0_[15] ),
        .O(\addr[15]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \addr[15]_INST_0_i_8 
       (.I0(\r_code[0]_i_1_n_0 ),
        .I1(\r_code[1]_i_1_n_0 ),
        .O(\addr[15]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \addr[15]_INST_0_i_9 
       (.I0(\r_code[1]_i_1_n_0 ),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\addr[15]_INST_0_i_20_n_0 ),
        .O(\addr[15]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8BBB8BBBBBBB8)) 
    \addr[1]_INST_0 
       (.I0(irqaddr[1]),
        .I1(\addr[15]_INST_0_i_5_n_0 ),
        .I2(\addr[1]_INST_0_i_1_n_0 ),
        .I3(\addr[1]_INST_0_i_2_n_0 ),
        .I4(\rrs[0] [1]),
        .I5(\addr[15]_INST_0_i_1_n_0 ),
        .O(addr[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    \addr[1]_INST_0_i_1 
       (.I0(data3[1]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[1]_INST_0_i_4_n_0 ),
        .I3(\addr[15]_INST_0_i_17_n_0 ),
        .I4(\addr[1]_INST_0_i_5_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0F0C000A000C000)) 
    \addr[1]_INST_0_i_10 
       (.I0(\r_reg[11] [1]),
        .I1(\r_reg[10] [1]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_9_n_0 ),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[15] [1]),
        .O(\addr[1]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h1000FFFF)) 
    \addr[1]_INST_0_i_11 
       (.I0(\addr[3]_INST_0_i_9_n_0 ),
        .I1(\r_code[1]_i_1_n_0 ),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(\r_reg[13] [1]),
        .I4(\r_code[3]_i_1_n_0 ),
        .O(\addr[1]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[1]_INST_0_i_12 
       (.I0(\addr[3]_INST_0_i_23_n_6 ),
        .I1(p_4_in),
        .I2(pc[1]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[1]),
        .O(\addr[1]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[1]_INST_0_i_13 
       (.I0(\r_reg[15] [1]),
        .I1(\r_reg[14] [1]),
        .I2(soc[2]),
        .I3(\r_reg[13] [1]),
        .I4(soc[1]),
        .I5(\r_reg[12] [1]),
        .O(\addr[1]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[1]_INST_0_i_14 
       (.I0(\r_reg[11] [1]),
        .I1(\r_reg[10] [1]),
        .I2(soc[2]),
        .I3(\r_reg[9] [1]),
        .I4(soc[1]),
        .I5(\r_reg[8] [1]),
        .O(\addr[1]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505FC0C0505FCFCF)) 
    \addr[1]_INST_0_i_15 
       (.I0(as[1]),
        .I1(\addr[1]_INST_0_i_18_n_0 ),
        .I2(soc[2]),
        .I3(sp_reg[1]),
        .I4(soc[1]),
        .I5(pc[1]),
        .O(\addr[1]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[1]_INST_0_i_16 
       (.I0(\r_reg[7] [1]),
        .I1(\r_reg[6] [1]),
        .I2(soc[2]),
        .I3(\r_reg[5] [1]),
        .I4(soc[1]),
        .I5(\r_reg[4] [1]),
        .O(\addr[1]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBABF8A80)) 
    \addr[1]_INST_0_i_17 
       (.I0(sp_reg[1]),
        .I1(din[0]),
        .I2(p_2_in88_in),
        .I3(r_code[0]),
        .I4(pc[1]),
        .O(\addr[1]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFBBFCB8FFFFFFFF)) 
    \addr[1]_INST_0_i_18 
       (.I0(din[4]),
        .I1(p_2_in88_in),
        .I2(r_code[4]),
        .I3(din[5]),
        .I4(r_code[5]),
        .I5(\sr_reg_n_0_[1] ),
        .O(\addr[1]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBABF8A80)) 
    \addr[1]_INST_0_i_19 
       (.I0(\r_reg[9] [1]),
        .I1(din[0]),
        .I2(p_2_in88_in),
        .I3(r_code[0]),
        .I4(\r_reg[8] [1]),
        .O(\addr[1]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000282020080)) 
    \addr[1]_INST_0_i_2 
       (.I0(sp_reg[1]),
        .I1(state[2]),
        .I2(state[3]),
        .I3(state[0]),
        .I4(state[1]),
        .I5(state[4]),
        .O(\addr[1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBFBFBFBFBFBFBAA)) 
    \addr[1]_INST_0_i_3 
       (.I0(\addr[1]_INST_0_i_6_n_0 ),
        .I1(\addr[1]_INST_0_i_7_n_0 ),
        .I2(\addr[1]_INST_0_i_8_n_0 ),
        .I3(\addr[1]_INST_0_i_9_n_0 ),
        .I4(\addr[1]_INST_0_i_10_n_0 ),
        .I5(\addr[1]_INST_0_i_11_n_0 ),
        .O(\rrs[0] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[1]_INST_0_i_4 
       (.I0(\addr[1]_INST_0_i_12_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[1]),
        .I3(state[0]),
        .I4(plusOp4_out[1]),
        .O(\addr[1]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFAFC0CFA0A0C0CF)) 
    \addr[1]_INST_0_i_5 
       (.I0(\addr[1]_INST_0_i_13_n_0 ),
        .I1(\addr[1]_INST_0_i_14_n_0 ),
        .I2(\r_code[11]_i_1_n_0 ),
        .I3(\addr[1]_INST_0_i_15_n_0 ),
        .I4(\r_code[10]_i_1_n_0 ),
        .I5(\addr[1]_INST_0_i_16_n_0 ),
        .O(\addr[1]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0880088AA880A88)) 
    \addr[1]_INST_0_i_6 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(\addr[1]_INST_0_i_17_n_0 ),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(as[1]),
        .I5(\addr[1]_INST_0_i_18_n_0 ),
        .O(\addr[1]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h54555555)) 
    \addr[1]_INST_0_i_7 
       (.I0(\r_code[3]_i_1_n_0 ),
        .I1(\addr[3]_INST_0_i_9_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_code[0]_i_1_n_0 ),
        .I4(\r_reg[5] [1]),
        .O(\addr[1]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00A000FC00A0000C)) 
    \addr[1]_INST_0_i_8 
       (.I0(\r_reg[7] [1]),
        .I1(\r_reg[4] [1]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_9_n_0 ),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[6] [1]),
        .O(\addr[1]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F000FAC000000AC)) 
    \addr[1]_INST_0_i_9 
       (.I0(\r_reg[14] [1]),
        .I1(\r_reg[12] [1]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_9_n_0 ),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\addr[1]_INST_0_i_19_n_0 ),
        .O(\addr[1]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8BBB8BBBBBBB8)) 
    \addr[2]_INST_0 
       (.I0(irqaddr[2]),
        .I1(\addr[15]_INST_0_i_5_n_0 ),
        .I2(\addr[2]_INST_0_i_1_n_0 ),
        .I3(\addr[2]_INST_0_i_2_n_0 ),
        .I4(\rrs[0] [2]),
        .I5(\addr[15]_INST_0_i_1_n_0 ),
        .O(addr[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000FFB8B8)) 
    \addr[2]_INST_0_i_1 
       (.I0(data3[2]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[2]_INST_0_i_4_n_0 ),
        .I3(\addr[2]_INST_0_i_5_n_0 ),
        .I4(\addr[15]_INST_0_i_17_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[2]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[2]_INST_0_i_10 
       (.I0(\addr[3]_INST_0_i_23_n_5 ),
        .I1(p_4_in),
        .I2(pc[2]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[2]),
        .O(\addr[2]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[2]_INST_0_i_11 
       (.I0(\r_reg[15] [2]),
        .I1(\r_reg[14] [2]),
        .I2(soc[2]),
        .I3(\r_reg[13] [2]),
        .I4(soc[1]),
        .I5(\r_reg[12] [2]),
        .O(\addr[2]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[2]_INST_0_i_12 
       (.I0(\r_reg[11] [2]),
        .I1(\r_reg[10] [2]),
        .I2(soc[2]),
        .I3(\r_reg[9] [2]),
        .I4(soc[1]),
        .I5(\r_reg[8] [2]),
        .O(\addr[2]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[2]_INST_0_i_13 
       (.I0(\r_reg[7] [2]),
        .I1(\r_reg[6] [2]),
        .I2(soc[2]),
        .I3(\r_reg[5] [2]),
        .I4(soc[1]),
        .I5(\r_reg[4] [2]),
        .O(\addr[2]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF000F0FF55335533)) 
    \addr[2]_INST_0_i_14 
       (.I0(sp_reg[2]),
        .I1(pc[2]),
        .I2(\addr[15]_INST_0_i_20_n_0 ),
        .I3(soc[1]),
        .I4(\addr[2]_INST_0_i_8_n_0 ),
        .I5(soc[2]),
        .O(\addr[2]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBABF8A80)) 
    \addr[2]_INST_0_i_15 
       (.I0(\r_reg[15] [2]),
        .I1(din[0]),
        .I2(p_2_in88_in),
        .I3(r_code[0]),
        .I4(\r_reg[14] [2]),
        .O(\addr[2]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBABF8A80)) 
    \addr[2]_INST_0_i_16 
       (.I0(\r_reg[13] [2]),
        .I1(din[0]),
        .I2(p_2_in88_in),
        .I3(r_code[0]),
        .I4(\r_reg[12] [2]),
        .O(\addr[2]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBABF8A80)) 
    \addr[2]_INST_0_i_17 
       (.I0(\r_reg[11] [2]),
        .I1(din[0]),
        .I2(p_2_in88_in),
        .I3(r_code[0]),
        .I4(\r_reg[10] [2]),
        .O(\addr[2]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBABF8A80)) 
    \addr[2]_INST_0_i_18 
       (.I0(\r_reg[9] [2]),
        .I1(din[0]),
        .I2(p_2_in88_in),
        .I3(r_code[0]),
        .I4(\r_reg[8] [2]),
        .O(\addr[2]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBABF8A80)) 
    \addr[2]_INST_0_i_19 
       (.I0(\r_reg[7] [2]),
        .I1(din[0]),
        .I2(p_2_in88_in),
        .I3(r_code[0]),
        .I4(\r_reg[6] [2]),
        .O(\addr[2]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000282020080)) 
    \addr[2]_INST_0_i_2 
       (.I0(sp_reg[2]),
        .I1(state[2]),
        .I2(state[3]),
        .I3(state[0]),
        .I4(state[1]),
        .I5(state[4]),
        .O(\addr[2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBABF8A80)) 
    \addr[2]_INST_0_i_20 
       (.I0(\r_reg[5] [2]),
        .I1(din[0]),
        .I2(p_2_in88_in),
        .I3(r_code[0]),
        .I4(\r_reg[4] [2]),
        .O(\addr[2]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEFECECEC)) 
    \addr[2]_INST_0_i_3 
       (.I0(\addr[2]_INST_0_i_6_n_0 ),
        .I1(\addr[2]_INST_0_i_7_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\addr[2]_INST_0_i_8_n_0 ),
        .I4(\addr[14]_INST_0_i_5_n_0 ),
        .I5(\addr[2]_INST_0_i_9_n_0 ),
        .O(\rrs[0] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[2]_INST_0_i_4 
       (.I0(\addr[2]_INST_0_i_10_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[2]),
        .I3(state[0]),
        .I4(plusOp4_out[2]),
        .O(\addr[2]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAACCAACCF0FFF000)) 
    \addr[2]_INST_0_i_5 
       (.I0(\addr[2]_INST_0_i_11_n_0 ),
        .I1(\addr[2]_INST_0_i_12_n_0 ),
        .I2(\addr[2]_INST_0_i_13_n_0 ),
        .I3(\r_code[10]_i_1_n_0 ),
        .I4(\addr[2]_INST_0_i_14_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\addr[2]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \addr[2]_INST_0_i_6 
       (.I0(\addr[2]_INST_0_i_15_n_0 ),
        .I1(\addr[2]_INST_0_i_16_n_0 ),
        .I2(\addr[3]_INST_0_i_9_n_0 ),
        .I3(\addr[2]_INST_0_i_17_n_0 ),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[2]_INST_0_i_18_n_0 ),
        .O(\addr[2]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000A808A0A0A808)) 
    \addr[2]_INST_0_i_7 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(pc[2]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(sp_reg[2]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_20_n_0 ),
        .O(\addr[2]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3355335530553000)) 
    \addr[2]_INST_0_i_8 
       (.I0(r_code[4]),
        .I1(din[4]),
        .I2(din[5]),
        .I3(p_2_in88_in),
        .I4(r_code[5]),
        .I5(p_1_in122_in),
        .O(\addr[2]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00004540)) 
    \addr[2]_INST_0_i_9 
       (.I0(\r_code[3]_i_1_n_0 ),
        .I1(\addr[2]_INST_0_i_19_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\addr[2]_INST_0_i_20_n_0 ),
        .I4(\addr[3]_INST_0_i_9_n_0 ),
        .O(\addr[2]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8BBB8BBBBBBB8)) 
    \addr[3]_INST_0 
       (.I0(irqaddr[3]),
        .I1(\addr[15]_INST_0_i_5_n_0 ),
        .I2(\addr[3]_INST_0_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_2_n_0 ),
        .I4(\rrs[0] [3]),
        .I5(\addr[15]_INST_0_i_1_n_0 ),
        .O(addr[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    \addr[3]_INST_0_i_1 
       (.I0(data3[3]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[3]_INST_0_i_5_n_0 ),
        .I3(\addr[15]_INST_0_i_17_n_0 ),
        .I4(\addr[3]_INST_0_i_6_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[3]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[3]_INST_0_i_10 
       (.I0(\r_reg[7] [3]),
        .I1(\r_reg[6] [3]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [3]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [3]),
        .O(\addr[3]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8988000000000000)) 
    \addr[3]_INST_0_i_11 
       (.I0(as[1]),
        .I1(as[0]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(p_1_in108_in),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[3]_INST_0_i_9_n_0 ),
        .O(\addr[3]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_12 
       (.I0(din[3]),
        .I1(\rrs[0] [3]),
        .O(\addr[3]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_13 
       (.I0(din[2]),
        .I1(\rrs[0] [2]),
        .O(\addr[3]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_14 
       (.I0(din[1]),
        .I1(\rrs[0] [1]),
        .O(\addr[3]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_15 
       (.I0(din[0]),
        .I1(\rrs[0] [0]),
        .O(\addr[3]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[3]_INST_0_i_16 
       (.I0(\addr[3]_INST_0_i_23_n_4 ),
        .I1(p_4_in),
        .I2(pc[3]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[3]),
        .O(\addr[3]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[3]_INST_0_i_17 
       (.CI(\<const0>__0__0 ),
        .CO({\addr[3]_INST_0_i_17_n_0 ,\addr[3]_INST_0_i_17_n_1 ,\addr[3]_INST_0_i_17_n_2 ,\addr[3]_INST_0_i_17_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(din[3:0]),
        .O(plusOp3_out[3:0]),
        .S({\addr[3]_INST_0_i_25_n_0 ,\addr[3]_INST_0_i_26_n_0 ,\addr[3]_INST_0_i_27_n_0 ,\addr[3]_INST_0_i_28_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[3]_INST_0_i_18 
       (.CI(\<const0>__0__0 ),
        .CO({\addr[3]_INST_0_i_18_n_0 ,\addr[3]_INST_0_i_18_n_1 ,\addr[3]_INST_0_i_18_n_2 ,\addr[3]_INST_0_i_18_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(din[3:0]),
        .O(plusOp4_out[3:0]),
        .S({\addr[3]_INST_0_i_29_n_0 ,\addr[3]_INST_0_i_30_n_0 ,\addr[3]_INST_0_i_31_n_0 ,\addr[3]_INST_0_i_32_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \addr[3]_INST_0_i_19 
       (.I0(\addr[3]_INST_0_i_33_n_0 ),
        .I1(\addr[3]_INST_0_i_34_n_0 ),
        .O(\addr[3]_INST_0_i_19_n_0 ),
        .S(\r_code[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000282020080)) 
    \addr[3]_INST_0_i_2 
       (.I0(sp_reg[3]),
        .I1(state[2]),
        .I2(state[3]),
        .I3(state[0]),
        .I4(state[1]),
        .I5(state[4]),
        .O(\addr[3]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \addr[3]_INST_0_i_20 
       (.I0(\addr[3]_INST_0_i_35_n_0 ),
        .I1(\addr[3]_INST_0_i_36_n_0 ),
        .O(\addr[3]_INST_0_i_20_n_0 ),
        .S(\r_code[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[3]_INST_0_i_21 
       (.I0(\r_reg[11] [3]),
        .I1(\r_reg[10] [3]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [3]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [3]),
        .O(\addr[3]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[3]_INST_0_i_22 
       (.I0(\r_reg[15] [3]),
        .I1(\r_reg[14] [3]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [3]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [3]),
        .O(\addr[3]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[3]_INST_0_i_23 
       (.CI(\<const0>__0__0 ),
        .CO({\addr[3]_INST_0_i_23_n_0 ,\addr[3]_INST_0_i_23_n_1 ,\addr[3]_INST_0_i_23_n_2 ,\addr[3]_INST_0_i_23_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(bsaddr__0[3:0]),
        .O({\addr[3]_INST_0_i_23_n_4 ,\addr[3]_INST_0_i_23_n_5 ,\addr[3]_INST_0_i_23_n_6 ,\addr[3]_INST_0_i_23_n_7 }),
        .S({\addr[3]_INST_0_i_37_n_0 ,\addr[3]_INST_0_i_38_n_0 ,\addr[3]_INST_0_i_39_n_0 ,\addr[3]_INST_0_i_40_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[3]_INST_0_i_24 
       (.CI(\<const0>__0__0 ),
        .CO({\addr[3]_INST_0_i_24_n_0 ,\addr[3]_INST_0_i_24_n_1 ,\addr[3]_INST_0_i_24_n_2 ,\addr[3]_INST_0_i_24_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(bsaddr__0[3:0]),
        .O(plusOp2_out[3:0]),
        .S({\addr[3]_INST_0_i_41_n_0 ,\addr[3]_INST_0_i_42_n_0 ,\addr[3]_INST_0_i_43_n_0 ,\addr[3]_INST_0_i_44_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_25 
       (.I0(din[3]),
        .I1(\rrd[0] [3]),
        .O(\addr[3]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_26 
       (.I0(din[2]),
        .I1(\rrd[0] [2]),
        .O(\addr[3]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555555566666AAA)) 
    \addr[3]_INST_0_i_27 
       (.I0(din[1]),
        .I1(\addr[15]_INST_0_i_11_n_0 ),
        .I2(\sr_reg_n_0_[1] ),
        .I3(\addr[3]_INST_0_i_47_n_0 ),
        .I4(\addr[3]_INST_0_i_48_n_0 ),
        .I5(\addr[3]_INST_0_i_49_n_0 ),
        .O(\addr[3]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h15EA)) 
    \addr[3]_INST_0_i_28 
       (.I0(lbe_INST_0_i_7_n_0),
        .I1(\addr[3]_INST_0_i_50_n_0 ),
        .I2(\addr[15]_INST_0_i_11_n_0 ),
        .I3(din[0]),
        .O(\addr[3]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_29 
       (.I0(din[3]),
        .I1(\addr[3]_INST_0_i_6_n_0 ),
        .O(\addr[3]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \addr[3]_INST_0_i_3 
       (.I0(\addr[3]_INST_0_i_7_n_0 ),
        .I1(\r_code[3]_i_1_n_0 ),
        .I2(\addr[3]_INST_0_i_8_n_0 ),
        .I3(\addr[3]_INST_0_i_9_n_0 ),
        .I4(\addr[3]_INST_0_i_10_n_0 ),
        .I5(\addr[3]_INST_0_i_11_n_0 ),
        .O(\rrs[0] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[3]_INST_0_i_30 
       (.I0(din[2]),
        .I1(\addr[2]_INST_0_i_5_n_0 ),
        .O(\addr[3]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_31 
       (.I0(din[1]),
        .I1(\addr[1]_INST_0_i_5_n_0 ),
        .O(\addr[3]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[3]_INST_0_i_32 
       (.I0(din[0]),
        .I1(lbe_INST_0_i_11_n_0),
        .O(\addr[3]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[3]_INST_0_i_33 
       (.I0(\addr[3]_INST_0_i_51_n_0 ),
        .I1(soc[2]),
        .I2(sp_reg[3]),
        .I3(soc[1]),
        .I4(pc[3]),
        .O(\addr[3]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[3]_INST_0_i_34 
       (.I0(\r_reg[7] [3]),
        .I1(\r_reg[6] [3]),
        .I2(soc[2]),
        .I3(\r_reg[5] [3]),
        .I4(soc[1]),
        .I5(\r_reg[4] [3]),
        .O(\addr[3]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[3]_INST_0_i_35 
       (.I0(\r_reg[11] [3]),
        .I1(\r_reg[10] [3]),
        .I2(soc[2]),
        .I3(\r_reg[9] [3]),
        .I4(soc[1]),
        .I5(\r_reg[8] [3]),
        .O(\addr[3]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[3]_INST_0_i_36 
       (.I0(\r_reg[15] [3]),
        .I1(\r_reg[14] [3]),
        .I2(soc[2]),
        .I3(\r_reg[13] [3]),
        .I4(soc[1]),
        .I5(\r_reg[12] [3]),
        .O(\addr[3]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_37 
       (.I0(bsaddr__0[3]),
        .I1(\addr[3]_INST_0_i_6_n_0 ),
        .O(\addr[3]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[3]_INST_0_i_38 
       (.I0(bsaddr__0[2]),
        .I1(\addr[2]_INST_0_i_5_n_0 ),
        .O(\addr[3]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_39 
       (.I0(bsaddr__0[1]),
        .I1(\addr[1]_INST_0_i_5_n_0 ),
        .O(\addr[3]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[3]_INST_0_i_4 
       (.CI(\<const0>__0__0 ),
        .CO({\addr[3]_INST_0_i_4_n_0 ,\addr[3]_INST_0_i_4_n_1 ,\addr[3]_INST_0_i_4_n_2 ,\addr[3]_INST_0_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(din[3:0]),
        .O(data3[3:0]),
        .S({\addr[3]_INST_0_i_12_n_0 ,\addr[3]_INST_0_i_13_n_0 ,\addr[3]_INST_0_i_14_n_0 ,\addr[3]_INST_0_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[3]_INST_0_i_40 
       (.I0(bsaddr__0[0]),
        .I1(lbe_INST_0_i_11_n_0),
        .O(\addr[3]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_41 
       (.I0(bsaddr__0[3]),
        .I1(\rrs[0] [3]),
        .O(\addr[3]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_42 
       (.I0(bsaddr__0[2]),
        .I1(\rrs[0] [2]),
        .O(\addr[3]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_43 
       (.I0(bsaddr__0[1]),
        .I1(\rrs[0] [1]),
        .O(\addr[3]_INST_0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[3]_INST_0_i_44 
       (.I0(bsaddr__0[0]),
        .I1(\rrs[0] [0]),
        .O(\addr[3]_INST_0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \addr[3]_INST_0_i_45 
       (.I0(\addr[3]_INST_0_i_22_n_0 ),
        .I1(\addr[3]_INST_0_i_21_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_52_n_0 ),
        .I4(\addr[3]_INST_0_i_9_n_0 ),
        .I5(\addr[3]_INST_0_i_10_n_0 ),
        .O(\rrd[0] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFAFC0AFCFA0C0A0)) 
    \addr[3]_INST_0_i_46 
       (.I0(\addr[3]_INST_0_i_53_n_0 ),
        .I1(\addr[3]_INST_0_i_54_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_9_n_0 ),
        .I4(\addr[3]_INST_0_i_55_n_0 ),
        .I5(\addr[3]_INST_0_i_56_n_0 ),
        .O(\rrd[0] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030553000)) 
    \addr[3]_INST_0_i_47 
       (.I0(r_code[7]),
        .I1(din[7]),
        .I2(din[1]),
        .I3(p_2_in88_in),
        .I4(r_code[1]),
        .I5(\r_code[0]_i_1_n_0 ),
        .O(\addr[3]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \addr[3]_INST_0_i_48 
       (.I0(pc[1]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(sp_reg[1]),
        .I3(\r_code[1]_i_1_n_0 ),
        .O(\addr[3]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFFFFFEFEFF00)) 
    \addr[3]_INST_0_i_49 
       (.I0(\addr[3]_INST_0_i_57_n_0 ),
        .I1(\addr[1]_INST_0_i_10_n_0 ),
        .I2(\addr[1]_INST_0_i_9_n_0 ),
        .I3(\addr[1]_INST_0_i_8_n_0 ),
        .I4(\r_code[3]_i_1_n_0 ),
        .I5(\addr[3]_INST_0_i_58_n_0 ),
        .O(\addr[3]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[3]_INST_0_i_5 
       (.I0(\addr[3]_INST_0_i_16_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[3]),
        .I3(state[0]),
        .I4(plusOp4_out[3]),
        .O(\addr[3]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC02F2FCFC02020)) 
    \addr[3]_INST_0_i_50 
       (.I0(sr_reg_n_0_),
        .I1(soc[0]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(sp_reg[0]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(pc[0]),
        .O(\addr[3]_INST_0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF002F0F0F0020202)) 
    \addr[3]_INST_0_i_51 
       (.I0(p_1_in108_in),
        .I1(soc[1]),
        .I2(as[0]),
        .I3(din[5]),
        .I4(p_2_in88_in),
        .I5(r_code[5]),
        .O(\addr[3]_INST_0_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AA0FCC00AA00CC)) 
    \addr[3]_INST_0_i_52 
       (.I0(sp_reg[3]),
        .I1(pc[3]),
        .I2(soc[0]),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(p_1_in108_in),
        .O(\addr[3]_INST_0_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[3]_INST_0_i_53 
       (.I0(\r_reg[15] [2]),
        .I1(\r_reg[14] [2]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [2]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [2]),
        .O(\addr[3]_INST_0_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[3]_INST_0_i_54 
       (.I0(\r_reg[11] [2]),
        .I1(\r_reg[10] [2]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [2]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [2]),
        .O(\addr[3]_INST_0_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000AAAA00F0CCCC)) 
    \addr[3]_INST_0_i_55 
       (.I0(sp_reg[2]),
        .I1(pc[2]),
        .I2(p_1_in122_in),
        .I3(soc[0]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\r_code[0]_i_1_n_0 ),
        .O(\addr[3]_INST_0_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[3]_INST_0_i_56 
       (.I0(\r_reg[7] [2]),
        .I1(\r_reg[6] [2]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [2]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [2]),
        .O(\addr[3]_INST_0_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0808080000000800)) 
    \addr[3]_INST_0_i_57 
       (.I0(\r_reg[13] [1]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(r_code[2]),
        .I4(p_2_in88_in),
        .I5(din[2]),
        .O(\addr[3]_INST_0_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0808080000000800)) 
    \addr[3]_INST_0_i_58 
       (.I0(\r_reg[5] [1]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(r_code[2]),
        .I4(p_2_in88_in),
        .I5(din[2]),
        .O(\addr[3]_INST_0_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \addr[3]_INST_0_i_6 
       (.I0(\addr[3]_INST_0_i_19_n_0 ),
        .I1(\addr[3]_INST_0_i_20_n_0 ),
        .O(\addr[3]_INST_0_i_6_n_0 ),
        .S(\r_code[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \addr[3]_INST_0_i_7 
       (.I0(\addr[3]_INST_0_i_21_n_0 ),
        .I1(\addr[3]_INST_0_i_22_n_0 ),
        .O(\addr[3]_INST_0_i_7_n_0 ),
        .S(\r_code[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \addr[3]_INST_0_i_8 
       (.I0(pc[3]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(sp_reg[3]),
        .I3(\r_code[1]_i_1_n_0 ),
        .O(\addr[3]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h47)) 
    \addr[3]_INST_0_i_9 
       (.I0(din[2]),
        .I1(p_2_in88_in),
        .I2(r_code[2]),
        .O(\addr[3]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "addr[3]_INST_0_i_9" *) 
  LUT3 #(
    .INIT(8'h47)) 
    \addr[3]_INST_0_i_9_replica 
       (.I0(din[2]),
        .I1(p_2_in88_in),
        .I2(r_code[2]),
        .O(\addr[3]_INST_0_i_9_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBB8BBB8BBBBBBB8)) 
    \addr[4]_INST_0 
       (.I0(irqaddr[4]),
        .I1(\addr[15]_INST_0_i_5_n_0 ),
        .I2(\addr[4]_INST_0_i_1_n_0 ),
        .I3(\addr[4]_INST_0_i_2_n_0 ),
        .I4(\rrs[0][4]_repN ),
        .I5(\addr[15]_INST_0_i_1_n_0 ),
        .O(addr[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000FFB8B8)) 
    \addr[4]_INST_0_i_1 
       (.I0(data3[4]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[4]_INST_0_i_4_n_0 ),
        .I3(\addr[4]_INST_0_i_5_n_0 ),
        .I4(\addr[15]_INST_0_i_17_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[4]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[4]_INST_0_i_10 
       (.I0(\addr[7]_INST_0_i_23_n_7 ),
        .I1(p_4_in),
        .I2(pc[4]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[4]),
        .O(\addr[4]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[4]_INST_0_i_11 
       (.I0(\r_reg[15] [4]),
        .I1(\r_reg[14] [4]),
        .I2(soc[2]),
        .I3(\r_reg[13] [4]),
        .I4(soc[1]),
        .I5(\r_reg[12] [4]),
        .O(\addr[4]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[4]_INST_0_i_12 
       (.I0(\r_reg[11] [4]),
        .I1(\r_reg[10] [4]),
        .I2(soc[2]),
        .I3(\r_reg[9] [4]),
        .I4(soc[1]),
        .I5(\r_reg[8] [4]),
        .O(\addr[4]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[4]_INST_0_i_13 
       (.I0(\r_reg[7] [4]),
        .I1(\r_reg[6] [4]),
        .I2(soc[2]),
        .I3(\r_reg[5] [4]),
        .I4(soc[1]),
        .I5(\r_reg[4] [4]),
        .O(\addr[4]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF000F0FF55335533)) 
    \addr[4]_INST_0_i_14 
       (.I0(sp_reg[4]),
        .I1(pc[4]),
        .I2(\addr[15]_INST_0_i_20_n_0 ),
        .I3(soc[1]),
        .I4(\addr[4]_INST_0_i_8_n_0 ),
        .I5(soc[2]),
        .O(\addr[4]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[4]_INST_0_i_15 
       (.I0(\r_reg[11] [4]),
        .I1(\r_reg[10] [4]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [4]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [4]),
        .O(\addr[4]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[4]_INST_0_i_16 
       (.I0(\r_reg[15] [4]),
        .I1(\r_reg[14] [4]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [4]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [4]),
        .O(\addr[4]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[4]_INST_0_i_17 
       (.I0(\r_reg[7] [4]),
        .I1(\r_reg[6] [4]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [4]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [4]),
        .O(\addr[4]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000282020080)) 
    \addr[4]_INST_0_i_2 
       (.I0(sp_reg[4]),
        .I1(state[2]),
        .I2(state[3]),
        .I3(state[0]),
        .I4(state[1]),
        .I5(state[4]),
        .O(\addr[4]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "addr[4]_INST_0_i_3" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEFEEEEEE)) 
    \addr[4]_INST_0_i_3_replica 
       (.I0(\addr[4]_INST_0_i_6_n_0 ),
        .I1(\addr[4]_INST_0_i_7_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\addr[4]_INST_0_i_8_n_0 ),
        .I4(\addr[14]_INST_0_i_5_n_0 ),
        .I5(\addr[4]_INST_0_i_9_n_0 ),
        .O(\rrs[0][4]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFBAAA)) 
    \addr[4]_INST_0_i_3_rewire 
       (.I0(\addr[4]_INST_0_i_6_n_0 ),
        .I1(\r_code[3]_i_1_n_0 ),
        .I2(\addr[4]_INST_0_i_8_n_0 ),
        .I3(\addr[14]_INST_0_i_5_n_0 ),
        .I4(\addr[4]_INST_0_i_9_n_0 ),
        .O(\rrs[0] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[4]_INST_0_i_4 
       (.I0(\addr[4]_INST_0_i_10_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[4]),
        .I3(state[0]),
        .I4(plusOp4_out[4]),
        .O(\addr[4]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAACCAACCF0FFF000)) 
    \addr[4]_INST_0_i_5 
       (.I0(\addr[4]_INST_0_i_11_n_0 ),
        .I1(\addr[4]_INST_0_i_12_n_0 ),
        .I2(\addr[4]_INST_0_i_13_n_0 ),
        .I3(\r_code[10]_i_1_n_0 ),
        .I4(\addr[4]_INST_0_i_14_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\addr[4]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEA202A00000000)) 
    \addr[4]_INST_0_i_6 
       (.I0(\addr[4]_INST_0_i_15_n_0 ),
        .I1(din[2]),
        .I2(p_2_in88_in),
        .I3(r_code[2]),
        .I4(\addr[4]_INST_0_i_16_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\addr[4]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA0000A808)) 
    \addr[4]_INST_0_i_7 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(pc[4]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(sp_reg[4]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_9_n_0 ),
        .O(\addr[4]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "addr[4]_INST_0_i_7" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA0000A808)) 
    \addr[4]_INST_0_i_7_replica 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(pc[4]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(sp_reg[4]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_9_n_0 ),
        .O(\addr[4]_INST_0_i_7_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00002020000A202A)) 
    \addr[4]_INST_0_i_8 
       (.I0(\sr_reg_n_0_[4] ),
        .I1(din[4]),
        .I2(p_2_in88_in),
        .I3(r_code[4]),
        .I4(din[5]),
        .I5(r_code[5]),
        .O(\addr[4]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000505030000000)) 
    \addr[4]_INST_0_i_9 
       (.I0(r_code[3]),
        .I1(din[3]),
        .I2(\addr[4]_INST_0_i_17_n_0 ),
        .I3(din[2]),
        .I4(p_2_in88_in),
        .I5(r_code[2]),
        .O(\addr[4]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4F44)) 
    \addr[5]_INST_0 
       (.I0(\addr[15]_INST_0_i_1_n_0 ),
        .I1(\rrs[0] [5]),
        .I2(\addr[15]_INST_0_i_3_n_0 ),
        .I3(sp_reg[5]),
        .I4(\addr[5]_INST_0_i_2_n_0 ),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(addr[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF00D5)) 
    \addr[5]_INST_0_i_1 
       (.I0(\addr[5]_INST_0_i_3_n_0 ),
        .I1(\addr[5]_INST_0_i_4_n_0 ),
        .I2(\addr[14]_INST_0_i_5_n_0 ),
        .I3(\r_code[3]_i_1_n_0 ),
        .I4(\addr[5]_INST_0_i_5_n_0 ),
        .I5(\addr[5]_INST_0_i_6_n_0 ),
        .O(\rrs[0] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[5]_INST_0_i_10 
       (.I0(\r_reg[11] [5]),
        .I1(\r_reg[10] [5]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [5]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [5]),
        .O(\addr[5]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[5]_INST_0_i_11 
       (.I0(\r_reg[15] [5]),
        .I1(\r_reg[14] [5]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [5]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [5]),
        .O(\addr[5]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[5]_INST_0_i_12 
       (.I0(\addr[7]_INST_0_i_23_n_6 ),
        .I1(p_4_in),
        .I2(pc[5]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[5]),
        .O(\addr[5]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[5]_INST_0_i_13 
       (.I0(\r_reg[15] [5]),
        .I1(\r_reg[14] [5]),
        .I2(soc[2]),
        .I3(\r_reg[13] [5]),
        .I4(soc[1]),
        .I5(\r_reg[12] [5]),
        .O(\addr[5]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[5]_INST_0_i_14 
       (.I0(\r_reg[11] [5]),
        .I1(\r_reg[10] [5]),
        .I2(soc[2]),
        .I3(\r_reg[9] [5]),
        .I4(soc[1]),
        .I5(\r_reg[8] [5]),
        .O(\addr[5]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5F50CFCF5F50C0C0)) 
    \addr[5]_INST_0_i_15 
       (.I0(\addr[15]_INST_0_i_20_n_0 ),
        .I1(\addr[5]_INST_0_i_4_n_0 ),
        .I2(soc[2]),
        .I3(sp_reg[5]),
        .I4(soc[1]),
        .I5(pc[5]),
        .O(\addr[5]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[5]_INST_0_i_16 
       (.I0(\r_reg[7] [5]),
        .I1(\r_reg[6] [5]),
        .I2(soc[2]),
        .I3(\r_reg[5] [5]),
        .I4(soc[1]),
        .I5(\r_reg[4] [5]),
        .O(\addr[5]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000FFB8B8)) 
    \addr[5]_INST_0_i_2 
       (.I0(data3[5]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[5]_INST_0_i_7_n_0 ),
        .I3(\addr[5]_INST_0_i_8_n_0 ),
        .I4(\addr[15]_INST_0_i_17_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[5]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    \addr[5]_INST_0_i_3 
       (.I0(r_code[2]),
        .I1(p_2_in88_in),
        .I2(din[2]),
        .I3(\addr[5]_INST_0_i_9_n_0 ),
        .O(\addr[5]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00002020000A202A)) 
    \addr[5]_INST_0_i_4 
       (.I0(\sr_reg_n_0_[5] ),
        .I1(din[4]),
        .I2(p_2_in88_in),
        .I3(r_code[4]),
        .I4(din[5]),
        .I5(r_code[5]),
        .O(\addr[5]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA0000A808)) 
    \addr[5]_INST_0_i_5 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(pc[5]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(sp_reg[5]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_9_n_0 ),
        .O(\addr[5]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEA202A00000000)) 
    \addr[5]_INST_0_i_6 
       (.I0(\addr[5]_INST_0_i_10_n_0 ),
        .I1(din[2]),
        .I2(p_2_in88_in),
        .I3(r_code[2]),
        .I4(\addr[5]_INST_0_i_11_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\addr[5]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[5]_INST_0_i_7 
       (.I0(\addr[5]_INST_0_i_12_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[5]),
        .I3(state[0]),
        .I4(plusOp4_out[5]),
        .O(\addr[5]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAACCCCFF000F0F)) 
    \addr[5]_INST_0_i_8 
       (.I0(\addr[5]_INST_0_i_13_n_0 ),
        .I1(\addr[5]_INST_0_i_14_n_0 ),
        .I2(\addr[5]_INST_0_i_15_n_0 ),
        .I3(\addr[5]_INST_0_i_16_n_0 ),
        .I4(\r_code[10]_i_1_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\addr[5]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[5]_INST_0_i_9 
       (.I0(\r_reg[7] [5]),
        .I1(\r_reg[6] [5]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [5]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [5]),
        .O(\addr[5]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4F44)) 
    \addr[6]_INST_0 
       (.I0(\addr[15]_INST_0_i_1_n_0 ),
        .I1(\rrs[0] [6]),
        .I2(\addr[15]_INST_0_i_3_n_0 ),
        .I3(sp_reg[6]),
        .I4(\addr[6]_INST_0_i_2_n_0 ),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(addr[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEFEEEEEE)) 
    \addr[6]_INST_0_i_1 
       (.I0(\addr[6]_INST_0_i_3_n_0 ),
        .I1(\addr[6]_INST_0_i_4_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\addr[6]_INST_0_i_5_n_0 ),
        .I4(\addr[14]_INST_0_i_5_n_0 ),
        .I5(\addr[6]_INST_0_i_6_n_0 ),
        .O(\rrs[0] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[6]_INST_0_i_10 
       (.I0(\r_reg[15] [6]),
        .I1(\r_reg[14] [6]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [6]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [6]),
        .O(\addr[6]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[6]_INST_0_i_11 
       (.I0(\r_reg[7] [6]),
        .I1(\r_reg[6] [6]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [6]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [6]),
        .O(\addr[6]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[6]_INST_0_i_12 
       (.I0(\addr[7]_INST_0_i_23_n_5 ),
        .I1(p_4_in),
        .I2(pc[6]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[6]),
        .O(\addr[6]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[6]_INST_0_i_13 
       (.I0(\r_reg[15] [6]),
        .I1(\r_reg[14] [6]),
        .I2(soc[2]),
        .I3(\r_reg[13] [6]),
        .I4(soc[1]),
        .I5(\r_reg[12] [6]),
        .O(\addr[6]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[6]_INST_0_i_14 
       (.I0(\r_reg[11] [6]),
        .I1(\r_reg[10] [6]),
        .I2(soc[2]),
        .I3(\r_reg[9] [6]),
        .I4(soc[1]),
        .I5(\r_reg[8] [6]),
        .O(\addr[6]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[6]_INST_0_i_15 
       (.I0(\r_reg[7] [6]),
        .I1(\r_reg[6] [6]),
        .I2(soc[2]),
        .I3(\r_reg[5] [6]),
        .I4(soc[1]),
        .I5(\r_reg[4] [6]),
        .O(\addr[6]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF000F0FF55335533)) 
    \addr[6]_INST_0_i_16 
       (.I0(sp_reg[6]),
        .I1(pc[6]),
        .I2(\addr[15]_INST_0_i_20_n_0 ),
        .I3(soc[1]),
        .I4(\addr[6]_INST_0_i_5_n_0 ),
        .I5(soc[2]),
        .O(\addr[6]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000FFB8B8)) 
    \addr[6]_INST_0_i_2 
       (.I0(data3[6]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[6]_INST_0_i_7_n_0 ),
        .I3(\addr[6]_INST_0_i_8_n_0 ),
        .I4(\addr[15]_INST_0_i_17_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[6]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEA202A00000000)) 
    \addr[6]_INST_0_i_3 
       (.I0(\addr[6]_INST_0_i_9_n_0 ),
        .I1(din[2]),
        .I2(p_2_in88_in),
        .I3(r_code[2]),
        .I4(\addr[6]_INST_0_i_10_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\addr[6]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA0000A808)) 
    \addr[6]_INST_0_i_4 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(pc[6]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(sp_reg[6]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_9_n_0 ),
        .O(\addr[6]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00002020000A202A)) 
    \addr[6]_INST_0_i_5 
       (.I0(\sr_reg_n_0_[6] ),
        .I1(din[4]),
        .I2(p_2_in88_in),
        .I3(r_code[4]),
        .I4(din[5]),
        .I5(r_code[5]),
        .O(\addr[6]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3000505030000000)) 
    \addr[6]_INST_0_i_6 
       (.I0(r_code[3]),
        .I1(din[3]),
        .I2(\addr[6]_INST_0_i_11_n_0 ),
        .I3(din[2]),
        .I4(p_2_in88_in),
        .I5(r_code[2]),
        .O(\addr[6]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[6]_INST_0_i_7 
       (.I0(\addr[6]_INST_0_i_12_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[6]),
        .I3(state[0]),
        .I4(plusOp4_out[6]),
        .O(\addr[6]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAACCAACCF0FFF000)) 
    \addr[6]_INST_0_i_8 
       (.I0(\addr[6]_INST_0_i_13_n_0 ),
        .I1(\addr[6]_INST_0_i_14_n_0 ),
        .I2(\addr[6]_INST_0_i_15_n_0 ),
        .I3(\r_code[10]_i_1_n_0 ),
        .I4(\addr[6]_INST_0_i_16_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\addr[6]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[6]_INST_0_i_9 
       (.I0(\r_reg[11] [6]),
        .I1(\r_reg[10] [6]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [6]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [6]),
        .O(\addr[6]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4F44)) 
    \addr[7]_INST_0 
       (.I0(\addr[15]_INST_0_i_1_n_0 ),
        .I1(\rrs[0][7]_repN ),
        .I2(\addr[15]_INST_0_i_3_n_0 ),
        .I3(sp_reg[7]),
        .I4(\addr[7]_INST_0_i_2_n_0 ),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(addr[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[7]_INST_0_i_10 
       (.I0(\r_reg[11] [7]),
        .I1(\r_reg[10] [7]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [7]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [7]),
        .O(\addr[7]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[7]_INST_0_i_11 
       (.I0(\r_reg[7] [7]),
        .I1(\r_reg[6] [7]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [7]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [7]),
        .O(\addr[7]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h36)) 
    \addr[7]_INST_0_i_12_rewire 
       (.I0(\addr[7]_INST_0_i_5_n_0 ),
        .I1(din[7]),
        .I2(\rrs[0] [7]),
        .O(\addr[7]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[7]_INST_0_i_13 
       (.I0(din[6]),
        .I1(\rrs[0] [6]),
        .O(\addr[7]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[7]_INST_0_i_14 
       (.I0(din[5]),
        .I1(\rrs[0] [5]),
        .O(\addr[7]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h36)) 
    \addr[7]_INST_0_i_15_rewire 
       (.I0(\addr[4]_INST_0_i_7_n_0 ),
        .I1(din[4]),
        .I2(\rrs[0] [4]),
        .O(\addr[7]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[7]_INST_0_i_16 
       (.I0(\addr[7]_INST_0_i_23_n_4 ),
        .I1(p_4_in),
        .I2(pc[7]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[7]),
        .O(\addr[7]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[7]_INST_0_i_17 
       (.CI(\addr[3]_INST_0_i_17_n_0 ),
        .CO({\addr[7]_INST_0_i_17_n_0 ,\addr[7]_INST_0_i_17_n_1 ,\addr[7]_INST_0_i_17_n_2 ,\addr[7]_INST_0_i_17_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(din[7:4]),
        .O(plusOp3_out[7:4]),
        .S({\addr[7]_INST_0_i_25_n_0 ,\addr[7]_INST_0_i_26_n_0 ,\addr[7]_INST_0_i_27_n_0 ,\addr[7]_INST_0_i_28_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[7]_INST_0_i_18 
       (.CI(\addr[3]_INST_0_i_18_n_0 ),
        .CO({\addr[7]_INST_0_i_18_n_0 ,\addr[7]_INST_0_i_18_n_1 ,\addr[7]_INST_0_i_18_n_2 ,\addr[7]_INST_0_i_18_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(din[7:4]),
        .O(plusOp4_out[7:4]),
        .S({\addr[7]_INST_0_i_29_n_0 ,\addr[7]_INST_0_i_30_n_0 ,\addr[7]_INST_0_i_31_n_0 ,\addr[7]_INST_0_i_32_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \addr[7]_INST_0_i_19 
       (.I0(\addr[7]_INST_0_i_33_n_0 ),
        .I1(\addr[7]_INST_0_i_34_n_0 ),
        .O(\addr[7]_INST_0_i_19_n_0 ),
        .S(\r_code[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "addr[7]_INST_0_i_1" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF10000)) 
    \addr[7]_INST_0_i_1_replica 
       (.I0(\addr[7]_INST_0_i_3_n_0 ),
        .I1(\addr[15]_INST_0_i_8_n_0 ),
        .I2(\addr[7]_INST_0_i_4_n_0 ),
        .I3(\addr[15]_INST_0_i_9_n_0 ),
        .I4(\addr[15]_INST_0_i_11_n_0 ),
        .I5(\addr[7]_INST_0_i_5_n_0 ),
        .O(\rrs[0][7]_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF10000)) 
    \addr[7]_INST_0_i_1_rewire 
       (.I0(\addr[7]_INST_0_i_3_n_0 ),
        .I1(\addr[15]_INST_0_i_8_n_0 ),
        .I2(\addr[7]_INST_0_i_4_n_0 ),
        .I3(\addr[15]_INST_0_i_9_n_0 ),
        .I4(\addr[15]_INST_0_i_11_n_0 ),
        .O(\rrs[0] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000FFB8B8)) 
    \addr[7]_INST_0_i_2 
       (.I0(data3[7]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[7]_INST_0_i_7_n_0 ),
        .I3(\addr[7]_INST_0_i_8_n_0 ),
        .I4(\addr[15]_INST_0_i_17_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[7]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000000E2)) 
    \addr[7]_INST_0_i_20 
       (.I0(pc[7]),
        .I1(soc[1]),
        .I2(sp_reg[7]),
        .I3(\r_code[10]_i_1_n_0 ),
        .I4(soc[2]),
        .O(\addr[7]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[7]_INST_0_i_21 
       (.I0(\r_reg[7] [7]),
        .I1(\r_reg[6] [7]),
        .I2(soc[2]),
        .I3(\r_reg[5] [7]),
        .I4(soc[1]),
        .I5(\r_reg[4] [7]),
        .O(\addr[7]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000002022220020)) 
    \addr[7]_INST_0_i_22 
       (.I0(soc[2]),
        .I1(\r_code[10]_i_1_n_0 ),
        .I2(\sr_reg_n_0_[7] ),
        .I3(lbe_INST_0_i_8_n_0),
        .I4(soc[1]),
        .I5(\addr[15]_INST_0_i_20_n_0 ),
        .O(\addr[7]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[7]_INST_0_i_23 
       (.CI(\addr[3]_INST_0_i_23_n_0 ),
        .CO({\addr[7]_INST_0_i_23_n_0 ,\addr[7]_INST_0_i_23_n_1 ,\addr[7]_INST_0_i_23_n_2 ,\addr[7]_INST_0_i_23_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(bsaddr__0[7:4]),
        .O({\addr[7]_INST_0_i_23_n_4 ,\addr[7]_INST_0_i_23_n_5 ,\addr[7]_INST_0_i_23_n_6 ,\addr[7]_INST_0_i_23_n_7 }),
        .S({\addr[7]_INST_0_i_35_n_0 ,\addr[7]_INST_0_i_36_n_0 ,\addr[7]_INST_0_i_37_n_0 ,\addr[7]_INST_0_i_38_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[7]_INST_0_i_24 
       (.CI(\addr[3]_INST_0_i_24_n_0 ),
        .CO({\addr[7]_INST_0_i_24_n_0 ,\addr[7]_INST_0_i_24_n_1 ,\addr[7]_INST_0_i_24_n_2 ,\addr[7]_INST_0_i_24_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(bsaddr__0[7:4]),
        .O(plusOp2_out[7:4]),
        .S({\addr[7]_INST_0_i_39_n_0 ,\addr[7]_INST_0_i_40_n_0 ,\addr[7]_INST_0_i_41_n_0 ,\addr[7]_INST_0_i_42_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[7]_INST_0_i_25 
       (.I0(din[7]),
        .I1(\rrd[0] [7]),
        .O(\addr[7]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[7]_INST_0_i_26 
       (.I0(din[6]),
        .I1(\rrd[0] [6]),
        .O(\addr[7]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h36)) 
    \addr[7]_INST_0_i_27_rewire 
       (.I0(\addr[5]_INST_0_i_6_n_0 ),
        .I1(din[5]),
        .I2(\rrd[0] [5]),
        .O(\addr[7]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[7]_INST_0_i_28 
       (.I0(din[4]),
        .I1(\rrd[0] [4]),
        .O(\addr[7]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[7]_INST_0_i_29 
       (.I0(din[7]),
        .I1(\addr[7]_INST_0_i_8_n_0 ),
        .O(\addr[7]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFBBFCB8FFFFFFFF)) 
    \addr[7]_INST_0_i_3 
       (.I0(din[4]),
        .I1(p_2_in88_in),
        .I2(r_code[4]),
        .I3(din[5]),
        .I4(r_code[5]),
        .I5(\sr_reg_n_0_[7] ),
        .O(\addr[7]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[7]_INST_0_i_30 
       (.I0(din[6]),
        .I1(\addr[6]_INST_0_i_8_n_0 ),
        .O(\addr[7]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[7]_INST_0_i_31 
       (.I0(din[5]),
        .I1(\addr[5]_INST_0_i_8_n_0 ),
        .O(\addr[7]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[7]_INST_0_i_32 
       (.I0(din[4]),
        .I1(\addr[4]_INST_0_i_5_n_0 ),
        .O(\addr[7]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[7]_INST_0_i_33 
       (.I0(\r_reg[11] [7]),
        .I1(\r_reg[10] [7]),
        .I2(soc[2]),
        .I3(\r_reg[9] [7]),
        .I4(soc[1]),
        .I5(\r_reg[8] [7]),
        .O(\addr[7]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[7]_INST_0_i_34 
       (.I0(\r_reg[15] [7]),
        .I1(\r_reg[14] [7]),
        .I2(soc[2]),
        .I3(\r_reg[13] [7]),
        .I4(soc[1]),
        .I5(\r_reg[12] [7]),
        .O(\addr[7]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[7]_INST_0_i_35 
       (.I0(bsaddr__0[7]),
        .I1(\addr[7]_INST_0_i_8_n_0 ),
        .O(\addr[7]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[7]_INST_0_i_36 
       (.I0(bsaddr__0[6]),
        .I1(\addr[6]_INST_0_i_8_n_0 ),
        .O(\addr[7]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[7]_INST_0_i_37 
       (.I0(bsaddr__0[5]),
        .I1(\addr[5]_INST_0_i_8_n_0 ),
        .O(\addr[7]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \addr[7]_INST_0_i_38 
       (.I0(bsaddr__0[4]),
        .I1(\addr[4]_INST_0_i_5_n_0 ),
        .O(\addr[7]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h36)) 
    \addr[7]_INST_0_i_39_rewire 
       (.I0(\addr[7]_INST_0_i_5_n_0 ),
        .I1(bsaddr__0[7]),
        .I2(\rrs[0] [7]),
        .O(\addr[7]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \addr[7]_INST_0_i_4 
       (.I0(pc[7]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(sp_reg[7]),
        .I3(\r_code[1]_i_1_n_0 ),
        .O(\addr[7]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[7]_INST_0_i_40 
       (.I0(bsaddr__0[6]),
        .I1(\rrs[0] [6]),
        .O(\addr[7]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \addr[7]_INST_0_i_41 
       (.I0(bsaddr__0[5]),
        .I1(\rrs[0] [5]),
        .O(\addr[7]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h36)) 
    \addr[7]_INST_0_i_42_rewire 
       (.I0(\addr[4]_INST_0_i_7_n_0 ),
        .I1(bsaddr__0[4]),
        .I2(\rrs[0] [4]),
        .O(\addr[7]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFEEEAAAA)) 
    \addr[7]_INST_0_i_43 
       (.I0(\addr[7]_INST_0_i_5_n_0 ),
        .I1(\addr[7]_INST_0_i_4_n_0 ),
        .I2(\addr[3]_INST_0_i_47_n_0 ),
        .I3(\sr_reg_n_0_[7] ),
        .I4(\addr[15]_INST_0_i_11_n_0 ),
        .O(\rrd[0] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEEAAA)) 
    \addr[7]_INST_0_i_44 
       (.I0(\addr[6]_INST_0_i_3_n_0 ),
        .I1(\addr[15]_INST_0_i_11_n_0 ),
        .I2(\sr_reg_n_0_[6] ),
        .I3(\addr[3]_INST_0_i_47_n_0 ),
        .I4(\addr[7]_INST_0_i_47_n_0 ),
        .I5(\addr[6]_INST_0_i_6_n_0 ),
        .O(\rrd[0] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h888F)) 
    \addr[7]_INST_0_i_45_rewire 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(\addr[7]_INST_0_i_48_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\addr[5]_INST_0_i_3_n_0 ),
        .O(\rrd[0] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEEAAA)) 
    \addr[7]_INST_0_i_46 
       (.I0(\addr[4]_INST_0_i_6_n_0 ),
        .I1(\addr[15]_INST_0_i_11_n_0 ),
        .I2(\addr[3]_INST_0_i_47_n_0 ),
        .I3(\sr_reg_n_0_[4] ),
        .I4(\addr[7]_INST_0_i_49_n_0 ),
        .I5(\addr[4]_INST_0_i_9_n_0 ),
        .O(\rrd[0] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \addr[7]_INST_0_i_47 
       (.I0(pc[6]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(sp_reg[6]),
        .I3(\r_code[1]_i_1_n_0 ),
        .O(\addr[7]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF454045404540)) 
    \addr[7]_INST_0_i_48 
       (.I0(\r_code[1]_i_1_n_0 ),
        .I1(sp_reg[5]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(pc[5]),
        .I4(\addr[3]_INST_0_i_47_n_0 ),
        .I5(\sr_reg_n_0_[5] ),
        .O(\addr[7]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \addr[7]_INST_0_i_49 
       (.I0(pc[4]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(sp_reg[4]),
        .I3(\r_code[1]_i_1_n_0 ),
        .O(\addr[7]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC0C0AFA0)) 
    \addr[7]_INST_0_i_5 
       (.I0(\addr[7]_INST_0_i_9_n_0 ),
        .I1(\addr[7]_INST_0_i_10_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\addr[7]_INST_0_i_11_n_0 ),
        .I4(\addr[3]_INST_0_i_9_n_0 ),
        .O(\addr[7]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \addr[7]_INST_0_i_6 
       (.CI(\addr[3]_INST_0_i_4_n_0 ),
        .CO({\addr[7]_INST_0_i_6_n_0 ,\addr[7]_INST_0_i_6_n_1 ,\addr[7]_INST_0_i_6_n_2 ,\addr[7]_INST_0_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(din[7:4]),
        .O(data3[7:4]),
        .S({\addr[7]_INST_0_i_12_n_0 ,\addr[7]_INST_0_i_13_n_0 ,\addr[7]_INST_0_i_14_n_0 ,\addr[7]_INST_0_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[7]_INST_0_i_7 
       (.I0(\addr[7]_INST_0_i_16_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[7]),
        .I3(state[0]),
        .I4(plusOp4_out[7]),
        .O(\addr[7]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888888888B8B8B)) 
    \addr[7]_INST_0_i_8 
       (.I0(\addr[7]_INST_0_i_19_n_0 ),
        .I1(\r_code[11]_i_1_n_0 ),
        .I2(\addr[7]_INST_0_i_20_n_0 ),
        .I3(\addr[7]_INST_0_i_21_n_0 ),
        .I4(\r_code[10]_i_1_n_0 ),
        .I5(\addr[7]_INST_0_i_22_n_0 ),
        .O(\addr[7]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[7]_INST_0_i_9 
       (.I0(\r_reg[15] [7]),
        .I1(\r_reg[14] [7]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [7]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [7]),
        .O(\addr[7]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4F44)) 
    \addr[8]_INST_0 
       (.I0(\addr[15]_INST_0_i_1_n_0 ),
        .I1(\rrs[0] [8]),
        .I2(\addr[15]_INST_0_i_3_n_0 ),
        .I3(sp_reg[8]),
        .I4(\addr[8]_INST_0_i_2_n_0 ),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(addr[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF00D5)) 
    \addr[8]_INST_0_i_1 
       (.I0(\addr[8]_INST_0_i_3_n_0 ),
        .I1(\addr[8]_INST_0_i_4_n_0 ),
        .I2(\addr[14]_INST_0_i_5_n_0 ),
        .I3(\r_code[3]_i_1_n_0 ),
        .I4(\addr[8]_INST_0_i_5_n_0 ),
        .I5(\addr[8]_INST_0_i_6_n_0 ),
        .O(\rrs[0] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[8]_INST_0_i_10 
       (.I0(\r_reg[11] [8]),
        .I1(\r_reg[10] [8]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [8]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [8]),
        .O(\addr[8]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[8]_INST_0_i_11 
       (.I0(\r_reg[15] [8]),
        .I1(\r_reg[14] [8]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [8]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [8]),
        .O(\addr[8]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[8]_INST_0_i_12 
       (.I0(\addr[11]_INST_0_i_24_n_7 ),
        .I1(p_4_in),
        .I2(pc[8]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[8]),
        .O(\addr[8]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[8]_INST_0_i_13 
       (.I0(\r_reg[15] [8]),
        .I1(\r_reg[14] [8]),
        .I2(soc[2]),
        .I3(\r_reg[13] [8]),
        .I4(soc[1]),
        .I5(\r_reg[12] [8]),
        .O(\addr[8]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[8]_INST_0_i_14 
       (.I0(\r_reg[11] [8]),
        .I1(\r_reg[10] [8]),
        .I2(soc[2]),
        .I3(\r_reg[9] [8]),
        .I4(soc[1]),
        .I5(\r_reg[8] [8]),
        .O(\addr[8]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5F50CFCF5F50C0C0)) 
    \addr[8]_INST_0_i_15 
       (.I0(\addr[15]_INST_0_i_20_n_0 ),
        .I1(\addr[8]_INST_0_i_4_n_0 ),
        .I2(soc[2]),
        .I3(sp_reg[8]),
        .I4(soc[1]),
        .I5(pc[8]),
        .O(\addr[8]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[8]_INST_0_i_16 
       (.I0(\r_reg[7] [8]),
        .I1(\r_reg[6] [8]),
        .I2(soc[2]),
        .I3(\r_reg[5] [8]),
        .I4(soc[1]),
        .I5(\r_reg[4] [8]),
        .O(\addr[8]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000FFB8B8)) 
    \addr[8]_INST_0_i_2 
       (.I0(data3[8]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[8]_INST_0_i_7_n_0 ),
        .I3(\addr[8]_INST_0_i_8_n_0 ),
        .I4(\addr[15]_INST_0_i_17_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[8]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    \addr[8]_INST_0_i_3 
       (.I0(r_code[2]),
        .I1(p_2_in88_in),
        .I2(din[2]),
        .I3(\addr[8]_INST_0_i_9_n_0 ),
        .O(\addr[8]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00002020000A202A)) 
    \addr[8]_INST_0_i_4 
       (.I0(\sr_reg_n_0_[8] ),
        .I1(din[4]),
        .I2(p_2_in88_in),
        .I3(r_code[4]),
        .I4(din[5]),
        .I5(r_code[5]),
        .O(\addr[8]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA0000A808)) 
    \addr[8]_INST_0_i_5 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(pc[8]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(sp_reg[8]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_9_n_0 ),
        .O(\addr[8]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEA202A00000000)) 
    \addr[8]_INST_0_i_6 
       (.I0(\addr[8]_INST_0_i_10_n_0 ),
        .I1(din[2]),
        .I2(p_2_in88_in),
        .I3(r_code[2]),
        .I4(\addr[8]_INST_0_i_11_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\addr[8]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[8]_INST_0_i_7 
       (.I0(\addr[8]_INST_0_i_12_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[8]),
        .I3(state[0]),
        .I4(plusOp4_out[8]),
        .O(\addr[8]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAACCCCFF000F0F)) 
    \addr[8]_INST_0_i_8 
       (.I0(\addr[8]_INST_0_i_13_n_0 ),
        .I1(\addr[8]_INST_0_i_14_n_0 ),
        .I2(\addr[8]_INST_0_i_15_n_0 ),
        .I3(\addr[8]_INST_0_i_16_n_0 ),
        .I4(\r_code[10]_i_1_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\addr[8]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[8]_INST_0_i_9 
       (.I0(\r_reg[7] [8]),
        .I1(\r_reg[6] [8]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [8]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [8]),
        .O(\addr[8]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4F44)) 
    \addr[9]_INST_0 
       (.I0(\addr[15]_INST_0_i_1_n_0 ),
        .I1(\rrs[0] [9]),
        .I2(\addr[15]_INST_0_i_3_n_0 ),
        .I3(sp_reg[9]),
        .I4(\addr[9]_INST_0_i_2_n_0 ),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(addr[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF00D5)) 
    \addr[9]_INST_0_i_1 
       (.I0(\addr[9]_INST_0_i_3_n_0 ),
        .I1(\addr[9]_INST_0_i_4_n_0 ),
        .I2(\addr[14]_INST_0_i_5_n_0 ),
        .I3(\r_code[3]_i_1_n_0 ),
        .I4(\addr[9]_INST_0_i_5_n_0 ),
        .I5(\addr[9]_INST_0_i_6_n_0 ),
        .O(\rrs[0] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[9]_INST_0_i_10 
       (.I0(\r_reg[11] [9]),
        .I1(\r_reg[10] [9]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[9] [9]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[8] [9]),
        .O(\addr[9]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[9]_INST_0_i_11 
       (.I0(\r_reg[15] [9]),
        .I1(\r_reg[14] [9]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[13] [9]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[12] [9]),
        .O(\addr[9]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \addr[9]_INST_0_i_12 
       (.I0(\addr[11]_INST_0_i_24_n_6 ),
        .I1(p_4_in),
        .I2(pc[9]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[9]),
        .O(\addr[9]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[9]_INST_0_i_13 
       (.I0(\r_reg[15] [9]),
        .I1(\r_reg[14] [9]),
        .I2(soc[2]),
        .I3(\r_reg[13] [9]),
        .I4(soc[1]),
        .I5(\r_reg[12] [9]),
        .O(\addr[9]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[9]_INST_0_i_14 
       (.I0(\r_reg[11] [9]),
        .I1(\r_reg[10] [9]),
        .I2(soc[2]),
        .I3(\r_reg[9] [9]),
        .I4(soc[1]),
        .I5(\r_reg[8] [9]),
        .O(\addr[9]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5F50CFCF5F50C0C0)) 
    \addr[9]_INST_0_i_15 
       (.I0(\addr[15]_INST_0_i_20_n_0 ),
        .I1(\addr[9]_INST_0_i_4_n_0 ),
        .I2(soc[2]),
        .I3(sp_reg[9]),
        .I4(soc[1]),
        .I5(pc[9]),
        .O(\addr[9]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \addr[9]_INST_0_i_16 
       (.I0(\r_reg[7] [9]),
        .I1(\r_reg[6] [9]),
        .I2(soc[2]),
        .I3(\r_reg[5] [9]),
        .I4(soc[1]),
        .I5(\r_reg[4] [9]),
        .O(\addr[9]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000FFB8B8)) 
    \addr[9]_INST_0_i_2 
       (.I0(data3[9]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(\addr[9]_INST_0_i_7_n_0 ),
        .I3(\addr[9]_INST_0_i_8_n_0 ),
        .I4(\addr[15]_INST_0_i_17_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(\addr[9]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1DFF)) 
    \addr[9]_INST_0_i_3 
       (.I0(r_code[2]),
        .I1(p_2_in88_in),
        .I2(din[2]),
        .I3(\addr[9]_INST_0_i_9_n_0 ),
        .O(\addr[9]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00002020000A202A)) 
    \addr[9]_INST_0_i_4 
       (.I0(\sr_reg_n_0_[9] ),
        .I1(din[4]),
        .I2(p_2_in88_in),
        .I3(r_code[4]),
        .I4(din[5]),
        .I5(r_code[5]),
        .O(\addr[9]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA0000A808)) 
    \addr[9]_INST_0_i_5 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(pc[9]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(sp_reg[9]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\addr[15]_INST_0_i_9_n_0 ),
        .O(\addr[9]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEA202A00000000)) 
    \addr[9]_INST_0_i_6 
       (.I0(\addr[9]_INST_0_i_10_n_0 ),
        .I1(din[2]),
        .I2(p_2_in88_in),
        .I3(r_code[2]),
        .I4(\addr[9]_INST_0_i_11_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\addr[9]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \addr[9]_INST_0_i_7 
       (.I0(\addr[9]_INST_0_i_12_n_0 ),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[9]),
        .I3(state[0]),
        .I4(plusOp4_out[9]),
        .O(\addr[9]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAACCCCFF000F0F)) 
    \addr[9]_INST_0_i_8 
       (.I0(\addr[9]_INST_0_i_13_n_0 ),
        .I1(\addr[9]_INST_0_i_14_n_0 ),
        .I2(\addr[9]_INST_0_i_15_n_0 ),
        .I3(\addr[9]_INST_0_i_16_n_0 ),
        .I4(\r_code[10]_i_1_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\addr[9]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \addr[9]_INST_0_i_9 
       (.I0(\r_reg[7] [9]),
        .I1(\r_reg[6] [9]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_reg[5] [9]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[4] [9]),
        .O(\addr[9]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[0]_i_1 
       (.I0(din[0]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[10]_i_1 
       (.I0(din[10]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[11]_i_1 
       (.I0(din[11]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[12]_i_1 
       (.I0(din[12]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[13]_i_1 
       (.I0(din[13]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[14]_i_1 
       (.I0(din[14]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000484)) 
    \bsaddr[15]_i_1 
       (.I0(state[1]),
        .I1(state[0]),
        .I2(state[2]),
        .I3(state[3]),
        .I4(state[4]),
        .I5(halt),
        .O(\bsaddr[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[15]_i_2 
       (.I0(din[15]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[1]_i_1 
       (.I0(din[1]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[2]_i_1 
       (.I0(din[2]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[3]_i_1 
       (.I0(din[3]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[4]_i_1 
       (.I0(din[4]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[5]_i_1 
       (.I0(din[5]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[6]_i_1 
       (.I0(din[6]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[7]_i_1 
       (.I0(din[7]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[8]_i_1 
       (.I0(din[8]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAA8AAAA)) 
    \bsaddr[9]_i_1 
       (.I0(din[9]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(bsaddr[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[0] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[0]),
        .Q(bsaddr__0[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[10] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[10]),
        .Q(bsaddr__0[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[11] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[11]),
        .Q(bsaddr__0[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[12] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[12]),
        .Q(bsaddr__0[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[13] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[13]),
        .Q(bsaddr__0[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[14] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[14]),
        .Q(bsaddr__0[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[15] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[15]),
        .Q(bsaddr__0[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[1] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[1]),
        .Q(bsaddr__0[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[2] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[2]),
        .Q(bsaddr__0[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[3] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[3]),
        .Q(bsaddr__0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[4] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[4]),
        .Q(bsaddr__0[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[5] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[5]),
        .Q(bsaddr__0[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[6] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[6]),
        .Q(bsaddr__0[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[7] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[7]),
        .Q(bsaddr__0[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[8] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[8]),
        .Q(bsaddr__0[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \bsaddr_reg[9] 
       (.C(clk),
        .CE(\bsaddr[15]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bsaddr[9]),
        .Q(bsaddr__0[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[0]_INST_0 
       (.I0(pc[0]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(sr_reg_n_0_),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[0]_INST_0_i_1_n_0 ),
        .O(dout[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dout[0]_INST_0_i_1 
       (.I0(\dout[8]_INST_0_i_2_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\dout[0]_INST_0_i_2_n_0 ),
        .O(\dout[0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h550055C0FFFF55C0)) 
    \dout[0]_INST_0_i_10 
       (.I0(\addr[1]_INST_0_i_5_n_0 ),
        .I1(\dout[0]_INST_0_i_13_n_0 ),
        .I2(\dout[0]_INST_0_i_14_n_0 ),
        .I3(\dout[5]_INST_0_i_10_n_0 ),
        .I4(\FSM_sequential_state[1]_i_12_n_0 ),
        .I5(\rrs[0] [1]),
        .O(\dout[0]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[0]_INST_0_i_11 
       (.I0(\dout[2]_INST_0_i_17_n_0 ),
        .I1(\dout[9]_INST_0_i_18_n_0 ),
        .O(\dout[0]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0CFF0C0C00000404)) 
    \dout[0]_INST_0_i_12 
       (.I0(\dout[15]_INST_0_i_11_n_0 ),
        .I1(doc[0]),
        .I2(\dout[15]_INST_0_i_37_n_0 ),
        .I3(\dout[2]_INST_0_i_42_n_0 ),
        .I4(\dout[9]_INST_0_i_18_n_0 ),
        .I5(\dout[2]_INST_0_i_17_n_0 ),
        .O(\dout[0]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7777777744474444)) 
    \dout[0]_INST_0_i_13 
       (.I0(\r_code[0]_i_1_n_0 ),
        .I1(eqOp93_in),
        .I2(\dout[13]_INST_0_i_3_n_0 ),
        .I3(rd_INST_0_i_16_n_0),
        .I4(rd_INST_0_i_21_n_0),
        .I5(\dout[2]_INST_0_i_38_n_0 ),
        .O(\dout[0]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFDFF)) 
    \dout[0]_INST_0_i_14 
       (.I0(src__0[1]),
        .I1(\dout[13]_INST_0_i_3_n_0 ),
        .I2(rd_INST_0_i_16_n_0),
        .I3(rd_INST_0_i_21_n_0),
        .O(\dout[0]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFEEE)) 
    \dout[0]_INST_0_i_2 
       (.I0(\dout[0]_INST_0_i_3_n_0 ),
        .I1(\dout[0]_INST_0_i_4_n_0 ),
        .I2(\dout[0]_INST_0_i_5_n_0 ),
        .I3(\dout[6]_INST_0_i_5_n_0 ),
        .I4(\dout[0]_INST_0_i_6_n_0 ),
        .O(\dout[0]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF222F222F222)) 
    \dout[0]_INST_0_i_3 
       (.I0(\dout[15]_INST_0_i_14_n_0 ),
        .I1(\dout[2]_INST_0_i_45_n_0 ),
        .I2(\dout[2]_INST_0_i_6_n_7 ),
        .I3(\dout[4]_INST_0_i_7_n_0 ),
        .I4(\dout[2]_INST_0_i_7_n_7 ),
        .I5(eqOp93_in),
        .O(\dout[0]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \dout[0]_INST_0_i_4 
       (.I0(\dout[0]_INST_0_i_7_n_0 ),
        .I1(\dout[0]_INST_0_i_8_n_0 ),
        .I2(\dout[15]_INST_0_i_23_n_0 ),
        .I3(\dout[2]_INST_0_i_11_n_7 ),
        .I4(\dout[15]_INST_0_i_19_n_0 ),
        .I5(\dout[0]_INST_0_i_9_n_0 ),
        .O(\dout[0]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \dout[0]_INST_0_i_5 
       (.I0(\dout[15]_INST_0_i_11_n_0 ),
        .I1(\dout[0]_INST_0_i_10_n_0 ),
        .O(\dout[0]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0505110000000000)) 
    \dout[0]_INST_0_i_6 
       (.I0(soc[1]),
        .I1(\dout[9]_INST_0_i_11_n_0 ),
        .I2(\dout[2]_INST_0_i_45_n_0 ),
        .I3(soc[0]),
        .I4(soc[2]),
        .I5(eqOp135_in),
        .O(\dout[0]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF444)) 
    \dout[0]_INST_0_i_7 
       (.I0(\dout[2]_INST_0_i_35_n_0 ),
        .I1(\dout[14]_INST_0_i_10_n_0 ),
        .I2(\dout[0]_INST_0_i_11_n_0 ),
        .I3(\dout[14]_INST_0_i_11_n_0 ),
        .I4(\dout[0]_INST_0_i_12_n_0 ),
        .O(\dout[0]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT4 #(
    .INIT(16'h1441)) 
    \dout[0]_INST_0_i_8 
       (.I0(bw),
        .I1(\dout[2]_INST_0_i_45_n_0 ),
        .I2(\dout[2]_INST_0_i_17_n_0 ),
        .I3(sr_reg_n_0_),
        .O(\dout[0]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55404040)) 
    \dout[0]_INST_0_i_9 
       (.I0(bw),
        .I1(\dout[2]_INST_0_i_30_n_7 ),
        .I2(\dout[15]_INST_0_i_20_n_0 ),
        .I3(\dout[2]_INST_0_i_31_n_7 ),
        .I4(\dout[15]_INST_0_i_31_n_0 ),
        .O(\dout[0]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[10]_INST_0 
       (.I0(pc[10]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[10] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[10]_INST_0_i_1_n_0 ),
        .O(dout[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00A2)) 
    \dout[10]_INST_0_i_1 
       (.I0(\dout[10]_INST_0_i_2_n_0 ),
        .I1(\dout[13]_INST_0_i_3_n_0 ),
        .I2(\dout[10]_INST_0_i_3_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[10]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7400FF74)) 
    \dout[10]_INST_0_i_10 
       (.I0(sr_reg_n_0_),
        .I1(bw),
        .I2(\dout[9]_INST_0_i_12_n_0 ),
        .I3(\dout[9]_INST_0_i_11_n_0 ),
        .I4(L[8]),
        .O(\dout[10]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[10]_INST_0_i_11 
       (.I0(L[9]),
        .I1(\dout[9]_INST_0_i_14_n_0 ),
        .O(\dout[15]_INST_0_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "dout[10]_INST_0_i_11" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[10]_INST_0_i_11_replica 
       (.I0(L[9]),
        .I1(\dout[9]_INST_0_i_14_n_0 ),
        .O(\dout[15]_INST_0_i_80_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[10]_INST_0_i_12 
       (.I0(L[9]),
        .I1(\dout[9]_INST_0_i_14_n_0 ),
        .O(\dout[10]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[10]_INST_0_i_13 
       (.I0(L[10]),
        .I1(\dout[2]_INST_0_i_12_n_0 ),
        .O(\dout[15]_INST_0_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \dout[10]_INST_0_i_14 
       (.I0(\dout[15]_INST_0_i_20_n_0 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_39_n_5 ),
        .O(\dout[10]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABAAABBB)) 
    \dout[10]_INST_0_i_15 
       (.I0(\dout[15]_INST_0_i_37_n_0 ),
        .I1(\dout[2]_INST_0_i_12_n_0 ),
        .I2(din[12]),
        .I3(p_2_in88_in),
        .I4(r_code[12]),
        .O(\dout[10]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB800B800B800)) 
    \dout[10]_INST_0_i_16 
       (.I0(\dout[15]_INST_0_i_66_n_5 ),
        .I1(bw),
        .I2(\dout[15]_INST_0_i_71_n_5 ),
        .I3(\dout[15]_INST_0_i_31_n_0 ),
        .I4(\dout[4]_INST_0_i_7_n_0 ),
        .I5(\dout[15]_INST_0_i_61_n_5 ),
        .O(\dout[10]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF33333222)) 
    \dout[10]_INST_0_i_2_rewire 
       (.I0(\dout[10]_INST_0_i_14_n_0 ),
        .I1(\dout[10]_INST_0_i_4_n_0 ),
        .I2(\dout[15]_INST_0_i_23_n_0 ),
        .I3(\dout[10]_INST_0_i_5_n_0 ),
        .I4(\dout[10]_INST_0_i_6_n_0 ),
        .I5(\dout[10]_INST_0_i_7_n_0 ),
        .O(\dout[10]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF8)) 
    \dout[10]_INST_0_i_3 
       (.I0(eqOp93_in),
        .I1(\dout[11]_INST_0_i_8_n_5 ),
        .I2(\dout[10]_INST_0_i_8_n_0 ),
        .I3(\dout[10]_INST_0_i_9_n_0 ),
        .O(\dout[10]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F444FFF44444444)) 
    \dout[10]_INST_0_i_4 
       (.I0(\dout[15]_INST_0_i_39_n_5 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_51_n_5 ),
        .I3(bw),
        .I4(\dout[15]_INST_0_i_56_n_5 ),
        .I5(\dout[15]_INST_0_i_20_n_0 ),
        .O(\dout[10]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h870078FF87FF7800)) 
    \dout[10]_INST_0_i_5 
       (.I0(\dout[10]_INST_0_i_10_n_0 ),
        .I1(\dout[15]_INST_0_i_80_n_0 ),
        .I2(\dout[10]_INST_0_i_12_n_0 ),
        .I3(\dout[9]_INST_0_i_5_n_0 ),
        .I4(\dout[15]_INST_0_i_79_n_0 ),
        .I5(\dout[11]_INST_0_i_14_n_0 ),
        .O(\dout[10]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0CAF0FF)) 
    \dout[10]_INST_0_i_6_rewire 
       (.I0(\dout[14]_INST_0_i_10_n_0 ),
        .I1(\dout[14]_INST_0_i_11_n_0 ),
        .I2(L[10]),
        .I3(\dout[2]_INST_0_i_12_n_0 ),
        .I4(\dout[10]_INST_0_i_15_n_0 ),
        .O(\dout[10]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEEFE)) 
    \dout[10]_INST_0_i_7 
       (.I0(\dout[10]_INST_0_i_3_n_0 ),
        .I1(\dout[10]_INST_0_i_16_n_0 ),
        .I2(\dout[15]_INST_0_i_14_n_0 ),
        .I3(\dout[2]_INST_0_i_12_n_0 ),
        .O(\dout[10]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0030005000000050)) 
    \dout[10]_INST_0_i_8 
       (.I0(\dout[11]_INST_0_i_16_n_0 ),
        .I1(soc[1]),
        .I2(eqOp135_in),
        .I3(soc[2]),
        .I4(soc[0]),
        .I5(\dout[2]_INST_0_i_5_n_0 ),
        .O(\dout[10]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCC80CC8000000C00)) 
    \dout[10]_INST_0_i_9 
       (.I0(soc[0]),
        .I1(eqOp135_in),
        .I2(soc[1]),
        .I3(soc[2]),
        .I4(\dout[2]_INST_0_i_12_n_0 ),
        .I5(\dout[13]_INST_0_i_21_n_0 ),
        .O(\dout[10]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[11]_INST_0 
       (.I0(pc[11]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[11] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[11]_INST_0_i_1_n_0 ),
        .O(dout[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00A2)) 
    \dout[11]_INST_0_i_1 
       (.I0(\dout[11]_INST_0_i_2_n_0 ),
        .I1(\dout[13]_INST_0_i_3_n_0 ),
        .I2(\dout[11]_INST_0_i_3_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[11]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCC80CC8000000C00)) 
    \dout[11]_INST_0_i_10 
       (.I0(soc[0]),
        .I1(eqOp135_in),
        .I2(soc[1]),
        .I3(soc[2]),
        .I4(\dout[11]_INST_0_i_16_n_0 ),
        .I5(\dout[13]_INST_0_i_21_n_0 ),
        .O(\dout[11]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h80F8)) 
    \dout[11]_INST_0_i_11 
       (.I0(\dout[10]_INST_0_i_10_n_0 ),
        .I1(\dout[15]_INST_0_i_80_n_0 ),
        .I2(\dout[15]_INST_0_i_79_n_0 ),
        .I3(\dout[10]_INST_0_i_12_n_0 ),
        .O(\dout[11]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[11]_INST_0_i_12 
       (.I0(L[11]),
        .I1(\dout[11]_INST_0_i_16_n_0 ),
        .O(\dout[15]_INST_0_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[11]_INST_0_i_13 
       (.I0(\dout[11]_INST_0_i_27_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\rrd[0] [10]),
        .I3(\dout[14]_INST_0_i_25_n_0 ),
        .I4(\dout[11]_INST_0_i_28_n_0 ),
        .O(L[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04545555FFFFFFFF)) 
    \dout[11]_INST_0_i_14 
       (.I0(\dout[11]_INST_0_i_29_n_0 ),
        .I1(\dout[9]_INST_0_i_12_n_0 ),
        .I2(bw),
        .I3(sr_reg_n_0_),
        .I4(\dout[11]_INST_0_i_30_n_0 ),
        .I5(\dout[11]_INST_0_i_31_n_0 ),
        .O(\dout[11]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \dout[11]_INST_0_i_15 
       (.I0(\dout[15]_INST_0_i_20_n_0 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_39_n_4 ),
        .O(\dout[11]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h2E)) 
    \dout[11]_INST_0_i_16 
       (.I0(\dout[11]_INST_0_i_32_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\dout[2]_INST_0_i_13_n_0 ),
        .O(\dout[11]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[11]_INST_0_i_17 
       (.I0(\dout[11]_INST_0_i_33_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\rrd[0] [11]),
        .I3(\dout[14]_INST_0_i_25_n_0 ),
        .I4(\dout[11]_INST_0_i_34_n_0 ),
        .O(L[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABAAABBB)) 
    \dout[11]_INST_0_i_18 
       (.I0(\dout[15]_INST_0_i_37_n_0 ),
        .I1(\dout[11]_INST_0_i_16_n_0 ),
        .I2(din[12]),
        .I3(p_2_in88_in),
        .I4(r_code[12]),
        .O(\dout[11]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB800B800B800)) 
    \dout[11]_INST_0_i_19 
       (.I0(\dout[15]_INST_0_i_66_n_4 ),
        .I1(bw),
        .I2(\dout[15]_INST_0_i_71_n_4 ),
        .I3(\dout[15]_INST_0_i_31_n_0 ),
        .I4(\dout[4]_INST_0_i_7_n_0 ),
        .I5(\dout[15]_INST_0_i_61_n_4 ),
        .O(\dout[11]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF5540)) 
    \dout[11]_INST_0_i_2 
       (.I0(\dout[11]_INST_0_i_4_n_0 ),
        .I1(\dout[15]_INST_0_i_23_n_0 ),
        .I2(\dout[11]_INST_0_i_5_n_0 ),
        .I3(\dout[11]_INST_0_i_6_n_0 ),
        .I4(\dout[11]_INST_0_i_7_n_0 ),
        .O(\dout[11]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[11]_INST_0_i_20 
       (.I0(\dout[11]_INST_0_i_35_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\rrd[0] [9]),
        .I3(\dout[14]_INST_0_i_25_n_0 ),
        .I4(\dout[11]_INST_0_i_36_n_0 ),
        .O(L[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[11]_INST_0_i_21 
       (.I0(\dout[11]_INST_0_i_37_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\rrd[0] [8]),
        .I3(\dout[14]_INST_0_i_25_n_0 ),
        .I4(\dout[11]_INST_0_i_38_n_0 ),
        .O(L[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \dout[11]_INST_0_i_22 
       (.I0(L[11]),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[11]_INST_0_i_16_n_0 ),
        .O(\dout[11]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \dout[11]_INST_0_i_23 
       (.I0(L[10]),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[2]_INST_0_i_12_n_0 ),
        .O(\dout[11]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \dout[11]_INST_0_i_24 
       (.I0(L[9]),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[9]_INST_0_i_14_n_0 ),
        .O(\dout[11]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \dout[11]_INST_0_i_25 
       (.I0(L[8]),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[9]_INST_0_i_11_n_0 ),
        .O(\dout[11]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000045450045)) 
    \dout[11]_INST_0_i_26 
       (.I0(\dout[2]_INST_0_i_37_n_0 ),
        .I1(\addr[3]_INST_0_i_6_n_0 ),
        .I2(\dout[5]_INST_0_i_10_n_0 ),
        .I3(\FSM_sequential_state[1]_i_12_n_0 ),
        .I4(\rrs[0] [3]),
        .I5(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[11]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[11]_INST_0_i_27 
       (.I0(\rrd[0] [2]),
        .I1(\dout[14]_INST_0_i_25_n_0 ),
        .I2(pc[2]),
        .I3(eqOp93_in),
        .I4(data4[2]),
        .O(\dout[11]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88B8B8B8)) 
    \dout[11]_INST_0_i_28 
       (.I0(pc[10]),
        .I1(eqOp93_in),
        .I2(din[10]),
        .I3(r_a0),
        .I4(bw),
        .O(\dout[11]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    \dout[11]_INST_0_i_29 
       (.I0(L[8]),
        .I1(\dout[9]_INST_0_i_11_n_0 ),
        .I2(\dout[10]_INST_0_i_12_n_0 ),
        .O(\dout[11]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF8)) 
    \dout[11]_INST_0_i_3 
       (.I0(eqOp93_in),
        .I1(\dout[11]_INST_0_i_8_n_4 ),
        .I2(\dout[11]_INST_0_i_9_n_0 ),
        .I3(\dout[11]_INST_0_i_10_n_0 ),
        .O(\dout[11]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \dout[11]_INST_0_i_30 
       (.I0(L[8]),
        .I1(\dout[9]_INST_0_i_11_n_0 ),
        .O(\dout[11]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \dout[11]_INST_0_i_31 
       (.I0(L[9]),
        .I1(\dout[9]_INST_0_i_14_n_0 ),
        .O(\dout[11]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h40405050CCCCFF00)) 
    \dout[11]_INST_0_i_32_rewire 
       (.I0(\addr[11]_INST_0_i_4_n_0 ),
        .I1(\addr[11]_INST_0_i_9_n_0 ),
        .I2(\addr[11]_INST_0_i_1_n_0 ),
        .I3(\dout[11]_INST_0_i_39_n_0 ),
        .I4(\dout[5]_INST_0_i_10_n_0 ),
        .I5(\FSM_sequential_state[1]_i_12_n_0 ),
        .O(\dout[11]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[11]_INST_0_i_33 
       (.I0(\rrd[0] [3]),
        .I1(\dout[14]_INST_0_i_25_n_0 ),
        .I2(pc[3]),
        .I3(eqOp93_in),
        .I4(data4[3]),
        .O(\dout[11]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88B8B8B8)) 
    \dout[11]_INST_0_i_34 
       (.I0(pc[11]),
        .I1(eqOp93_in),
        .I2(din[11]),
        .I3(r_a0),
        .I4(bw),
        .O(\dout[11]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB888B8BB)) 
    \dout[11]_INST_0_i_35 
       (.I0(\rrd[0] [1]),
        .I1(\dout[14]_INST_0_i_25_n_0 ),
        .I2(pc[1]),
        .I3(eqOp93_in),
        .I4(\dout[2]_INST_0_i_38_n_0 ),
        .O(\dout[11]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88B8B8B8)) 
    \dout[11]_INST_0_i_36 
       (.I0(pc[9]),
        .I1(eqOp93_in),
        .I2(din[9]),
        .I3(r_a0),
        .I4(bw),
        .O(\dout[11]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEFE0EFE0E0E0EF)) 
    \dout[11]_INST_0_i_37 
       (.I0(lbe_INST_0_i_7_n_0),
        .I1(\dout[11]_INST_0_i_40_n_0 ),
        .I2(\dout[14]_INST_0_i_25_n_0 ),
        .I3(\dout[11]_INST_0_i_41_n_0 ),
        .I4(eqOp93_in),
        .I5(pc[0]),
        .O(\dout[11]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88B8B8B8)) 
    \dout[11]_INST_0_i_38 
       (.I0(pc[8]),
        .I1(eqOp93_in),
        .I2(din[8]),
        .I3(r_a0),
        .I4(bw),
        .O(\dout[11]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000477777774777)) 
    \dout[11]_INST_0_i_39 
       (.I0(soc[2]),
        .I1(eqOp93_in),
        .I2(din[11]),
        .I3(\dout[15]_INST_0_i_109_n_0 ),
        .I4(\dout[5]_INST_0_i_14_n_0 ),
        .I5(src__0[11]),
        .O(\dout[11]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F444FFF44444444)) 
    \dout[11]_INST_0_i_4 
       (.I0(\dout[15]_INST_0_i_39_n_4 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_51_n_4 ),
        .I3(bw),
        .I4(\dout[15]_INST_0_i_56_n_4 ),
        .I5(\dout[15]_INST_0_i_20_n_0 ),
        .O(\dout[11]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA808A80808A80808)) 
    \dout[11]_INST_0_i_40 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(\dout[11]_INST_0_i_42_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(soc[0]),
        .I4(sr_reg_n_0_),
        .I5(\r_code[0]_i_1_n_0 ),
        .O(\dout[11]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h15D5)) 
    \dout[11]_INST_0_i_41 
       (.I0(din[0]),
        .I1(bw),
        .I2(r_a0),
        .I3(din[8]),
        .O(\dout[11]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dout[11]_INST_0_i_42 
       (.I0(sp_reg[0]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(pc[0]),
        .O(\dout[11]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h87877887B48778B4)) 
    \dout[11]_INST_0_i_5 
       (.I0(\dout[11]_INST_0_i_11_n_0 ),
        .I1(\dout[9]_INST_0_i_5_n_0 ),
        .I2(\dout[15]_INST_0_i_78_n_0 ),
        .I3(L[10]),
        .I4(\dout[2]_INST_0_i_12_n_0 ),
        .I5(\dout[11]_INST_0_i_14_n_0 ),
        .O(\dout[11]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFAFCF0FAFFFFF0FF)) 
    \dout[11]_INST_0_i_6 
       (.I0(\dout[14]_INST_0_i_10_n_0 ),
        .I1(\dout[14]_INST_0_i_11_n_0 ),
        .I2(\dout[11]_INST_0_i_15_n_0 ),
        .I3(\dout[11]_INST_0_i_16_n_0 ),
        .I4(L[11]),
        .I5(\dout[11]_INST_0_i_18_n_0 ),
        .O(\dout[11]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEEFE)) 
    \dout[11]_INST_0_i_7 
       (.I0(\dout[11]_INST_0_i_3_n_0 ),
        .I1(\dout[11]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_14_n_0 ),
        .I3(\dout[11]_INST_0_i_16_n_0 ),
        .O(\dout[11]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[11]_INST_0_i_8 
       (.CI(\dout[4]_INST_0_i_8_n_0 ),
        .CO({\dout[11]_INST_0_i_8_n_0 ,\dout[11]_INST_0_i_8_n_1 ,\dout[11]_INST_0_i_8_n_2 ,\dout[11]_INST_0_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(L[11:8]),
        .O({\dout[11]_INST_0_i_8_n_4 ,\dout[11]_INST_0_i_8_n_5 ,\dout[11]_INST_0_i_8_n_6 ,\dout[11]_INST_0_i_8_n_7 }),
        .S({\dout[11]_INST_0_i_22_n_0 ,\dout[11]_INST_0_i_23_n_0 ,\dout[11]_INST_0_i_24_n_0 ,\dout[11]_INST_0_i_25_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0030005000000050)) 
    \dout[11]_INST_0_i_9 
       (.I0(\dout[4]_INST_0_i_13_n_0 ),
        .I1(soc[1]),
        .I2(eqOp135_in),
        .I3(soc[2]),
        .I4(soc[0]),
        .I5(\dout[11]_INST_0_i_26_n_0 ),
        .O(\dout[11]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[12]_INST_0 
       (.I0(pc[12]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[12] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[12]_INST_0_i_1_n_0 ),
        .O(dout[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00A2)) 
    \dout[12]_INST_0_i_1 
       (.I0(\dout[12]_INST_0_i_2_n_0 ),
        .I1(\dout[13]_INST_0_i_3_n_0 ),
        .I2(\dout[12]_INST_0_i_3_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[12]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \dout[12]_INST_0_i_10 
       (.I0(\dout[15]_INST_0_i_20_n_0 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_21_n_7 ),
        .O(\dout[12]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABAAABBB)) 
    \dout[12]_INST_0_i_11 
       (.I0(\dout[15]_INST_0_i_37_n_0 ),
        .I1(\dout[4]_INST_0_i_13_n_0 ),
        .I2(din[12]),
        .I3(p_2_in88_in),
        .I4(r_code[12]),
        .O(\dout[12]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB800B800B800)) 
    \dout[12]_INST_0_i_12 
       (.I0(\dout[15]_INST_0_i_29_n_7 ),
        .I1(bw),
        .I2(\dout[15]_INST_0_i_30_n_7 ),
        .I3(\dout[15]_INST_0_i_31_n_0 ),
        .I4(\dout[4]_INST_0_i_7_n_0 ),
        .I5(\dout[15]_INST_0_i_28_n_7 ),
        .O(\dout[12]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF5510)) 
    \dout[12]_INST_0_i_2 
       (.I0(\dout[12]_INST_0_i_4_n_0 ),
        .I1(\dout[12]_INST_0_i_5_n_0 ),
        .I2(\dout[15]_INST_0_i_23_n_0 ),
        .I3(\dout[12]_INST_0_i_6_n_0 ),
        .I4(\dout[12]_INST_0_i_7_n_0 ),
        .O(\dout[12]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF8)) 
    \dout[12]_INST_0_i_3 
       (.I0(eqOp93_in),
        .I1(\dout[13]_INST_0_i_10_n_7 ),
        .I2(\dout[12]_INST_0_i_8_n_0 ),
        .I3(\dout[12]_INST_0_i_9_n_0 ),
        .O(\dout[12]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F444FFF44444444)) 
    \dout[12]_INST_0_i_4 
       (.I0(\dout[15]_INST_0_i_21_n_7 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_25_n_7 ),
        .I3(bw),
        .I4(\dout[15]_INST_0_i_26_n_7 ),
        .I5(\dout[15]_INST_0_i_20_n_0 ),
        .O(\dout[12]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h96)) 
    \dout[12]_INST_0_i_5 
       (.I0(\dout[9]_INST_0_i_5_n_0 ),
        .I1(L[12]),
        .I2(\dout[4]_INST_0_i_13_n_0 ),
        .O(\dout[12]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFAFCF0FAFFFFF0FF)) 
    \dout[12]_INST_0_i_6 
       (.I0(\dout[14]_INST_0_i_10_n_0 ),
        .I1(\dout[14]_INST_0_i_11_n_0 ),
        .I2(\dout[12]_INST_0_i_10_n_0 ),
        .I3(\dout[4]_INST_0_i_13_n_0 ),
        .I4(L[12]),
        .I5(\dout[12]_INST_0_i_11_n_0 ),
        .O(\dout[12]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEEFE)) 
    \dout[12]_INST_0_i_7 
       (.I0(\dout[12]_INST_0_i_3_n_0 ),
        .I1(\dout[12]_INST_0_i_12_n_0 ),
        .I2(\dout[15]_INST_0_i_14_n_0 ),
        .I3(\dout[4]_INST_0_i_13_n_0 ),
        .O(\dout[12]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h003000A0000000A0)) 
    \dout[12]_INST_0_i_8 
       (.I0(\dout[14]_INST_0_i_27_n_0 ),
        .I1(soc[1]),
        .I2(eqOp135_in),
        .I3(soc[2]),
        .I4(soc[0]),
        .I5(\dout[4]_INST_0_i_5_n_0 ),
        .O(\dout[12]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCC80CC8000000C00)) 
    \dout[12]_INST_0_i_9 
       (.I0(soc[0]),
        .I1(eqOp135_in),
        .I2(soc[1]),
        .I3(soc[2]),
        .I4(\dout[4]_INST_0_i_13_n_0 ),
        .I5(\dout[13]_INST_0_i_21_n_0 ),
        .O(\dout[12]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[13]_INST_0 
       (.I0(pc[13]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[13] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[13]_INST_0_i_1_n_0 ),
        .O(dout[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00A2)) 
    \dout[13]_INST_0_i_1 
       (.I0(\dout[13]_INST_0_i_2_n_0 ),
        .I1(\dout[13]_INST_0_i_3_n_0 ),
        .I2(\dout[13]_INST_0_i_4_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[13]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[13]_INST_0_i_10 
       (.CI(\dout[11]_INST_0_i_8_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,L[14:12]}),
        .O({\dout[13]_INST_0_i_10_n_4 ,\dout[13]_INST_0_i_10_n_5 ,\dout[13]_INST_0_i_10_n_6 ,\dout[13]_INST_0_i_10_n_7 }),
        .S({\dout[13]_INST_0_i_16_n_0 ,\dout[13]_INST_0_i_17_n_0 ,\dout[13]_INST_0_i_18_n_0 ,\dout[13]_INST_0_i_19_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0030005000000050)) 
    \dout[13]_INST_0_i_11 
       (.I0(\dout[14]_INST_0_i_9_n_0 ),
        .I1(soc[1]),
        .I2(eqOp135_in),
        .I3(soc[2]),
        .I4(soc[0]),
        .I5(\dout[13]_INST_0_i_20_n_0_repN ),
        .O(\dout[13]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCC880000C00000)) 
    \dout[13]_INST_0_i_12 
       (.I0(soc[0]),
        .I1(eqOp135_in),
        .I2(\dout[14]_INST_0_i_27_n_0 ),
        .I3(soc[1]),
        .I4(soc[2]),
        .I5(\dout[13]_INST_0_i_21_n_0 ),
        .O(\dout[13]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \dout[13]_INST_0_i_13 
       (.I0(\dout[15]_INST_0_i_20_n_0 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_21_n_6 ),
        .O(\dout[13]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \dout[13]_INST_0_i_14 
       (.I0(\dout[15]_INST_0_i_37_n_0 ),
        .I1(din[12]),
        .I2(p_2_in88_in),
        .I3(r_code[12]),
        .I4(\dout[14]_INST_0_i_27_n_0 ),
        .O(\dout[13]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFAC00AC00AC00)) 
    \dout[13]_INST_0_i_15 
       (.I0(\dout[15]_INST_0_i_29_n_6 ),
        .I1(\dout[15]_INST_0_i_30_n_6 ),
        .I2(bw),
        .I3(\dout[15]_INST_0_i_31_n_0 ),
        .I4(\dout[4]_INST_0_i_7_n_0 ),
        .I5(\dout[15]_INST_0_i_28_n_6 ),
        .O(\dout[13]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \dout[13]_INST_0_i_16 
       (.I0(L[15]),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[15]_INST_0_i_15_n_0 ),
        .O(\dout[13]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \dout[13]_INST_0_i_17 
       (.I0(L[14]),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[14]_INST_0_i_9_n_0 ),
        .O(\dout[13]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h9A)) 
    \dout[13]_INST_0_i_18 
       (.I0(L[13]),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[14]_INST_0_i_27_n_0 ),
        .O(\dout[13]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \dout[13]_INST_0_i_19 
       (.I0(L[12]),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[4]_INST_0_i_13_n_0 ),
        .O(\dout[13]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF5510)) 
    \dout[13]_INST_0_i_2 
       (.I0(\dout[13]_INST_0_i_5_n_0 ),
        .I1(\dout[13]_INST_0_i_6_n_0 ),
        .I2(\dout[15]_INST_0_i_23_n_0 ),
        .I3(\dout[13]_INST_0_i_7_n_0 ),
        .I4(\dout[13]_INST_0_i_8_n_0 ),
        .O(\dout[13]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0070)) 
    \dout[13]_INST_0_i_20_rewire_replica_rewire 
       (.I0(\dout[5]_INST_0_i_15_n_0 ),
        .I1(\dout[4]_INST_0_i_46_n_0 ),
        .I2(\dout[4]_INST_0_i_16_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[13]_INST_0_i_20_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h07)) 
    \dout[13]_INST_0_i_20_rewire_rewire_rewire 
       (.I0(\dout[5]_INST_0_i_15_n_0 ),
        .I1(\dout[4]_INST_0_i_46_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[13]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2220002000000000)) 
    \dout[13]_INST_0_i_21 
       (.I0(\dout[7]_INST_0_i_7_n_0_repN ),
        .I1(soc[2]),
        .I2(r_code[7]),
        .I3(p_2_in88_in),
        .I4(din[7]),
        .I5(soc[1]),
        .O(\dout[13]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h060095FF06FF9500)) 
    \dout[13]_INST_0_i_22 
       (.I0(p_1_in122_in),
        .I1(\sr_reg_n_0_[8] ),
        .I2(\r_code[11]_i_1_n_0 ),
        .I3(doc[0]),
        .I4(\r_code[10]_i_1_n_0 ),
        .I5(\dout[13]_INST_0_i_23_n_0 ),
        .O(\dout[13]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dout[13]_INST_0_i_23 
       (.I0(sr_reg_n_0_),
        .I1(\r_code[11]_i_1_n_0 ),
        .I2(\sr_reg_n_0_[1] ),
        .O(\dout[13]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00053305)) 
    \dout[13]_INST_0_i_3 
       (.I0(r_code[15]),
        .I1(din[15]),
        .I2(r_code[14]),
        .I3(p_2_in88_in),
        .I4(din[14]),
        .O(\dout[13]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF8)) 
    \dout[13]_INST_0_i_4 
       (.I0(eqOp93_in),
        .I1(\dout[13]_INST_0_i_10_n_6 ),
        .I2(\dout[13]_INST_0_i_11_n_0 ),
        .I3(\dout[13]_INST_0_i_12_n_0 ),
        .O(\dout[13]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F444FFF44444444)) 
    \dout[13]_INST_0_i_5 
       (.I0(\dout[15]_INST_0_i_21_n_6 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_25_n_6 ),
        .I3(bw),
        .I4(\dout[15]_INST_0_i_26_n_6 ),
        .I5(\dout[15]_INST_0_i_20_n_0 ),
        .O(\dout[13]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAEA7E57AAAAAAEA)) 
    \dout[13]_INST_0_i_6 
       (.I0(\dout[14]_INST_0_i_29_n_0_repN ),
        .I1(\dout[14]_INST_0_i_19_n_0 ),
        .I2(\dout[14]_INST_0_i_9_n_0 ),
        .I3(L[14]),
        .I4(L[15]),
        .I5(\dout[15]_INST_0_i_15_n_0 ),
        .O(\dout[13]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFAFAF0FFFFFFF0)) 
    \dout[13]_INST_0_i_7 
       (.I0(\dout[14]_INST_0_i_10_n_0 ),
        .I1(\dout[14]_INST_0_i_11_n_0 ),
        .I2(\dout[13]_INST_0_i_13_n_0 ),
        .I3(L[13]),
        .I4(\dout[14]_INST_0_i_27_n_0 ),
        .I5(\dout[13]_INST_0_i_14_n_0 ),
        .O(\dout[13]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFEEE)) 
    \dout[13]_INST_0_i_8 
       (.I0(\dout[13]_INST_0_i_4_n_0 ),
        .I1(\dout[13]_INST_0_i_15_n_0 ),
        .I2(\dout[14]_INST_0_i_27_n_0 ),
        .I3(\dout[15]_INST_0_i_14_n_0 ),
        .O(\dout[13]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \dout[13]_INST_0_i_9 
       (.I0(r_code[13]),
        .I1(p_2_in88_in),
        .I2(din[13]),
        .I3(\dout[13]_INST_0_i_3_n_0 ),
        .O(eqOp93_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[14]_INST_0 
       (.I0(pc[14]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[14] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[14]_INST_0_i_1_n_0 ),
        .O(dout[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AAFE)) 
    \dout[14]_INST_0_i_1 
       (.I0(\dout[14]_INST_0_i_2_n_0 ),
        .I1(\dout[14]_INST_0_i_3_n_0 ),
        .I2(\dout[14]_INST_0_i_4_n_0 ),
        .I3(\dout[14]_INST_0_i_5_n_0 ),
        .I4(\dout[14]_INST_0_i_6_n_0 ),
        .I5(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[14]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000B80000000000)) 
    \dout[14]_INST_0_i_10 
       (.I0(din[14]),
        .I1(p_2_in88_in),
        .I2(r_code[14]),
        .I3(doc[3]),
        .I4(doc[0]),
        .I5(doc[1]),
        .O(\dout[14]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB830880000000000)) 
    \dout[14]_INST_0_i_11 
       (.I0(din[13]),
        .I1(p_2_in88_in),
        .I2(r_code[13]),
        .I3(din[15]),
        .I4(r_code[15]),
        .I5(doc[0]),
        .O(\dout[14]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \dout[14]_INST_0_i_12 
       (.I0(\dout[15]_INST_0_i_20_n_0 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_21_n_5 ),
        .O(\dout[14]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[14]_INST_0_i_13 
       (.I0(\dout[14]_INST_0_i_23_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\rrd[0] [14]),
        .I3(\dout[14]_INST_0_i_25_n_0 ),
        .I4(\dout[14]_INST_0_i_26_n_0 ),
        .O(L[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABAAABBB)) 
    \dout[14]_INST_0_i_14 
       (.I0(\dout[15]_INST_0_i_37_n_0 ),
        .I1(\dout[14]_INST_0_i_9_n_0 ),
        .I2(din[12]),
        .I3(p_2_in88_in),
        .I4(r_code[12]),
        .O(\dout[14]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[14]_INST_0_i_15 
       (.I0(L[14]),
        .I1(\dout[14]_INST_0_i_9_n_0 ),
        .O(\dout[15]_INST_0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \dout[14]_INST_0_i_16 
       (.I0(\dout[14]_INST_0_i_27_n_0 ),
        .I1(L[13]),
        .O(\dout[14]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hDF5D)) 
    \dout[14]_INST_0_i_17 
       (.I0(\dout[15]_INST_0_i_45_n_0 ),
        .I1(L[12]),
        .I2(\dout[4]_INST_0_i_13_n_0 ),
        .I3(\dout[9]_INST_0_i_5_n_0 ),
        .O(\dout[14]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h220202002B222202)) 
    \dout[14]_INST_0_i_18 
       (.I0(\dout[15]_INST_0_i_15_n_0 ),
        .I1(L[15]),
        .I2(L[14]),
        .I3(\dout[14]_INST_0_i_9_n_0 ),
        .I4(\dout[14]_INST_0_i_19_n_0 ),
        .I5(\dout[14]_INST_0_i_29_n_0 ),
        .O(\dout[14]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "dout[14]_INST_0_i_18" *) 
  LUT6 #(
    .INIT(64'h220202002B222202)) 
    \dout[14]_INST_0_i_18_replica 
       (.I0(\dout[15]_INST_0_i_15_n_0 ),
        .I1(L[15]),
        .I2(L[14]),
        .I3(\dout[14]_INST_0_i_9_n_0 ),
        .I4(\dout[14]_INST_0_i_19_n_0 ),
        .I5(\dout[14]_INST_0_i_29_n_0 ),
        .O(\dout[14]_INST_0_i_18_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h004D4DFF)) 
    \dout[14]_INST_0_i_19 
       (.I0(\dout[9]_INST_0_i_5_n_0 ),
        .I1(\dout[4]_INST_0_i_13_n_0 ),
        .I2(L[12]),
        .I3(L[13]),
        .I4(\dout[14]_INST_0_i_27_n_0 ),
        .O(\dout[14]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEEFE)) 
    \dout[14]_INST_0_i_2 
       (.I0(\dout[14]_INST_0_i_7_n_0 ),
        .I1(\dout[14]_INST_0_i_8_n_0 ),
        .I2(\dout[15]_INST_0_i_14_n_0 ),
        .I3(\dout[14]_INST_0_i_9_n_0 ),
        .O(\dout[14]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0030005000000050)) 
    \dout[14]_INST_0_i_20 
       (.I0(\dout[15]_INST_0_i_15_n_0 ),
        .I1(soc[1]),
        .I2(eqOp135_in),
        .I3(soc[2]),
        .I4(soc[0]),
        .I5(\dout[6]_INST_0_i_7_n_0_repN ),
        .O(\dout[14]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h337F337FFFFFF3FF))
    \dout[14]_INST_0_i_21 
       (.I0(soc[0]),
        .I1(eqOp135_in),
        .I2(soc[1]),
        .I3(soc[2]),
        .I4(\dout[14]_INST_0_i_9_n_0 ),
        .I5(\dout[13]_INST_0_i_21_n_0 ),
        .O(\dout[14]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44CC55F0)) 
    \dout[14]_INST_0_i_22 
       (.I0(\addr[14]_INST_0_i_9_n_0 ),
        .I1(\addr[14]_INST_0_i_1_n_0 ),
        .I2(\dout[14]_INST_0_i_30_n_0 ),
        .I3(\dout[5]_INST_0_i_10_n_0 ),
        .I4(\FSM_sequential_state[1]_i_12_n_0 ),
        .O(\dout[14]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[14]_INST_0_i_23 
       (.I0(\rrd[0] [6]),
        .I1(\dout[14]_INST_0_i_25_n_0 ),
        .I2(pc[6]),
        .I3(eqOp93_in),
        .I4(data4[6]),
        .O(\dout[14]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEAEAEAFF)) 
    \dout[14]_INST_0_i_24 
       (.I0(\addr[14]_INST_0_i_7_n_0 ),
        .I1(\addr[15]_INST_0_i_11_n_0 ),
        .I2(\dout[14]_INST_0_i_31_n_0 ),
        .I3(\r_code[3]_i_1_n_0 ),
        .I4(\addr[14]_INST_0_i_3_n_0 ),
        .O(\rrd[0] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA8A8AAAA08A80)) 
    \dout[14]_INST_0_i_25 
       (.I0(rd_INST_0_i_16_n_0),
        .I1(din[14]),
        .I2(p_2_in88_in),
        .I3(r_code[14]),
        .I4(din[15]),
        .I5(r_code[15]),
        .O(\dout[14]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88B8B8B8)) 
    \dout[14]_INST_0_i_26 
       (.I0(pc[14]),
        .I1(eqOp93_in),
        .I2(din[14]),
        .I3(r_a0),
        .I4(bw),
        .O(\dout[14]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h07000F0F)) 
    \dout[14]_INST_0_i_27_rewire_rewire 
       (.I0(\dout[5]_INST_0_i_15_n_0 ),
        .I1(\dout[4]_INST_0_i_46_n_0 ),
        .I2(\dout[14]_INST_0_i_32_n_0 ),
        .I3(\dout[4]_INST_0_i_16_n_0 ),
        .I4(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[14]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[14]_INST_0_i_28 
       (.I0(L[13]),
        .I1(\dout[14]_INST_0_i_27_n_0 ),
        .O(\dout[15]_INST_0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9A59)) 
    \dout[14]_INST_0_i_29 
       (.I0(\dout[15]_INST_0_i_45_n_0 ),
        .I1(L[12]),
        .I2(\dout[4]_INST_0_i_13_n_0 ),
        .I3(\dout[9]_INST_0_i_5_n_0 ),
        .O(\dout[14]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "dout[14]_INST_0_i_29" *) 
  LUT4 #(
    .INIT(16'h9A59)) 
    \dout[14]_INST_0_i_29_replica 
       (.I0(\dout[15]_INST_0_i_45_n_0 ),
        .I1(L[12]),
        .I2(\dout[4]_INST_0_i_13_n_0 ),
        .I3(\dout[9]_INST_0_i_5_n_0 ),
        .O(\dout[14]_INST_0_i_29_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFAF0FCFAFFF0FFFF)) 
    \dout[14]_INST_0_i_3 
       (.I0(\dout[14]_INST_0_i_10_n_0 ),
        .I1(\dout[14]_INST_0_i_11_n_0 ),
        .I2(\dout[14]_INST_0_i_12_n_0 ),
        .I3(L[14]),
        .I4(\dout[14]_INST_0_i_9_n_0 ),
        .I5(\dout[14]_INST_0_i_14_n_0 ),
        .O(\dout[14]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000477777774777)) 
    \dout[14]_INST_0_i_30 
       (.I0(soc[2]),
        .I1(eqOp93_in),
        .I2(din[14]),
        .I3(\dout[15]_INST_0_i_109_n_0 ),
        .I4(\dout[5]_INST_0_i_14_n_0 ),
        .I5(src__0[14]),
        .O(\dout[14]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF454045404540)) 
    \dout[14]_INST_0_i_31 
       (.I0(\r_code[1]_i_1_n_0 ),
        .I1(sp_reg[14]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(pc[14]),
        .I4(\addr[3]_INST_0_i_47_n_0 ),
        .I5(\sr_reg_n_0_[14] ),
        .O(\dout[14]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1101330311013000)) 
    \dout[14]_INST_0_i_32 
       (.I0(\rrs[0] [13]),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\dout[5]_INST_0_i_10_n_0 ),
        .I3(\addr[13]_INST_0_i_8_n_0 ),
        .I4(\FSM_sequential_state[1]_i_12_n_0 ),
        .I5(\dout[14]_INST_0_i_33_n_0 ),
        .O(\dout[14]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000477777774777)) 
    \dout[14]_INST_0_i_33 
       (.I0(soc[2]),
        .I1(eqOp93_in),
        .I2(din[13]),
        .I3(\dout[15]_INST_0_i_109_n_0 ),
        .I4(\dout[5]_INST_0_i_14_n_0 ),
        .I5(src__0[13]),
        .O(\dout[14]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5569AA6900000000)) 
    \dout[14]_INST_0_i_4 
       (.I0(\dout[15]_INST_0_i_44_n_0 ),
        .I1(\dout[14]_INST_0_i_16_n_0 ),
        .I2(\dout[14]_INST_0_i_17_n_0 ),
        .I3(\dout[14]_INST_0_i_18_n_0_repN ),
        .I4(\dout[14]_INST_0_i_19_n_0 ),
        .I5(\dout[15]_INST_0_i_23_n_0 ),
        .O(\dout[14]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F444FFF44444444)) 
    \dout[14]_INST_0_i_5 
       (.I0(\dout[15]_INST_0_i_21_n_5 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_25_n_5 ),
        .I3(bw),
        .I4(\dout[15]_INST_0_i_26_n_5 ),
        .I5(\dout[15]_INST_0_i_20_n_0 ),
        .O(\dout[14]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000440347)) 
    \dout[14]_INST_0_i_6 
       (.I0(din[14]),
        .I1(p_2_in88_in),
        .I2(r_code[14]),
        .I3(din[15]),
        .I4(r_code[15]),
        .I5(\dout[14]_INST_0_i_7_n_0 ),
        .O(\dout[14]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF8)) 
    \dout[14]_INST_0_i_7 
       (.I0(eqOp93_in),
        .I1(\dout[13]_INST_0_i_10_n_5 ),
        .I2(\dout[14]_INST_0_i_20_n_0 ),
        .I3(\dout[14]_INST_0_i_21_n_0 ),
        .O(\dout[14]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB800B800B800)) 
    \dout[14]_INST_0_i_8 
       (.I0(\dout[15]_INST_0_i_29_n_5 ),
        .I1(bw),
        .I2(\dout[15]_INST_0_i_30_n_5 ),
        .I3(\dout[15]_INST_0_i_31_n_0 ),
        .I4(\dout[4]_INST_0_i_7_n_0 ),
        .I5(\dout[15]_INST_0_i_28_n_5 ),
        .O(\dout[14]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACFC)) 
    \dout[14]_INST_0_i_9_rewire 
       (.I0(\dout[5]_INST_0_i_11_n_0 ),
        .I1(\dout[14]_INST_0_i_22_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .I3(\dout[5]_INST_0_i_5_n_0 ),
        .O(\dout[14]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[15]_INST_0 
       (.I0(pc[15]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[15] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[15]_INST_0_i_3_n_0 ),
        .O(dout[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0009000800080008)) 
    \dout[15]_INST_0_i_1 
       (.I0(state[2]),
        .I1(state[3]),
        .I2(state[4]),
        .I3(\dout[15]_INST_0_i_4_n_0 ),
        .I4(soc[0]),
        .I5(nstate1),
        .O(\dout[15]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000440347)) 
    \dout[15]_INST_0_i_10 
       (.I0(din[14]),
        .I1(p_2_in88_in),
        .I2(r_code[14]),
        .I3(din[15]),
        .I4(r_code[15]),
        .I5(\dout[15]_INST_0_i_12_n_0 ),
        .O(\dout[15]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \dout[15]_INST_0_i_100 
       (.I0(\dout[9]_INST_0_i_11_n_0 ),
        .O(\dout[15]_INST_0_i_100_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_101 
       (.I0(L[11]),
        .I1(\dout[11]_INST_0_i_16_n_0 ),
        .O(\dout[15]_INST_0_i_101_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_102 
       (.I0(L[10]),
        .I1(\dout[2]_INST_0_i_12_n_0 ),
        .O(\dout[15]_INST_0_i_102_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_103 
       (.I0(L[9]),
        .I1(\dout[9]_INST_0_i_14_n_0 ),
        .O(\dout[15]_INST_0_i_103_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[15]_INST_0_i_104 
       (.I0(L[8]),
        .I1(sr_reg_n_0_),
        .O(\dout[15]_INST_0_i_104_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \dout[15]_INST_0_i_109 
       (.I0(bw),
        .I1(r_a0),
        .O(\dout[15]_INST_0_i_109_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h22222222222222A2)) 
    \dout[15]_INST_0_i_11 
       (.I0(bw),
        .I1(\dout[13]_INST_0_i_3_n_0 ),
        .I2(doc[0]),
        .I3(doc[1]),
        .I4(\r_code[11]_i_1_n_0 ),
        .I5(\r_code[10]_i_1_n_0 ),
        .O(\dout[15]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFF080808)) 
    \dout[15]_INST_0_i_12 
       (.I0(\dout[6]_INST_0_i_5_n_0 ),
        .I1(sr_reg_n_0_),
        .I2(soc[1]),
        .I3(\dout[13]_INST_0_i_10_n_4 ),
        .I4(eqOp93_in),
        .I5(\dout[15]_INST_0_i_27_n_0 ),
        .O(\dout[15]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8FFF88888888888)) 
    \dout[15]_INST_0_i_13 
       (.I0(p_13_in),
        .I1(\dout[4]_INST_0_i_7_n_0 ),
        .I2(\dout[15]_INST_0_i_29_n_4 ),
        .I3(bw),
        .I4(\dout[15]_INST_0_i_30_n_4 ),
        .I5(\dout[15]_INST_0_i_31_n_0 ),
        .O(\dout[15]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0044034700000000)) 
    \dout[15]_INST_0_i_14 
       (.I0(din[12]),
        .I1(p_2_in88_in),
        .I2(r_code[12]),
        .I3(din[13]),
        .I4(r_code[13]),
        .I5(\dout[15]_INST_0_i_32_n_0 ),
        .O(\dout[15]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h74)) 
    \dout[15]_INST_0_i_15 
       (.I0(\dout[15]_INST_0_i_33_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\dout[15]_INST_0_i_34_n_0 ),
        .O(\dout[15]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h74)) 
    \dout[15]_INST_0_i_16 
       (.I0(\dout[15]_INST_0_i_43_n_0 ),
        .I1(\dout[14]_INST_0_i_10_n_0 ),
        .I2(\dout[15]_INST_0_i_36_n_0 ),
        .O(\dout[15]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8880888888808080)) 
    \dout[15]_INST_0_i_17 
       (.I0(doc[1]),
        .I1(doc[3]),
        .I2(doc[0]),
        .I3(din[14]),
        .I4(p_2_in88_in),
        .I5(r_code[14]),
        .O(\dout[15]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000FFE2)) 
    \dout[15]_INST_0_i_18 
       (.I0(r_code[12]),
        .I1(p_2_in88_in),
        .I2(din[12]),
        .I3(\dout[15]_INST_0_i_15_n_0 ),
        .I4(\dout[15]_INST_0_i_37_n_0 ),
        .I5(\dout[15]_INST_0_i_38_n_0 ),
        .O(\dout[15]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000C0000000C0A0A)) 
    \dout[15]_INST_0_i_19 
       (.I0(r_code[15]),
        .I1(din[15]),
        .I2(doc[1]),
        .I3(din[14]),
        .I4(p_2_in88_in),
        .I5(r_code[14]),
        .O(\dout[15]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010000)) 
    \dout[15]_INST_0_i_2 
       (.I0(state[2]),
        .I1(state[3]),
        .I2(state[0]),
        .I3(state[1]),
        .I4(state[4]),
        .O(\dout[15]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB830880000000000)) 
    \dout[15]_INST_0_i_20 
       (.I0(din[12]),
        .I1(p_2_in88_in),
        .I2(r_code[12]),
        .I3(din[13]),
        .I4(r_code[13]),
        .I5(\dout[15]_INST_0_i_32_n_0 ),
        .O(\dout[15]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[15]_INST_0_i_21 
       (.CI(\dout[15]_INST_0_i_39_n_0 ),
        .CO({\dout[15]_INST_0_i_21_n_0 ,\dout[15]_INST_0_i_21_n_1 ,\dout[15]_INST_0_i_21_n_2 ,\dout[15]_INST_0_i_21_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(L[15:12]),
        .O({\dout[15]_INST_0_i_21_n_4 ,\dout[15]_INST_0_i_21_n_5 ,\dout[15]_INST_0_i_21_n_6 ,\dout[15]_INST_0_i_21_n_7 }),
        .S({\dout[15]_INST_0_i_43_n_0 ,\dout[15]_INST_0_i_44_n_0 ,\dout[15]_INST_0_i_45_n_0 ,\dout[15]_INST_0_i_46_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3CC33DC3C13CED3E)) 
    \dout[15]_INST_0_i_22 
       (.I0(\dout[15]_INST_0_i_47_n_0 ),
        .I1(\dout[15]_INST_0_i_48_n_0 ),
        .I2(L[15]),
        .I3(\dout[15]_INST_0_i_15_n_0 ),
        .I4(\dout[15]_INST_0_i_49_n_0 ),
        .I5(\dout[15]_INST_0_i_50_n_0 ),
        .O(\dout[15]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0008000000080808)) 
    \dout[15]_INST_0_i_23 
       (.I0(doc[1]),
        .I1(doc[3]),
        .I2(doc[0]),
        .I3(din[14]),
        .I4(p_2_in88_in),
        .I5(r_code[14]),
        .O(\dout[15]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000101000051015)) 
    \dout[15]_INST_0_i_24 
       (.I0(\dout[15]_INST_0_i_21_n_4 ),
        .I1(din[13]),
        .I2(p_2_in88_in),
        .I3(r_code[13]),
        .I4(din[14]),
        .I5(r_code[14]),
        .O(\dout[15]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[15]_INST_0_i_25 
       (.CI(\dout[15]_INST_0_i_51_n_0 ),
        .CO({\dout[15]_INST_0_i_25_n_0 ,\dout[15]_INST_0_i_25_n_1 ,\dout[15]_INST_0_i_25_n_2 ,\dout[15]_INST_0_i_25_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(L[15:12]),
        .O({\dout[15]_INST_0_i_25_n_4 ,\dout[15]_INST_0_i_25_n_5 ,\dout[15]_INST_0_i_25_n_6 ,\dout[15]_INST_0_i_25_n_7 }),
        .S({\dout[15]_INST_0_i_43_n_0 ,\dout[15]_INST_0_i_44_n_0 ,\dout[15]_INST_0_i_45_n_0 ,\dout[15]_INST_0_i_55_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[15]_INST_0_i_26 
       (.CI(\dout[15]_INST_0_i_56_n_0 ),
        .CO({\dout[15]_INST_0_i_26_n_0 ,\dout[15]_INST_0_i_26_n_1 ,\dout[15]_INST_0_i_26_n_2 ,\dout[15]_INST_0_i_26_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(L[15:12]),
        .O({\dout[15]_INST_0_i_26_n_4 ,\dout[15]_INST_0_i_26_n_5 ,\dout[15]_INST_0_i_26_n_6 ,\dout[15]_INST_0_i_26_n_7 }),
        .S({\dout[15]_INST_0_i_43_n_0 ,\dout[15]_INST_0_i_44_n_0 ,\dout[15]_INST_0_i_45_n_0 ,\dout[15]_INST_0_i_60_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h11F4000011040000)) 
    \dout[15]_INST_0_i_27 
       (.I0(\dout[15]_INST_0_i_15_n_0 ),
        .I1(soc[1]),
        .I2(soc[0]),
        .I3(soc[2]),
        .I4(eqOp135_in),
        .I5(\dout[7]_INST_0_i_7_n_0_repN ),
        .O(\dout[15]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[15]_INST_0_i_28 
       (.CI(\dout[15]_INST_0_i_61_n_0 ),
        .CO({\dout[15]_INST_0_i_28_n_0 ,\dout[15]_INST_0_i_28_n_1 ,\dout[15]_INST_0_i_28_n_2 ,\dout[15]_INST_0_i_28_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(L[15:12]),
        .O({p_13_in,\dout[15]_INST_0_i_28_n_5 ,\dout[15]_INST_0_i_28_n_6 ,\dout[15]_INST_0_i_28_n_7 }),
        .S({\dout[15]_INST_0_i_62_n_0 ,\dout[15]_INST_0_i_63_n_0 ,\dout[15]_INST_0_i_64_n_0 ,\dout[15]_INST_0_i_65_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[15]_INST_0_i_29 
       (.CI(\dout[15]_INST_0_i_66_n_0 ),
        .CO({\dout[15]_INST_0_i_29_n_0 ,\dout[15]_INST_0_i_29_n_1 ,\dout[15]_INST_0_i_29_n_2 ,\dout[15]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(L[15:12]),
        .O({\dout[15]_INST_0_i_29_n_4 ,\dout[15]_INST_0_i_29_n_5 ,\dout[15]_INST_0_i_29_n_6 ,\dout[15]_INST_0_i_29_n_7 }),
        .S({\dout[15]_INST_0_i_67_n_0 ,\dout[15]_INST_0_i_68_n_0 ,\dout[15]_INST_0_i_69_n_0 ,\dout[15]_INST_0_i_70_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AAFE)) 
    \dout[15]_INST_0_i_3 
       (.I0(\dout[15]_INST_0_i_6_n_0 ),
        .I1(\dout[15]_INST_0_i_7_n_0 ),
        .I2(\dout[15]_INST_0_i_8_n_0 ),
        .I3(\dout[15]_INST_0_i_9_n_0 ),
        .I4(\dout[15]_INST_0_i_10_n_0 ),
        .I5(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[15]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[15]_INST_0_i_30 
       (.CI(\dout[15]_INST_0_i_71_n_0 ),
        .CO({\dout[15]_INST_0_i_30_n_0 ,\dout[15]_INST_0_i_30_n_1 ,\dout[15]_INST_0_i_30_n_2 ,\dout[15]_INST_0_i_30_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\dout[15]_INST_0_i_30_n_4 ,\dout[15]_INST_0_i_30_n_5 ,\dout[15]_INST_0_i_30_n_6 ,\dout[15]_INST_0_i_30_n_7 }),
        .S({p_13_in,\dout[15]_INST_0_i_28_n_5 ,\dout[15]_INST_0_i_28_n_6 ,\dout[15]_INST_0_i_28_n_7 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4703440000000000)) 
    \dout[15]_INST_0_i_31 
       (.I0(din[12]),
        .I1(p_2_in88_in),
        .I2(r_code[12]),
        .I3(din[13]),
        .I4(r_code[13]),
        .I5(\dout[15]_INST_0_i_32_n_0 ),
        .O(\dout[15]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000ACC0A)) 
    \dout[15]_INST_0_i_32 
       (.I0(r_code[14]),
        .I1(din[14]),
        .I2(r_code[15]),
        .I3(p_2_in88_in),
        .I4(din[15]),
        .O(\dout[15]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000EFEFEF)) 
    \dout[15]_INST_0_i_33_rewire 
       (.I0(\addr[7]_INST_0_i_5_n_0 ),
        .I1(\rrs[0] [7]),
        .I2(\FSM_sequential_state[1]_i_12_n_0 ),
        .I3(\addr[7]_INST_0_i_8_n_0 ),
        .I4(\dout[5]_INST_0_i_10_n_0 ),
        .I5(\dout[15]_INST_0_i_76_n_0 ),
        .O(\dout[15]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4455CCF0)) 
    \dout[15]_INST_0_i_34 
       (.I0(\addr[15]_INST_0_i_2_n_0 ),
        .I1(\addr[15]_INST_0_i_16_n_0 ),
        .I2(\dout[15]_INST_0_i_77_n_0 ),
        .I3(\dout[5]_INST_0_i_10_n_0 ),
        .I4(\FSM_sequential_state[1]_i_12_n_0 ),
        .O(\dout[15]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[15]_INST_0_i_35 
       (.I0(L[15]),
        .I1(\dout[15]_INST_0_i_15_n_0 ),
        .O(\dout[15]_INST_0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[15]_INST_0_i_36 
       (.I0(L[15]),
        .I1(\dout[15]_INST_0_i_15_n_0 ),
        .O(\dout[15]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF3FFF5F5F3FFFFFF)) 
    \dout[15]_INST_0_i_37 
       (.I0(r_code[15]),
        .I1(din[15]),
        .I2(doc[1]),
        .I3(din[14]),
        .I4(p_2_in88_in),
        .I5(r_code[14]),
        .O(\dout[15]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[15]_INST_0_i_38 
       (.I0(\dout[15]_INST_0_i_15_n_0 ),
        .I1(L[15]),
        .O(\dout[15]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[15]_INST_0_i_39 
       (.CI(\dout[4]_INST_0_i_11_n_0 ),
        .CO({\dout[15]_INST_0_i_39_n_0 ,\dout[15]_INST_0_i_39_n_1 ,\dout[15]_INST_0_i_39_n_2 ,\dout[15]_INST_0_i_39_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(L[11:8]),
        .O({\dout[15]_INST_0_i_39_n_4 ,\dout[15]_INST_0_i_39_n_5 ,\dout[15]_INST_0_i_39_n_6 ,\dout[15]_INST_0_i_39_n_7 }),
        .S({\dout[15]_INST_0_i_78_n_0 ,\dout[15]_INST_0_i_79_n_0 ,\dout[15]_INST_0_i_80_n_0 ,\dout[15]_INST_0_i_81_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \dout[15]_INST_0_i_4 
       (.I0(state[0]),
        .I1(state[1]),
        .O(\dout[15]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[15]_INST_0_i_40 
       (.I0(\dout[15]_INST_0_i_82_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\addr[15]_INST_0_i_62_n_0 ),
        .I3(\dout[14]_INST_0_i_25_n_0 ),
        .I4(\dout[15]_INST_0_i_83_n_0 ),
        .O(L[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[15]_INST_0_i_41 
       (.I0(\dout[15]_INST_0_i_84_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\rrd[0] [13]),
        .I3(\dout[14]_INST_0_i_25_n_0 ),
        .I4(\dout[15]_INST_0_i_85_n_0 ),
        .O(L[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[15]_INST_0_i_42 
       (.I0(\dout[4]_INST_0_i_34_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\rrd[0] [12]),
        .I3(\dout[14]_INST_0_i_25_n_0 ),
        .I4(\dout[15]_INST_0_i_86_n_0 ),
        .O(L[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[15]_INST_0_i_46 
       (.I0(L[12]),
        .I1(\dout[4]_INST_0_i_13_n_0 ),
        .O(\dout[15]_INST_0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF17117717)) 
    \dout[15]_INST_0_i_47 
       (.I0(\dout[14]_INST_0_i_27_n_0 ),
        .I1(L[13]),
        .I2(L[12]),
        .I3(\dout[4]_INST_0_i_13_n_0 ),
        .I4(\dout[9]_INST_0_i_5_n_0 ),
        .I5(\dout[15]_INST_0_i_87_n_0 ),
        .O(\dout[15]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[15]_INST_0_i_48 
       (.I0(L[14]),
        .I1(\dout[14]_INST_0_i_9_n_0 ),
        .O(\dout[15]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFB2B24D4DFF)) 
    \dout[15]_INST_0_i_49 
       (.I0(\dout[9]_INST_0_i_5_n_0 ),
        .I1(\dout[4]_INST_0_i_13_n_0 ),
        .I2(L[12]),
        .I3(L[13]),
        .I4(\dout[14]_INST_0_i_27_n_0 ),
        .I5(\dout[15]_INST_0_i_44_n_0 ),
        .O(\dout[15]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[15]_INST_0_i_5 
       (.I0(soc[2]),
        .I1(soc[1]),
        .O(nstate1));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDF5D0000FFFFDF5D)) 
    \dout[15]_INST_0_i_50 
       (.I0(\dout[15]_INST_0_i_45_n_0 ),
        .I1(L[12]),
        .I2(\dout[4]_INST_0_i_13_n_0 ),
        .I3(\dout[9]_INST_0_i_5_n_0 ),
        .I4(\dout[14]_INST_0_i_16_n_0 ),
        .I5(\dout[15]_INST_0_i_44_n_0 ),
        .O(\dout[15]_INST_0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[15]_INST_0_i_51 
       (.CI(\<const0>__0__0 ),
        .CO({\dout[15]_INST_0_i_51_n_0 ,\dout[15]_INST_0_i_51_n_1 ,\dout[15]_INST_0_i_51_n_2 ,\dout[15]_INST_0_i_51_n_3 }),
        .CYINIT(\dout[9]_INST_0_i_11_n_0 ),
        .DI(L[11:8]),
        .O({\dout[15]_INST_0_i_51_n_4 ,\dout[15]_INST_0_i_51_n_5 ,\dout[15]_INST_0_i_51_n_6 ,\dout[15]_INST_0_i_51_n_7 }),
        .S({\dout[15]_INST_0_i_78_n_0 ,\dout[15]_INST_0_i_79_n_0 ,\dout[15]_INST_0_i_80_n_0_repN ,\dout[15]_INST_0_i_91_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[15]_INST_0_i_55 
       (.I0(L[12]),
        .I1(\dout[4]_INST_0_i_13_n_0 ),
        .O(\dout[15]_INST_0_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[15]_INST_0_i_56 
       (.CI(\dout[4]_INST_0_i_43_n_0 ),
        .CO({\dout[15]_INST_0_i_56_n_0 ,\dout[15]_INST_0_i_56_n_1 ,\dout[15]_INST_0_i_56_n_2 ,\dout[15]_INST_0_i_56_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(L[11:8]),
        .O({\dout[15]_INST_0_i_56_n_4 ,\dout[15]_INST_0_i_56_n_5 ,\dout[15]_INST_0_i_56_n_6 ,\dout[15]_INST_0_i_56_n_7 }),
        .S({\dout[15]_INST_0_i_78_n_0 ,\dout[15]_INST_0_i_79_n_0 ,\dout[15]_INST_0_i_80_n_0 ,\dout[15]_INST_0_i_95_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEEFE)) 
    \dout[15]_INST_0_i_6 
       (.I0(\dout[15]_INST_0_i_12_n_0 ),
        .I1(\dout[15]_INST_0_i_13_n_0 ),
        .I2(\dout[15]_INST_0_i_14_n_0 ),
        .I3(\dout[15]_INST_0_i_15_n_0 ),
        .O(\dout[15]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[15]_INST_0_i_60 
       (.I0(L[12]),
        .I1(\dout[4]_INST_0_i_13_n_0 ),
        .O(\dout[15]_INST_0_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[15]_INST_0_i_61 
       (.CI(\dout[4]_INST_0_i_6_n_0 ),
        .CO({\dout[15]_INST_0_i_61_n_0 ,\dout[15]_INST_0_i_61_n_1 ,\dout[15]_INST_0_i_61_n_2 ,\dout[15]_INST_0_i_61_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(L[11:8]),
        .O({\dout[15]_INST_0_i_61_n_4 ,\dout[15]_INST_0_i_61_n_5 ,\dout[15]_INST_0_i_61_n_6 ,\dout[15]_INST_0_i_61_n_7 }),
        .S({\dout[15]_INST_0_i_96_n_0 ,\dout[15]_INST_0_i_97_n_0 ,\dout[15]_INST_0_i_98_n_0 ,\dout[15]_INST_0_i_99_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_62 
       (.I0(L[15]),
        .I1(\dout[15]_INST_0_i_15_n_0 ),
        .O(\dout[15]_INST_0_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_63 
       (.I0(L[14]),
        .I1(\dout[14]_INST_0_i_9_n_0 ),
        .O(\dout[15]_INST_0_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[15]_INST_0_i_64 
       (.I0(L[13]),
        .I1(\dout[14]_INST_0_i_27_n_0 ),
        .O(\dout[15]_INST_0_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_65 
       (.I0(L[12]),
        .I1(\dout[4]_INST_0_i_13_n_0 ),
        .O(\dout[15]_INST_0_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[15]_INST_0_i_66 
       (.CI(\<const0>__0__0 ),
        .CO({\dout[15]_INST_0_i_66_n_0 ,\dout[15]_INST_0_i_66_n_1 ,\dout[15]_INST_0_i_66_n_2 ,\dout[15]_INST_0_i_66_n_3 }),
        .CYINIT(\dout[15]_INST_0_i_100_n_0 ),
        .DI(L[11:8]),
        .O({\dout[15]_INST_0_i_66_n_4 ,\dout[15]_INST_0_i_66_n_5 ,\dout[15]_INST_0_i_66_n_6 ,\dout[15]_INST_0_i_66_n_7 }),
        .S({\dout[15]_INST_0_i_101_n_0 ,\dout[15]_INST_0_i_102_n_0 ,\dout[15]_INST_0_i_103_n_0 ,\dout[15]_INST_0_i_104_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_67 
       (.I0(L[15]),
        .I1(\dout[15]_INST_0_i_15_n_0 ),
        .O(\dout[15]_INST_0_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_68 
       (.I0(L[14]),
        .I1(\dout[14]_INST_0_i_9_n_0 ),
        .O(\dout[15]_INST_0_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[15]_INST_0_i_69 
       (.I0(L[13]),
        .I1(\dout[14]_INST_0_i_27_n_0 ),
        .O(\dout[15]_INST_0_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFF8FFFFF8F8)) 
    \dout[15]_INST_0_i_7 
       (.I0(\dout[15]_INST_0_i_16_n_0 ),
        .I1(\dout[15]_INST_0_i_17_n_0 ),
        .I2(\dout[15]_INST_0_i_18_n_0 ),
        .I3(\dout[15]_INST_0_i_19_n_0 ),
        .I4(\dout[15]_INST_0_i_20_n_0 ),
        .I5(\dout[15]_INST_0_i_21_n_4 ),
        .O(\dout[15]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_70 
       (.I0(L[12]),
        .I1(\dout[4]_INST_0_i_13_n_0 ),
        .O(\dout[15]_INST_0_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[15]_INST_0_i_71 
       (.CI(\dout[4]_INST_0_i_44_n_0 ),
        .CO({\dout[15]_INST_0_i_71_n_0 ,\dout[15]_INST_0_i_71_n_1 ,\dout[15]_INST_0_i_71_n_2 ,\dout[15]_INST_0_i_71_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\dout[15]_INST_0_i_71_n_4 ,\dout[15]_INST_0_i_71_n_5 ,\dout[15]_INST_0_i_71_n_6 ,\dout[15]_INST_0_i_71_n_7 }),
        .S({\dout[15]_INST_0_i_61_n_4 ,\dout[15]_INST_0_i_61_n_5 ,\dout[15]_INST_0_i_61_n_6 ,\dout[15]_INST_0_i_61_n_7 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h003F1D1D00000000)) 
    \dout[15]_INST_0_i_76 
       (.I0(data4[7]),
        .I1(eqOp93_in),
        .I2(bw),
        .I3(src__0[7]),
        .I4(\dout[5]_INST_0_i_14_n_0 ),
        .I5(\dout[5]_INST_0_i_15_n_0 ),
        .O(\dout[15]_INST_0_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000477777774777)) 
    \dout[15]_INST_0_i_77 
       (.I0(soc[2]),
        .I1(eqOp93_in),
        .I2(\dout[15]_INST_0_i_109_n_0 ),
        .I3(din[15]),
        .I4(\dout[5]_INST_0_i_14_n_0 ),
        .I5(src__0[15]),
        .O(\dout[15]_INST_0_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \dout[15]_INST_0_i_8 
       (.I0(\dout[15]_INST_0_i_22_n_0 ),
        .I1(\dout[15]_INST_0_i_23_n_0 ),
        .O(\dout[15]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[15]_INST_0_i_81 
       (.I0(L[8]),
        .I1(\dout[9]_INST_0_i_11_n_0 ),
        .O(\dout[15]_INST_0_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[15]_INST_0_i_82 
       (.I0(\rrd[0] [7]),
        .I1(\dout[14]_INST_0_i_25_n_0 ),
        .I2(pc[7]),
        .I3(eqOp93_in),
        .I4(data4[7]),
        .O(\dout[15]_INST_0_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8BBB8888)) 
    \dout[15]_INST_0_i_83 
       (.I0(pc[15]),
        .I1(eqOp93_in),
        .I2(r_a0),
        .I3(bw),
        .I4(din[15]),
        .O(\dout[15]_INST_0_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFE0EFEFEFE0E0E0)) 
    \dout[15]_INST_0_i_84_rewire 
       (.I0(\addr[5]_INST_0_i_6_n_0 ),
        .I1(\rrd[0] [5]),
        .I2(\dout[14]_INST_0_i_25_n_0 ),
        .I3(pc[5]),
        .I4(eqOp93_in),
        .I5(data4[5]),
        .O(\dout[15]_INST_0_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88B8B8B8)) 
    \dout[15]_INST_0_i_85 
       (.I0(pc[13]),
        .I1(eqOp93_in),
        .I2(din[13]),
        .I3(r_a0),
        .I4(bw),
        .O(\dout[15]_INST_0_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88B8B8B8)) 
    \dout[15]_INST_0_i_86 
       (.I0(pc[12]),
        .I1(eqOp93_in),
        .I2(din[12]),
        .I3(r_a0),
        .I4(bw),
        .O(\dout[15]_INST_0_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[15]_INST_0_i_87 
       (.I0(\dout[14]_INST_0_i_9_n_0 ),
        .I1(L[14]),
        .O(\dout[15]_INST_0_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F888FFF88888888)) 
    \dout[15]_INST_0_i_9 
       (.I0(\dout[15]_INST_0_i_24_n_0 ),
        .I1(doc[3]),
        .I2(\dout[15]_INST_0_i_25_n_4 ),
        .I3(bw),
        .I4(\dout[15]_INST_0_i_26_n_4 ),
        .I5(\dout[15]_INST_0_i_20_n_0 ),
        .O(\dout[15]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[15]_INST_0_i_91 
       (.I0(L[8]),
        .I1(sr_reg_n_0_),
        .O(\dout[15]_INST_0_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[15]_INST_0_i_95 
       (.I0(L[8]),
        .I1(\dout[9]_INST_0_i_11_n_0 ),
        .O(\dout[15]_INST_0_i_95_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_96 
       (.I0(L[11]),
        .I1(\dout[11]_INST_0_i_16_n_0 ),
        .O(\dout[15]_INST_0_i_96_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_97 
       (.I0(L[10]),
        .I1(\dout[2]_INST_0_i_12_n_0 ),
        .O(\dout[15]_INST_0_i_97_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_98 
       (.I0(L[9]),
        .I1(\dout[9]_INST_0_i_14_n_0 ),
        .O(\dout[15]_INST_0_i_98_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[15]_INST_0_i_99 
       (.I0(L[8]),
        .I1(\dout[9]_INST_0_i_11_n_0 ),
        .O(\dout[15]_INST_0_i_99_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[1]_INST_0 
       (.I0(pc[1]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[1] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[1]_INST_0_i_1_n_0 ),
        .O(dout[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4447444477777777)) 
    \dout[1]_INST_0_i_10 
       (.I0(\r_code[1]_i_1_n_0 ),
        .I1(eqOp93_in),
        .I2(\dout[13]_INST_0_i_3_n_0 ),
        .I3(rd_INST_0_i_16_n_0),
        .I4(rd_INST_0_i_21_n_0),
        .I5(data4[2]),
        .O(\dout[1]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFDFF)) 
    \dout[1]_INST_0_i_11 
       (.I0(src__0[2]),
        .I1(\dout[13]_INST_0_i_3_n_0 ),
        .I2(rd_INST_0_i_16_n_0),
        .I3(rd_INST_0_i_21_n_0),
        .O(\dout[1]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h22FF000022220202)) 
    \dout[1]_INST_0_i_12 
       (.I0(doc[0]),
        .I1(\dout[15]_INST_0_i_37_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .I3(\dout[2]_INST_0_i_42_n_0 ),
        .I4(\dout[2]_INST_0_i_16_n_0 ),
        .I5(\dout[0]_INST_0_i_10_n_0 ),
        .O(\dout[1]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFEFFFE00)) 
    \dout[1]_INST_0_i_1_rewire_rewire 
       (.I0(\dout[9]_INST_0_i_16_n_0 ),
        .I1(\dout[9]_INST_0_i_8_n_0 ),
        .I2(\dout[9]_INST_0_i_2_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .I4(\dout[1]_INST_0_i_2_n_0 ),
        .O(\dout[1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFEEFE)) 
    \dout[1]_INST_0_i_2 
       (.I0(\dout[1]_INST_0_i_3_n_0 ),
        .I1(\dout[1]_INST_0_i_4_n_0 ),
        .I2(\dout[6]_INST_0_i_5_n_0 ),
        .I3(\dout[1]_INST_0_i_5_n_0 ),
        .I4(\dout[1]_INST_0_i_6_n_0 ),
        .O(\dout[1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \dout[1]_INST_0_i_3 
       (.I0(\dout[15]_INST_0_i_14_n_0 ),
        .I1(\dout[0]_INST_0_i_5_n_0 ),
        .I2(\dout[2]_INST_0_i_6_n_6 ),
        .I3(\dout[4]_INST_0_i_7_n_0 ),
        .I4(\dout[2]_INST_0_i_7_n_6 ),
        .I5(eqOp93_in),
        .O(\dout[1]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \dout[1]_INST_0_i_4 
       (.I0(\dout[1]_INST_0_i_7_n_0 ),
        .I1(\dout[1]_INST_0_i_8_n_0 ),
        .I2(\dout[15]_INST_0_i_23_n_0 ),
        .I3(\dout[1]_INST_0_i_9_n_0 ),
        .I4(\dout[2]_INST_0_i_11_n_6 ),
        .I5(\dout[15]_INST_0_i_19_n_0 ),
        .O(\dout[1]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAA00AAC0FFFFAAC0)) 
    \dout[1]_INST_0_i_5 
       (.I0(\addr[2]_INST_0_i_5_n_0 ),
        .I1(\dout[1]_INST_0_i_10_n_0 ),
        .I2(\dout[1]_INST_0_i_11_n_0 ),
        .I3(\dout[5]_INST_0_i_10_n_0 ),
        .I4(\FSM_sequential_state[1]_i_12_n_0 ),
        .I5(\rrs[0] [2]),
        .O(\dout[1]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h008800A800000020)) 
    \dout[1]_INST_0_i_6 
       (.I0(eqOp135_in),
        .I1(soc[2]),
        .I2(soc[0]),
        .I3(soc[1]),
        .I4(\dout[9]_INST_0_i_14_n_0 ),
        .I5(\dout[0]_INST_0_i_5_n_0 ),
        .O(\dout[1]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF444)) 
    \dout[1]_INST_0_i_7 
       (.I0(\dout[2]_INST_0_i_34_n_0 ),
        .I1(\dout[14]_INST_0_i_10_n_0 ),
        .I2(\dout[2]_INST_0_i_43_n_0 ),
        .I3(\dout[14]_INST_0_i_11_n_0 ),
        .I4(\dout[1]_INST_0_i_12_n_0 ),
        .O(\dout[1]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0069)) 
    \dout[1]_INST_0_i_8 
       (.I0(\dout[4]_INST_0_i_35_n_0 ),
        .I1(\dout[2]_INST_0_i_34_n_0 ),
        .I2(\dout[2]_INST_0_i_44_n_0 ),
        .I3(bw),
        .O(\dout[1]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55404040)) 
    \dout[1]_INST_0_i_9 
       (.I0(bw),
        .I1(\dout[2]_INST_0_i_30_n_6 ),
        .I2(\dout[15]_INST_0_i_20_n_0 ),
        .I3(\dout[2]_INST_0_i_31_n_6 ),
        .I4(\dout[15]_INST_0_i_31_n_0 ),
        .O(\dout[1]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[2]_INST_0 
       (.I0(pc[2]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(p_1_in122_in),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[2]_INST_0_i_1_n_0 ),
        .O(dout[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBBBB8)) 
    \dout[2]_INST_0_i_1 
       (.I0(\dout[10]_INST_0_i_2_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\dout[2]_INST_0_i_2_n_0 ),
        .I3(\dout[2]_INST_0_i_3_n_0 ),
        .I4(\dout[2]_INST_0_i_4_n_0 ),
        .O(\dout[2]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55404040)) 
    \dout[2]_INST_0_i_10 
       (.I0(bw),
        .I1(\dout[2]_INST_0_i_30_n_5 ),
        .I2(\dout[15]_INST_0_i_20_n_0 ),
        .I3(\dout[2]_INST_0_i_31_n_5 ),
        .I4(\dout[15]_INST_0_i_31_n_0 ),
        .O(\dout[2]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[2]_INST_0_i_11 
       (.CI(\<const0>__0__0 ),
        .CO({\dout[2]_INST_0_i_11_n_0 ,\dout[2]_INST_0_i_11_n_1 ,\dout[2]_INST_0_i_11_n_2 ,\dout[2]_INST_0_i_11_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\dout[2]_INST_0_i_14_n_0 ,\dout[2]_INST_0_i_15_n_0 ,\dout[2]_INST_0_i_16_n_0 ,\dout[2]_INST_0_i_17_n_0 }),
        .O({\dout[2]_INST_0_i_11_n_4 ,\dout[2]_INST_0_i_11_n_5 ,\dout[2]_INST_0_i_11_n_6 ,\dout[2]_INST_0_i_11_n_7 }),
        .S({\dout[2]_INST_0_i_32_n_0 ,\dout[2]_INST_0_i_33_n_0 ,\dout[2]_INST_0_i_34_n_0 ,\dout[2]_INST_0_i_35_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \dout[2]_INST_0_i_12 
       (.I0(\dout[2]_INST_0_i_36_n_0 ),
        .I1(\dout[1]_INST_0_i_5_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[2]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000BB0B)) 
    \dout[2]_INST_0_i_13 
       (.I0(\rrs[0] [3]),
        .I1(\FSM_sequential_state[1]_i_12_n_0 ),
        .I2(\dout[5]_INST_0_i_10_n_0 ),
        .I3(\addr[3]_INST_0_i_6_n_0 ),
        .I4(\dout[2]_INST_0_i_37_n_0 ),
        .O(\dout[2]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \dout[2]_INST_0_i_14 
       (.I0(data4[3]),
        .I1(eqOp93_in),
        .I2(pc[3]),
        .I3(\dout[14]_INST_0_i_25_n_0 ),
        .I4(\rrd[0] [3]),
        .I5(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[2]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \dout[2]_INST_0_i_15 
       (.I0(data4[2]),
        .I1(eqOp93_in),
        .I2(pc[2]),
        .I3(\dout[14]_INST_0_i_25_n_0 ),
        .I4(\rrd[0] [2]),
        .I5(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[2]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFD100D1)) 
    \dout[2]_INST_0_i_16 
       (.I0(\dout[2]_INST_0_i_38_n_0 ),
        .I1(eqOp93_in),
        .I2(pc[1]),
        .I3(\dout[14]_INST_0_i_25_n_0 ),
        .I4(\rrd[0] [1]),
        .I5(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[2]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEEEE222)) 
    \dout[2]_INST_0_i_17 
       (.I0(\dout[2]_INST_0_i_40_n_0 ),
        .I1(\dout[14]_INST_0_i_25_n_0 ),
        .I2(\addr[15]_INST_0_i_11_n_0 ),
        .I3(\addr[3]_INST_0_i_50_n_0 ),
        .I4(lbe_INST_0_i_7_n_0),
        .I5(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[2]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAA9A99)) 
    \dout[2]_INST_0_i_18 
       (.I0(\dout[2]_INST_0_i_14_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\rrs[0] [3]),
        .I3(\FSM_sequential_state[1]_i_12_n_0 ),
        .I4(\dout[2]_INST_0_i_41_n_0 ),
        .I5(\dout[2]_INST_0_i_37_n_0 ),
        .O(\dout[2]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \dout[2]_INST_0_i_19 
       (.I0(\dout[2]_INST_0_i_15_n_0 ),
        .I1(\dout[1]_INST_0_i_5_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[2]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \dout[2]_INST_0_i_2 
       (.I0(\dout[15]_INST_0_i_14_n_0 ),
        .I1(\dout[2]_INST_0_i_5_n_0 ),
        .I2(\dout[2]_INST_0_i_6_n_5 ),
        .I3(\dout[4]_INST_0_i_7_n_0 ),
        .I4(\dout[2]_INST_0_i_7_n_5 ),
        .I5(eqOp93_in),
        .O(\dout[2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \dout[2]_INST_0_i_20 
       (.I0(\dout[2]_INST_0_i_16_n_0 ),
        .I1(\dout[0]_INST_0_i_10_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[2]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[2]_INST_0_i_21 
       (.I0(\dout[2]_INST_0_i_17_n_0 ),
        .I1(\dout[2]_INST_0_i_45_n_0 ),
        .O(\dout[2]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h9A)) 
    \dout[2]_INST_0_i_22 
       (.I0(\dout[2]_INST_0_i_14_n_0 ),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[11]_INST_0_i_26_n_0 ),
        .O(\dout[2]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h9A)) 
    \dout[2]_INST_0_i_23 
       (.I0(\dout[2]_INST_0_i_15_n_0 ),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[2]_INST_0_i_5_n_0 ),
        .O(\dout[2]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h9A)) 
    \dout[2]_INST_0_i_24 
       (.I0(\dout[2]_INST_0_i_16_n_0 ),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[0]_INST_0_i_5_n_0 ),
        .O(\dout[2]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hA9)) 
    \dout[2]_INST_0_i_25 
       (.I0(\dout[2]_INST_0_i_17_n_0 ),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[2]_INST_0_i_45_n_0 ),
        .O(\dout[2]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h56)) 
    \dout[2]_INST_0_i_26 
       (.I0(\dout[2]_INST_0_i_15_n_0 ),
        .I1(\dout[1]_INST_0_i_5_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[2]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[2]_INST_0_i_27 
       (.I0(\dout[2]_INST_0_i_15_n_0 ),
        .I1(\dout[1]_INST_0_i_5_n_0 ),
        .O(\dout[2]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h22FF000022220202)) 
    \dout[2]_INST_0_i_28 
       (.I0(doc[0]),
        .I1(\dout[15]_INST_0_i_37_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .I3(\dout[2]_INST_0_i_42_n_0 ),
        .I4(\dout[2]_INST_0_i_15_n_0 ),
        .I5(\dout[1]_INST_0_i_5_n_0 ),
        .O(\dout[2]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h933C93969396C66C)) 
    \dout[2]_INST_0_i_29 
       (.I0(\dout[4]_INST_0_i_35_n_0 ),
        .I1(\dout[2]_INST_0_i_33_n_0 ),
        .I2(\dout[2]_INST_0_i_43_n_0 ),
        .I3(\dout[2]_INST_0_i_44_n_0 ),
        .I4(\dout[0]_INST_0_i_5_n_0 ),
        .I5(\dout[2]_INST_0_i_16_n_0 ),
        .O(\dout[2]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \dout[2]_INST_0_i_3 
       (.I0(\dout[2]_INST_0_i_8_n_0 ),
        .I1(\dout[2]_INST_0_i_9_n_0 ),
        .I2(\dout[15]_INST_0_i_23_n_0 ),
        .I3(\dout[2]_INST_0_i_10_n_0 ),
        .I4(\dout[2]_INST_0_i_11_n_5 ),
        .I5(\dout[15]_INST_0_i_19_n_0 ),
        .O(\dout[2]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[2]_INST_0_i_30 
       (.CI(\<const0>__0__0 ),
        .CO({\dout[2]_INST_0_i_30_n_0 ,\dout[2]_INST_0_i_30_n_1 ,\dout[2]_INST_0_i_30_n_2 ,\dout[2]_INST_0_i_30_n_3 }),
        .CYINIT(\dout[2]_INST_0_i_45_n_0 ),
        .DI({\dout[2]_INST_0_i_14_n_0 ,\dout[2]_INST_0_i_15_n_0 ,\dout[2]_INST_0_i_16_n_0 ,\dout[2]_INST_0_i_17_n_0 }),
        .O({\dout[2]_INST_0_i_30_n_4 ,\dout[2]_INST_0_i_30_n_5 ,\dout[2]_INST_0_i_30_n_6 ,\dout[2]_INST_0_i_30_n_7 }),
        .S({\dout[2]_INST_0_i_46_n_0 ,\dout[2]_INST_0_i_33_n_0 ,\dout[2]_INST_0_i_34_n_0 ,\dout[2]_INST_0_i_49_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[2]_INST_0_i_31 
       (.CI(\<const0>__0__0 ),
        .CO({\dout[2]_INST_0_i_31_n_0 ,\dout[2]_INST_0_i_31_n_1 ,\dout[2]_INST_0_i_31_n_2 ,\dout[2]_INST_0_i_31_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\dout[2]_INST_0_i_6_n_7 }),
        .O({\dout[2]_INST_0_i_31_n_4 ,\dout[2]_INST_0_i_31_n_5 ,\dout[2]_INST_0_i_31_n_6 ,\dout[2]_INST_0_i_31_n_7 }),
        .S({\dout[2]_INST_0_i_6_n_4 ,\dout[2]_INST_0_i_6_n_5 ,\dout[2]_INST_0_i_6_n_6 ,\dout[2]_INST_0_i_53_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[2]_INST_0_i_32 
       (.I0(\dout[11]_INST_0_i_26_n_0 ),
        .I1(\dout[2]_INST_0_i_14_n_0 ),
        .O(\dout[2]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h101050503333FF00)) 
    \dout[2]_INST_0_i_36_rewire 
       (.I0(\addr[10]_INST_0_i_4_n_0 ),
        .I1(\addr[10]_INST_0_i_8_n_0 ),
        .I2(\addr[10]_INST_0_i_1_n_0 ),
        .I3(\dout[2]_INST_0_i_56_n_0 ),
        .I4(\dout[5]_INST_0_i_10_n_0 ),
        .I5(\FSM_sequential_state[1]_i_12_n_0 ),
        .O(\dout[2]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00F3D1D100000000)) 
    \dout[2]_INST_0_i_37 
       (.I0(data4[3]),
        .I1(eqOp93_in),
        .I2(\addr[3]_INST_0_i_9_n_0 ),
        .I3(src__0[3]),
        .I4(\dout[5]_INST_0_i_14_n_0 ),
        .I5(\dout[5]_INST_0_i_15_n_0 ),
        .O(\dout[2]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h15D5)) 
    \dout[2]_INST_0_i_38 
       (.I0(din[1]),
        .I1(bw),
        .I2(r_a0),
        .I3(din[9]),
        .O(\dout[2]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFDDDDDDD0)) 
    \dout[2]_INST_0_i_39 
       (.I0(\addr[1]_INST_0_i_7_n_0 ),
        .I1(\addr[1]_INST_0_i_8_n_0 ),
        .I2(\addr[1]_INST_0_i_9_n_0 ),
        .I3(\addr[1]_INST_0_i_10_n_0 ),
        .I4(\addr[1]_INST_0_i_11_n_0 ),
        .I5(\dout[2]_INST_0_i_57_n_0 ),
        .O(\rrd[0] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF11F111F111F1)) 
    \dout[2]_INST_0_i_4 
       (.I0(\dout[2]_INST_0_i_12_n_0 ),
        .I1(\dout[4]_INST_0_i_14_n_0 ),
        .I2(\dout[2]_INST_0_i_5_n_0 ),
        .I3(\dout[4]_INST_0_i_15_n_0 ),
        .I4(\dout[2]_INST_0_i_13_n_0 ),
        .I5(\dout[6]_INST_0_i_5_n_0 ),
        .O(\dout[2]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFEA2A0000EA2A)) 
    \dout[2]_INST_0_i_40 
       (.I0(din[0]),
        .I1(bw),
        .I2(r_a0),
        .I3(din[8]),
        .I4(eqOp93_in),
        .I5(pc[0]),
        .O(\dout[2]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \dout[2]_INST_0_i_41 
       (.I0(\dout[5]_INST_0_i_10_n_0 ),
        .I1(\addr[3]_INST_0_i_33_n_0 ),
        .I2(\r_code[10]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_34_n_0 ),
        .I4(\r_code[11]_i_1_n_0 ),
        .I5(\addr[3]_INST_0_i_20_n_0 ),
        .O(\dout[2]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF47FF)) 
    \dout[2]_INST_0_i_42 
       (.I0(din[14]),
        .I1(p_2_in88_in),
        .I2(r_code[14]),
        .I3(doc[3]),
        .I4(doc[0]),
        .I5(doc[1]),
        .O(\dout[2]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[2]_INST_0_i_43 
       (.I0(\dout[2]_INST_0_i_16_n_0 ),
        .I1(\dout[0]_INST_0_i_10_n_0 ),
        .O(\dout[2]_INST_0_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hAB22)) 
    \dout[2]_INST_0_i_44 
       (.I0(\dout[2]_INST_0_i_17_n_0 ),
        .I1(\dout[9]_INST_0_i_18_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .I3(sr_reg_n_0_),
        .O(\dout[2]_INST_0_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[2]_INST_0_i_46 
       (.I0(\dout[11]_INST_0_i_26_n_0 ),
        .I1(\dout[2]_INST_0_i_14_n_0 ),
        .O(\dout[2]_INST_0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[2]_INST_0_i_49 
       (.I0(\dout[2]_INST_0_i_17_n_0 ),
        .I1(sr_reg_n_0_),
        .O(\dout[2]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \dout[2]_INST_0_i_5 
       (.I0(\dout[15]_INST_0_i_11_n_0 ),
        .I1(\dout[1]_INST_0_i_5_n_0 ),
        .O(\dout[2]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[2]_INST_0_i_53 
       (.I0(\dout[2]_INST_0_i_6_n_7 ),
        .I1(sr_reg_n_0_),
        .O(\dout[2]_INST_0_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h56)) 
    \dout[2]_INST_0_i_54 
       (.I0(\dout[2]_INST_0_i_16_n_0 ),
        .I1(\dout[0]_INST_0_i_10_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[2]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[2]_INST_0_i_55 
       (.I0(\dout[2]_INST_0_i_17_n_0 ),
        .I1(\dout[2]_INST_0_i_45_n_0 ),
        .O(\dout[2]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000477777774777)) 
    \dout[2]_INST_0_i_56 
       (.I0(soc[2]),
        .I1(eqOp93_in),
        .I2(din[10]),
        .I3(\dout[15]_INST_0_i_109_n_0 ),
        .I4(\dout[5]_INST_0_i_14_n_0 ),
        .I5(src__0[10]),
        .O(\dout[2]_INST_0_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00AA08AA00000800)) 
    \dout[2]_INST_0_i_57 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(\sr_reg_n_0_[1] ),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(soc[0]),
        .I5(\addr[1]_INST_0_i_17_n_0 ),
        .O(\dout[2]_INST_0_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[2]_INST_0_i_6 
       (.CI(\<const0>__0__0 ),
        .CO({\dout[2]_INST_0_i_6_n_0 ,\dout[2]_INST_0_i_6_n_1 ,\dout[2]_INST_0_i_6_n_2 ,\dout[2]_INST_0_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\dout[2]_INST_0_i_14_n_0 ,\dout[2]_INST_0_i_15_n_0 ,\dout[2]_INST_0_i_16_n_0 ,\dout[2]_INST_0_i_17_n_0 }),
        .O({\dout[2]_INST_0_i_6_n_4 ,\dout[2]_INST_0_i_6_n_5 ,\dout[2]_INST_0_i_6_n_6 ,\dout[2]_INST_0_i_6_n_7 }),
        .S({\dout[2]_INST_0_i_18_n_0 ,\dout[2]_INST_0_i_19_n_0 ,\dout[2]_INST_0_i_20_n_0 ,\dout[2]_INST_0_i_21_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[2]_INST_0_i_7 
       (.CI(\<const0>__0__0 ),
        .CO({\dout[2]_INST_0_i_7_n_0 ,\dout[2]_INST_0_i_7_n_1 ,\dout[2]_INST_0_i_7_n_2 ,\dout[2]_INST_0_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\dout[2]_INST_0_i_14_n_0 ,\dout[2]_INST_0_i_15_n_0 ,\dout[2]_INST_0_i_16_n_0 ,\dout[2]_INST_0_i_17_n_0 }),
        .O({\dout[2]_INST_0_i_7_n_4 ,\dout[2]_INST_0_i_7_n_5 ,\dout[2]_INST_0_i_7_n_6 ,\dout[2]_INST_0_i_7_n_7 }),
        .S({\dout[2]_INST_0_i_22_n_0 ,\dout[2]_INST_0_i_23_n_0 ,\dout[2]_INST_0_i_24_n_0 ,\dout[2]_INST_0_i_25_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF222)) 
    \dout[2]_INST_0_i_8 
       (.I0(\dout[14]_INST_0_i_10_n_0 ),
        .I1(\dout[2]_INST_0_i_33_n_0 ),
        .I2(\dout[2]_INST_0_i_27_n_0 ),
        .I3(\dout[14]_INST_0_i_11_n_0 ),
        .I4(\dout[2]_INST_0_i_28_n_0 ),
        .O(\dout[2]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \dout[2]_INST_0_i_9 
       (.I0(bw),
        .I1(\dout[2]_INST_0_i_29_n_0 ),
        .O(\dout[2]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[3]_INST_0 
       (.I0(pc[3]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(p_1_in108_in),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[3]_INST_0_i_1_n_0 ),
        .O(dout[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h003F1D1D00000000)) 
    \dout[3]_INST_0_i_10 
       (.I0(data4[4]),
        .I1(eqOp93_in),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(src__0[4]),
        .I4(\dout[5]_INST_0_i_14_n_0 ),
        .I5(\dout[5]_INST_0_i_15_n_0 ),
        .O(\dout[3]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCEFFFFFFCFFFFFFF)) 
    \dout[3]_INST_0_i_11 
       (.I0(\dout[2]_INST_0_i_13_n_0 ),
        .I1(doc[1]),
        .I2(doc[0]),
        .I3(doc[3]),
        .I4(doc[2]),
        .I5(\dout[2]_INST_0_i_14_n_0 ),
        .O(\dout[3]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9999999999966666)) 
    \dout[3]_INST_0_i_12 
       (.I0(\dout[11]_INST_0_i_26_n_0 ),
        .I1(\dout[2]_INST_0_i_14_n_0 ),
        .I2(\dout[2]_INST_0_i_5_n_0 ),
        .I3(\dout[2]_INST_0_i_15_n_0 ),
        .I4(\dout[4]_INST_0_i_61_n_0 ),
        .I5(\dout[2]_INST_0_i_27_n_0 ),
        .O(\dout[3]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8E71718E718E8E71)) 
    \dout[3]_INST_0_i_13 
       (.I0(\dout[3]_INST_0_i_14_n_0 ),
        .I1(\dout[2]_INST_0_i_43_n_0 ),
        .I2(\dout[2]_INST_0_i_33_n_0 ),
        .I3(\dout[2]_INST_0_i_27_n_0 ),
        .I4(\dout[2]_INST_0_i_14_n_0 ),
        .I5(\dout[11]_INST_0_i_26_n_0 ),
        .O(\dout[3]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hD)) 
    \dout[3]_INST_0_i_14 
       (.I0(\dout[2]_INST_0_i_34_n_0 ),
        .I1(\dout[2]_INST_0_i_44_n_0 ),
        .O(\dout[3]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCFCA)) 
    \dout[3]_INST_0_i_1_rewire 
       (.I0(\dout[3]_INST_0_i_4_n_0 ),
        .I1(\dout[11]_INST_0_i_2_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .I3(\dout[3]_INST_0_i_2_n_0 ),
        .O(\dout[3]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFDCCC)) 
    \dout[3]_INST_0_i_2_rewire_rewire 
       (.I0(\dout[3]_INST_0_i_10_n_0 ),
        .I1(\dout[3]_INST_0_i_3_n_0 ),
        .I2(\dout[3]_INST_0_i_5_n_0 ),
        .I3(\dout[6]_INST_0_i_5_n_0 ),
        .I4(\dout[3]_INST_0_i_6_n_0 ),
        .O(\dout[3]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \dout[3]_INST_0_i_3 
       (.I0(\dout[15]_INST_0_i_14_n_0 ),
        .I1(\dout[11]_INST_0_i_26_n_0 ),
        .I2(\dout[2]_INST_0_i_7_n_4 ),
        .I3(eqOp93_in),
        .I4(\dout[2]_INST_0_i_6_n_4 ),
        .I5(\dout[4]_INST_0_i_7_n_0 ),
        .O(\dout[3]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \dout[3]_INST_0_i_4 
       (.I0(\dout[3]_INST_0_i_7_n_0 ),
        .I1(\dout[3]_INST_0_i_8_n_0 ),
        .I2(\dout[15]_INST_0_i_23_n_0 ),
        .I3(\dout[3]_INST_0_i_9_n_0 ),
        .I4(\dout[2]_INST_0_i_11_n_4 ),
        .I5(\dout[15]_INST_0_i_19_n_0 ),
        .O(\dout[3]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3F3F2A3F)) 
    \dout[3]_INST_0_i_5_rewire_rewire 
       (.I0(\addr[4]_INST_0_i_7_n_0 ),
        .I1(\dout[5]_INST_0_i_10_n_0 ),
        .I2(\addr[4]_INST_0_i_5_n_0 ),
        .I3(\FSM_sequential_state[1]_i_12_n_0 ),
        .I4(\rrs[0] [4]),
        .O(\dout[3]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "dout[3]_INST_0_i_5_rewire_rewire" *) 
  LUT5 #(
    .INIT(32'h3F3F2A3F)) 
    \dout[3]_INST_0_i_5_rewire_rewire_replica 
       (.I0(\addr[4]_INST_0_i_7_n_0_repN ),
        .I1(\dout[5]_INST_0_i_10_n_0 ),
        .I2(\addr[4]_INST_0_i_5_n_0 ),
        .I3(\FSM_sequential_state[1]_i_12_n_0 ),
        .I4(\rrs[0] [4]),
        .O(\dout[3]_INST_0_i_5_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h008800A800000020)) 
    \dout[3]_INST_0_i_6 
       (.I0(eqOp135_in),
        .I1(soc[2]),
        .I2(soc[0]),
        .I3(soc[1]),
        .I4(\dout[11]_INST_0_i_16_n_0 ),
        .I5(\dout[11]_INST_0_i_26_n_0 ),
        .O(\dout[3]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFDFD00D0DD5D00D0)) 
    \dout[3]_INST_0_i_7 
       (.I0(\dout[3]_INST_0_i_11_n_0 ),
        .I1(\dout[14]_INST_0_i_10_n_0 ),
        .I2(\dout[2]_INST_0_i_13_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .I4(\dout[2]_INST_0_i_14_n_0 ),
        .I5(\dout[14]_INST_0_i_11_n_0 ),
        .O(\dout[3]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \dout[3]_INST_0_i_8 
       (.I0(\dout[3]_INST_0_i_12_n_0 ),
        .I1(\dout[4]_INST_0_i_35_n_0 ),
        .I2(\dout[3]_INST_0_i_13_n_0 ),
        .I3(bw),
        .O(\dout[3]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55404040)) 
    \dout[3]_INST_0_i_9 
       (.I0(bw),
        .I1(\dout[2]_INST_0_i_30_n_4 ),
        .I2(\dout[15]_INST_0_i_20_n_0 ),
        .I3(\dout[2]_INST_0_i_31_n_4 ),
        .I4(\dout[15]_INST_0_i_31_n_0 ),
        .O(\dout[3]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[4]_INST_0 
       (.I0(pc[4]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[4] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[4]_INST_0_i_1_n_0 ),
        .O(dout[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBBBB8)) 
    \dout[4]_INST_0_i_1 
       (.I0(\dout[12]_INST_0_i_2_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\dout[4]_INST_0_i_2_n_0 ),
        .I3(\dout[4]_INST_0_i_3_n_0 ),
        .I4(\dout[4]_INST_0_i_4_n_0 ),
        .O(\dout[4]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4114)) 
    \dout[4]_INST_0_i_10 
       (.I0(bw),
        .I1(\dout[4]_INST_0_i_34_n_0 ),
        .I2(\dout[4]_INST_0_i_5_n_0 ),
        .I3(\dout[4]_INST_0_i_35_n_0 ),
        .O(\dout[4]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[4]_INST_0_i_11 
       (.CI(\dout[2]_INST_0_i_11_n_0 ),
        .CO({\dout[4]_INST_0_i_11_n_0 ,\dout[4]_INST_0_i_11_n_1 ,\dout[4]_INST_0_i_11_n_2 ,\dout[4]_INST_0_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\dout[4]_INST_0_i_36_n_0 ,\dout[4]_INST_0_i_37_n_0 ,\dout[4]_INST_0_i_38_n_0 ,\dout[4]_INST_0_i_20_n_0 }),
        .O({\dout[4]_INST_0_i_11_n_4 ,\dout[4]_INST_0_i_11_n_5 ,\dout[4]_INST_0_i_11_n_6 ,\dout[4]_INST_0_i_11_n_7 }),
        .S({\dout[4]_INST_0_i_39_n_0 ,\dout[4]_INST_0_i_40_n_0 ,\dout[4]_INST_0_i_41_n_0 ,\dout[4]_INST_0_i_42_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55404040)) 
    \dout[4]_INST_0_i_12 
       (.I0(bw),
        .I1(\dout[4]_INST_0_i_43_n_7 ),
        .I2(\dout[15]_INST_0_i_20_n_0 ),
        .I3(\dout[4]_INST_0_i_44_n_7 ),
        .I4(\dout[15]_INST_0_i_31_n_0 ),
        .O(\dout[4]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBFB0)) 
    \dout[4]_INST_0_i_13_rewire 
       (.I0(\dout[3]_INST_0_i_10_n_0 ),
        .I1(\dout[3]_INST_0_i_5_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .I3(\dout[4]_INST_0_i_45_n_0 ),
        .O(\dout[4]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBFBFBFFFFFFFBFF)) 
    \dout[4]_INST_0_i_14 
       (.I0(soc[1]),
        .I1(eqOp135_in),
        .I2(soc[2]),
        .I3(r_code[7]),
        .I4(p_2_in88_in),
        .I5(din[7]),
        .O(\dout[4]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \dout[4]_INST_0_i_15 
       (.I0(soc[1]),
        .I1(soc[2]),
        .I2(eqOp135_in),
        .O(\dout[4]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000045CF45CF45CF)) 
    \dout[4]_INST_0_i_16_replica_rewire 
       (.I0(\dout[5]_INST_0_i_15_n_0 ),
        .I1(\rrs[0] [5]),
        .I2(\FSM_sequential_state[1]_i_12_n_0 ),
        .I3(\dout[4]_INST_0_i_46_n_0 ),
        .I4(\addr[5]_INST_0_i_8_n_0 ),
        .I5(\dout[5]_INST_0_i_10_n_0 ),
        .O(\dout[4]_INST_0_i_16_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0BBB)) 
    \dout[4]_INST_0_i_16_rewire 
       (.I0(\rrs[0] [5]),
        .I1(\FSM_sequential_state[1]_i_12_n_0 ),
        .I2(\addr[5]_INST_0_i_8_n_0 ),
        .I3(\dout[5]_INST_0_i_10_n_0 ),
        .O(\dout[4]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[4]_INST_0_i_17 
       (.I0(\dout[15]_INST_0_i_82_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[4]_INST_0_i_18 
       (.I0(\dout[14]_INST_0_i_23_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[4]_INST_0_i_19 
       (.I0(\dout[15]_INST_0_i_84_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \dout[4]_INST_0_i_2 
       (.I0(\dout[15]_INST_0_i_14_n_0 ),
        .I1(\dout[4]_INST_0_i_5_n_0 ),
        .I2(\dout[4]_INST_0_i_6_n_7 ),
        .I3(\dout[4]_INST_0_i_7_n_0 ),
        .I4(\dout[4]_INST_0_i_8_n_7 ),
        .I5(eqOp93_in),
        .O(\dout[4]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \dout[4]_INST_0_i_20 
       (.I0(data4[4]),
        .I1(eqOp93_in),
        .I2(pc[4]),
        .I3(\dout[14]_INST_0_i_25_n_0 ),
        .I4(\rrd[0] [4]),
        .I5(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6AC0)) 
    \dout[4]_INST_0_i_21_rewire_rewire 
       (.I0(\dout[15]_INST_0_i_33_n_0 ),
        .I1(\dout[15]_INST_0_i_82_n_0 ),
        .I2(\dout[9]_INST_0_i_22_n_0 ),
        .I3(\dout[7]_INST_0_i_7_n_0 ),
        .O(\dout[4]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44B400F0)) 
    \dout[4]_INST_0_i_22_rewire_rewire 
       (.I0(\dout[5]_INST_0_i_11_n_0 ),
        .I1(\dout[5]_INST_0_i_5_n_0 ),
        .I2(\dout[14]_INST_0_i_23_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .I4(\dout[6]_INST_0_i_7_n_0 ),
        .O(\dout[4]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6AC0)) 
    \dout[4]_INST_0_i_23_rewire_rewire 
       (.I0(\dout[4]_INST_0_i_16_n_0 ),
        .I1(\dout[15]_INST_0_i_84_n_0 ),
        .I2(\dout[5]_INST_0_i_12_n_0 ),
        .I3(\dout[13]_INST_0_i_20_n_0 ),
        .O(\dout[4]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \dout[4]_INST_0_i_24 
       (.I0(\dout[4]_INST_0_i_20_n_0 ),
        .I1(\dout[4]_INST_0_i_5_n_0 ),
        .O(\dout[4]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[4]_INST_0_i_25 
       (.I0(\dout[15]_INST_0_i_82_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[4]_INST_0_i_26 
       (.I0(\dout[14]_INST_0_i_23_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[4]_INST_0_i_27 
       (.I0(\dout[15]_INST_0_i_84_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC06AC0C0)) 
    \dout[4]_INST_0_i_28_rewire_rewire 
       (.I0(\dout[15]_INST_0_i_33_n_0 ),
        .I1(\dout[15]_INST_0_i_82_n_0 ),
        .I2(\dout[9]_INST_0_i_22_n_0 ),
        .I3(\dout[13]_INST_0_i_22_n_0 ),
        .I4(\dout[7]_INST_0_i_7_n_0 ),
        .O(\dout[4]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00F044B400F000F0)) 
    \dout[4]_INST_0_i_29_rewire_rewire 
       (.I0(\dout[5]_INST_0_i_11_n_0 ),
        .I1(\dout[5]_INST_0_i_5_n_0 ),
        .I2(\dout[14]_INST_0_i_23_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .I4(\dout[13]_INST_0_i_22_n_0 ),
        .I5(\dout[6]_INST_0_i_7_n_0 ),
        .O(\dout[4]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \dout[4]_INST_0_i_3 
       (.I0(\dout[4]_INST_0_i_9_n_0 ),
        .I1(\dout[4]_INST_0_i_10_n_0 ),
        .I2(\dout[15]_INST_0_i_23_n_0 ),
        .I3(\dout[4]_INST_0_i_11_n_7 ),
        .I4(\dout[15]_INST_0_i_19_n_0 ),
        .I5(\dout[4]_INST_0_i_12_n_0 ),
        .O(\dout[4]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC06AC0C0)) 
    \dout[4]_INST_0_i_30_rewire_rewire 
       (.I0(\dout[4]_INST_0_i_16_n_0 ),
        .I1(\dout[15]_INST_0_i_84_n_0 ),
        .I2(\dout[5]_INST_0_i_12_n_0 ),
        .I3(\dout[13]_INST_0_i_22_n_0 ),
        .I4(\dout[13]_INST_0_i_20_n_0 ),
        .O(\dout[4]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h9A)) 
    \dout[4]_INST_0_i_31 
       (.I0(\dout[4]_INST_0_i_20_n_0 ),
        .I1(\dout[13]_INST_0_i_22_n_0 ),
        .I2(\dout[4]_INST_0_i_5_n_0 ),
        .O(\dout[4]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \dout[4]_INST_0_i_32_rewire 
       (.I0(\dout[3]_INST_0_i_10_n_0 ),
        .I1(\dout[4]_INST_0_i_20_n_0 ),
        .I2(\dout[3]_INST_0_i_5_n_0 ),
        .O(\dout[4]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FA00FF00100000)) 
    \dout[4]_INST_0_i_33_rewire 
       (.I0(\dout[3]_INST_0_i_10_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(doc[0]),
        .I3(\dout[15]_INST_0_i_37_n_0 ),
        .I4(\dout[3]_INST_0_i_5_n_0 ),
        .I5(\dout[4]_INST_0_i_20_n_0 ),
        .O(\dout[4]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[4]_INST_0_i_34 
       (.I0(\rrd[0] [4]),
        .I1(\dout[14]_INST_0_i_25_n_0 ),
        .I2(pc[4]),
        .I3(eqOp93_in),
        .I4(data4[4]),
        .O(\dout[4]_INST_0_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hDD04FF5D)) 
    \dout[4]_INST_0_i_35 
       (.I0(\dout[4]_INST_0_i_47_n_0 ),
        .I1(\dout[2]_INST_0_i_13_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .I3(\dout[2]_INST_0_i_14_n_0 ),
        .I4(\dout[4]_INST_0_i_48_n_0 ),
        .O(\dout[4]_INST_0_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[4]_INST_0_i_36 
       (.I0(\dout[15]_INST_0_i_82_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[4]_INST_0_i_37 
       (.I0(\dout[14]_INST_0_i_23_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[4]_INST_0_i_38 
       (.I0(\dout[15]_INST_0_i_84_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF11F111F111F1)) 
    \dout[4]_INST_0_i_4 
       (.I0(\dout[4]_INST_0_i_13_n_0 ),
        .I1(\dout[4]_INST_0_i_14_n_0 ),
        .I2(\dout[4]_INST_0_i_5_n_0 ),
        .I3(\dout[4]_INST_0_i_15_n_0 ),
        .I4(\dout[4]_INST_0_i_16_n_0_repN ),
        .I5(\dout[6]_INST_0_i_5_n_0 ),
        .O(\dout[4]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h953F)) 
    \dout[4]_INST_0_i_41_rewire_rewire 
       (.I0(\dout[4]_INST_0_i_16_n_0 ),
        .I1(\dout[15]_INST_0_i_84_n_0 ),
        .I2(\dout[5]_INST_0_i_12_n_0 ),
        .I3(\dout[13]_INST_0_i_20_n_0 ),
        .O(\dout[4]_INST_0_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[4]_INST_0_i_42 
       (.I0(\dout[4]_INST_0_i_20_n_0 ),
        .I1(\dout[4]_INST_0_i_5_n_0 ),
        .O(\dout[4]_INST_0_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[4]_INST_0_i_43 
       (.CI(\dout[2]_INST_0_i_30_n_0 ),
        .CO({\dout[4]_INST_0_i_43_n_0 ,\dout[4]_INST_0_i_43_n_1 ,\dout[4]_INST_0_i_43_n_2 ,\dout[4]_INST_0_i_43_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\dout[4]_INST_0_i_49_n_0 ,\dout[4]_INST_0_i_50_n_0 ,\dout[4]_INST_0_i_51_n_0 ,\dout[4]_INST_0_i_20_n_0 }),
        .O({\dout[4]_INST_0_i_43_n_4 ,\dout[4]_INST_0_i_43_n_5 ,\dout[4]_INST_0_i_43_n_6 ,\dout[4]_INST_0_i_43_n_7 }),
        .S({\dout[4]_INST_0_i_39_n_0 ,\dout[4]_INST_0_i_40_n_0 ,\dout[4]_INST_0_i_54_n_0 ,\dout[4]_INST_0_i_55_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[4]_INST_0_i_44 
       (.CI(\dout[2]_INST_0_i_31_n_0 ),
        .CO({\dout[4]_INST_0_i_44_n_0 ,\dout[4]_INST_0_i_44_n_1 ,\dout[4]_INST_0_i_44_n_2 ,\dout[4]_INST_0_i_44_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\dout[4]_INST_0_i_44_n_4 ,\dout[4]_INST_0_i_44_n_5 ,\dout[4]_INST_0_i_44_n_6 ,\dout[4]_INST_0_i_44_n_7 }),
        .S({\dout[4]_INST_0_i_6_n_4 ,\dout[4]_INST_0_i_6_n_5 ,\dout[4]_INST_0_i_6_n_6 ,\dout[4]_INST_0_i_6_n_7 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h05FF05CC000005CC)) 
    \dout[4]_INST_0_i_45_rewire 
       (.I0(\addr[12]_INST_0_i_4_n_0 ),
        .I1(\dout[4]_INST_0_i_60_n_0 ),
        .I2(\rrs[0] [12]),
        .I3(\FSM_sequential_state[1]_i_12_n_0 ),
        .I4(\dout[5]_INST_0_i_10_n_0 ),
        .I5(\addr[12]_INST_0_i_8_n_0 ),
        .O(\dout[4]_INST_0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h003F1D1D)) 
    \dout[4]_INST_0_i_46_rewire 
       (.I0(data4[5]),
        .I1(eqOp93_in),
        .I2(as[0]),
        .I3(src__0[5]),
        .I4(\dout[5]_INST_0_i_14_n_0 ),
        .O(\dout[4]_INST_0_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0630300C)) 
    \dout[4]_INST_0_i_47 
       (.I0(\dout[2]_INST_0_i_43_n_0 ),
        .I1(\dout[2]_INST_0_i_33_n_0 ),
        .I2(\dout[2]_INST_0_i_44_n_0 ),
        .I3(\dout[2]_INST_0_i_16_n_0 ),
        .I4(\dout[0]_INST_0_i_5_n_0 ),
        .O(\dout[4]_INST_0_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1115)) 
    \dout[4]_INST_0_i_48 
       (.I0(\dout[2]_INST_0_i_27_n_0 ),
        .I1(\dout[4]_INST_0_i_61_n_0 ),
        .I2(\dout[2]_INST_0_i_15_n_0 ),
        .I3(\dout[2]_INST_0_i_5_n_0 ),
        .O(\dout[4]_INST_0_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[4]_INST_0_i_49 
       (.I0(\dout[15]_INST_0_i_82_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[4]_INST_0_i_50 
       (.I0(\dout[14]_INST_0_i_23_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[4]_INST_0_i_51 
       (.I0(\dout[15]_INST_0_i_84_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h953F)) 
    \dout[4]_INST_0_i_54_rewire_rewire 
       (.I0(\dout[4]_INST_0_i_16_n_0 ),
        .I1(\dout[15]_INST_0_i_84_n_0 ),
        .I2(\dout[5]_INST_0_i_12_n_0 ),
        .I3(\dout[13]_INST_0_i_20_n_0 ),
        .O(\dout[4]_INST_0_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \dout[4]_INST_0_i_55 
       (.I0(\dout[4]_INST_0_i_20_n_0 ),
        .I1(\dout[4]_INST_0_i_5_n_0 ),
        .O(\dout[4]_INST_0_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \dout[4]_INST_0_i_5_rewire 
       (.I0(\dout[3]_INST_0_i_10_n_0 ),
        .I1(\dout[3]_INST_0_i_5_n_0_repN ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[4]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[4]_INST_0_i_6 
       (.CI(\dout[2]_INST_0_i_6_n_0 ),
        .CO({\dout[4]_INST_0_i_6_n_0 ,\dout[4]_INST_0_i_6_n_1 ,\dout[4]_INST_0_i_6_n_2 ,\dout[4]_INST_0_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\dout[4]_INST_0_i_17_n_0 ,\dout[4]_INST_0_i_18_n_0 ,\dout[4]_INST_0_i_19_n_0 ,\dout[4]_INST_0_i_20_n_0 }),
        .O({\dout[4]_INST_0_i_6_n_4 ,\dout[4]_INST_0_i_6_n_5 ,\dout[4]_INST_0_i_6_n_6 ,\dout[4]_INST_0_i_6_n_7 }),
        .S({\dout[4]_INST_0_i_21_n_0 ,\dout[4]_INST_0_i_22_n_0 ,\dout[4]_INST_0_i_23_n_0 ,\dout[4]_INST_0_i_24_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000477777774777)) 
    \dout[4]_INST_0_i_60 
       (.I0(soc[2]),
        .I1(eqOp93_in),
        .I2(din[12]),
        .I3(\dout[15]_INST_0_i_109_n_0 ),
        .I4(\dout[5]_INST_0_i_14_n_0 ),
        .I5(src__0[12]),
        .O(\dout[4]_INST_0_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAB220000FFFF0B02)) 
    \dout[4]_INST_0_i_61 
       (.I0(\dout[2]_INST_0_i_17_n_0 ),
        .I1(\dout[9]_INST_0_i_18_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .I3(sr_reg_n_0_),
        .I4(\dout[2]_INST_0_i_16_n_0 ),
        .I5(\dout[0]_INST_0_i_10_n_0 ),
        .O(\dout[4]_INST_0_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000080800A008A80)) 
    \dout[4]_INST_0_i_7 
       (.I0(\dout[15]_INST_0_i_32_n_0 ),
        .I1(din[12]),
        .I2(p_2_in88_in),
        .I3(r_code[12]),
        .I4(din[13]),
        .I5(r_code[13]),
        .O(\dout[4]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \dout[4]_INST_0_i_8 
       (.CI(\dout[2]_INST_0_i_7_n_0 ),
        .CO({\dout[4]_INST_0_i_8_n_0 ,\dout[4]_INST_0_i_8_n_1 ,\dout[4]_INST_0_i_8_n_2 ,\dout[4]_INST_0_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\dout[4]_INST_0_i_25_n_0 ,\dout[4]_INST_0_i_26_n_0 ,\dout[4]_INST_0_i_27_n_0 ,\dout[4]_INST_0_i_20_n_0 }),
        .O({\dout[4]_INST_0_i_8_n_4 ,\dout[4]_INST_0_i_8_n_5 ,\dout[4]_INST_0_i_8_n_6 ,\dout[4]_INST_0_i_8_n_7 }),
        .S({\dout[4]_INST_0_i_28_n_0 ,\dout[4]_INST_0_i_29_n_0 ,\dout[4]_INST_0_i_30_n_0 ,\dout[4]_INST_0_i_31_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFF606060)) 
    \dout[4]_INST_0_i_9 
       (.I0(\dout[4]_INST_0_i_20_n_0 ),
        .I1(\dout[4]_INST_0_i_5_n_0 ),
        .I2(\dout[14]_INST_0_i_10_n_0 ),
        .I3(\dout[14]_INST_0_i_11_n_0 ),
        .I4(\dout[4]_INST_0_i_32_n_0 ),
        .I5(\dout[4]_INST_0_i_33_n_0 ),
        .O(\dout[4]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[5]_INST_0 
       (.I0(pc[5]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[5] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[5]_INST_0_i_1_n_0 ),
        .O(dout[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dout[5]_INST_0_i_1 
       (.I0(\dout[13]_INST_0_i_2_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\dout[5]_INST_0_i_2_n_0 ),
        .O(\dout[5]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0101010055555555)) 
    \dout[5]_INST_0_i_10 
       (.I0(\dout[13]_INST_0_i_3_n_0 ),
        .I1(\r[10][0]_i_5_n_0 ),
        .I2(\r_code[11]_i_1_n_0 ),
        .I3(soc[1]),
        .I4(as[1]),
        .I5(lbe_INST_0_i_8_n_0),
        .O(\dout[5]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h003F1D1D00000000)) 
    \dout[5]_INST_0_i_11 
       (.I0(data4[6]),
        .I1(eqOp93_in),
        .I2(as[1]),
        .I3(src__0[6]),
        .I4(\dout[5]_INST_0_i_14_n_0 ),
        .I5(\dout[5]_INST_0_i_15_n_0 ),
        .O(\dout[5]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "dout[5]_INST_0_i_12" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[5]_INST_0_i_12_replica 
       (.I0(\dout[15]_INST_0_i_84_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[5]_INST_0_i_12_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \dout[5]_INST_0_i_12_rewire 
       (.I0(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[5]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000B0AA3000)) 
    \dout[5]_INST_0_i_13_rewire 
       (.I0(\dout[15]_INST_0_i_84_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(doc[0]),
        .I3(\dout[4]_INST_0_i_16_n_0_repN ),
        .I4(\dout[5]_INST_0_i_12_n_0 ),
        .I5(\dout[15]_INST_0_i_37_n_0 ),
        .O(\dout[5]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \dout[5]_INST_0_i_14 
       (.I0(rd_INST_0_i_21_n_0),
        .I1(rd_INST_0_i_16_n_0),
        .I2(\dout[13]_INST_0_i_3_n_0 ),
        .O(\dout[5]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h45)) 
    \dout[5]_INST_0_i_15 
       (.I0(\dout[5]_INST_0_i_10_n_0 ),
        .I1(rd_INST_0_i_19_n_0),
        .I2(eqOp135_in),
        .O(\dout[5]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFDFCFCFC)) 
    \dout[5]_INST_0_i_2_rewire 
       (.I0(\dout[5]_INST_0_i_11_n_0 ),
        .I1(\dout[5]_INST_0_i_3_n_0 ),
        .I2(\dout[5]_INST_0_i_4_n_0 ),
        .I3(\dout[5]_INST_0_i_5_n_0 ),
        .I4(\dout[6]_INST_0_i_5_n_0 ),
        .I5(\dout[5]_INST_0_i_6_n_0 ),
        .O(\dout[5]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \dout[5]_INST_0_i_3 
       (.I0(\dout[15]_INST_0_i_14_n_0 ),
        .I1(\dout[13]_INST_0_i_20_n_0_repN ),
        .I2(\dout[4]_INST_0_i_6_n_6 ),
        .I3(\dout[4]_INST_0_i_7_n_0 ),
        .I4(\dout[4]_INST_0_i_8_n_6 ),
        .I5(eqOp93_in),
        .O(\dout[5]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \dout[5]_INST_0_i_4 
       (.I0(\dout[5]_INST_0_i_7_n_0 ),
        .I1(\dout[5]_INST_0_i_8_n_0 ),
        .I2(\dout[15]_INST_0_i_23_n_0 ),
        .I3(\dout[5]_INST_0_i_9_n_0 ),
        .I4(\dout[4]_INST_0_i_11_n_6 ),
        .I5(\dout[15]_INST_0_i_19_n_0 ),
        .O(\dout[5]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7707)) 
    \dout[5]_INST_0_i_5_rewire 
       (.I0(\dout[5]_INST_0_i_10_n_0 ),
        .I1(\addr[6]_INST_0_i_8_n_0 ),
        .I2(\FSM_sequential_state[1]_i_12_n_0 ),
        .I3(\rrs[0] [6]),
        .O(\dout[5]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00A8008800200000)) 
    \dout[5]_INST_0_i_6 
       (.I0(eqOp135_in),
        .I1(soc[2]),
        .I2(soc[0]),
        .I3(soc[1]),
        .I4(\dout[14]_INST_0_i_27_n_0 ),
        .I5(\dout[13]_INST_0_i_20_n_0_repN ),
        .O(\dout[5]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFF606060)) 
    \dout[5]_INST_0_i_7 
       (.I0(\dout[5]_INST_0_i_12_n_0_repN ),
        .I1(\dout[13]_INST_0_i_20_n_0_repN ),
        .I2(\dout[14]_INST_0_i_10_n_0 ),
        .I3(\dout[14]_INST_0_i_11_n_0 ),
        .I4(\dout[6]_INST_0_i_13_n_0 ),
        .I5(\dout[5]_INST_0_i_13_n_0 ),
        .O(\dout[5]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h41)) 
    \dout[5]_INST_0_i_8 
       (.I0(bw),
        .I1(\dout[9]_INST_0_i_12_n_0 ),
        .I2(\dout[9]_INST_0_i_21_n_0 ),
        .O(\dout[5]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55404040)) 
    \dout[5]_INST_0_i_9 
       (.I0(bw),
        .I1(\dout[4]_INST_0_i_43_n_6 ),
        .I2(\dout[15]_INST_0_i_20_n_0 ),
        .I3(\dout[4]_INST_0_i_44_n_6 ),
        .I4(\dout[15]_INST_0_i_31_n_0 ),
        .O(\dout[5]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[6]_INST_0 
       (.I0(pc[6]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[6] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[6]_INST_0_i_1_n_0 ),
        .O(dout[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF54FFFFFF540000)) 
    \dout[6]_INST_0_i_1 
       (.I0(\dout[14]_INST_0_i_5_n_0 ),
        .I1(\dout[14]_INST_0_i_4_n_0 ),
        .I2(\dout[14]_INST_0_i_3_n_0 ),
        .I3(\dout[14]_INST_0_i_2_n_0 ),
        .I4(\dout[15]_INST_0_i_11_n_0 ),
        .I5(\dout[6]_INST_0_i_2_n_0 ),
        .O(\dout[6]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55404040)) 
    \dout[6]_INST_0_i_10 
       (.I0(bw),
        .I1(\dout[4]_INST_0_i_43_n_5 ),
        .I2(\dout[15]_INST_0_i_20_n_0 ),
        .I3(\dout[4]_INST_0_i_44_n_5 ),
        .I4(\dout[15]_INST_0_i_31_n_0 ),
        .O(\dout[6]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBB4BFF0F)) 
    \dout[6]_INST_0_i_11_rewire_rewire 
       (.I0(\dout[5]_INST_0_i_11_n_0 ),
        .I1(\dout[5]_INST_0_i_5_n_0 ),
        .I2(\dout[14]_INST_0_i_23_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .I4(\dout[6]_INST_0_i_7_n_0 ),
        .O(\dout[4]_INST_0_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000D0C0000080C)) 
    \dout[6]_INST_0_i_12_rewire 
       (.I0(\dout[5]_INST_0_i_11_n_0 ),
        .I1(\dout[14]_INST_0_i_23_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .I3(\dout[5]_INST_0_i_5_n_0 ),
        .I4(\dout[15]_INST_0_i_37_n_0 ),
        .I5(doc[0]),
        .O(\dout[6]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h07000000)) 
    \dout[6]_INST_0_i_13_rewire_rewire 
       (.I0(\dout[5]_INST_0_i_15_n_0 ),
        .I1(\dout[4]_INST_0_i_46_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .I3(\dout[15]_INST_0_i_84_n_0 ),
        .I4(\dout[4]_INST_0_i_16_n_0 ),
        .O(\dout[6]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000009090999)) 
    \dout[6]_INST_0_i_14 
       (.I0(\dout[5]_INST_0_i_12_n_0_repN ),
        .I1(\dout[13]_INST_0_i_20_n_0_repN ),
        .I2(\dout[4]_INST_0_i_35_n_0 ),
        .I3(\dout[4]_INST_0_i_5_n_0 ),
        .I4(\dout[4]_INST_0_i_20_n_0 ),
        .I5(\dout[4]_INST_0_i_32_n_0 ),
        .O(\dout[6]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "dout[6]_INST_0_i_1" *) 
  LUT6 #(
    .INIT(64'hFF54FFFFFF540000)) 
    \dout[6]_INST_0_i_1_replica 
       (.I0(\dout[14]_INST_0_i_5_n_0 ),
        .I1(\dout[14]_INST_0_i_4_n_0 ),
        .I2(\dout[14]_INST_0_i_3_n_0 ),
        .I3(\dout[14]_INST_0_i_2_n_0 ),
        .I4(\dout[15]_INST_0_i_11_n_0 ),
        .I5(\dout[6]_INST_0_i_2_n_0 ),
        .O(\dout[6]_INST_0_i_1_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFCFCFC)) 
    \dout[6]_INST_0_i_2_rewire 
       (.I0(\dout[15]_INST_0_i_33_n_0 ),
        .I1(\dout[6]_INST_0_i_3_n_0 ),
        .I2(\dout[6]_INST_0_i_4_n_0 ),
        .I3(\dout[7]_INST_0_i_7_n_0 ),
        .I4(\dout[6]_INST_0_i_5_n_0 ),
        .I5(\dout[6]_INST_0_i_6_n_0 ),
        .O(\dout[6]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \dout[6]_INST_0_i_3 
       (.I0(\dout[15]_INST_0_i_14_n_0 ),
        .I1(\dout[6]_INST_0_i_7_n_0_repN ),
        .I2(\dout[4]_INST_0_i_6_n_5 ),
        .I3(\dout[4]_INST_0_i_7_n_0 ),
        .I4(\dout[4]_INST_0_i_8_n_5 ),
        .I5(eqOp93_in),
        .O(\dout[6]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \dout[6]_INST_0_i_4 
       (.I0(\dout[6]_INST_0_i_8_n_0 ),
        .I1(\dout[6]_INST_0_i_9_n_0 ),
        .I2(\dout[15]_INST_0_i_23_n_0 ),
        .I3(\dout[6]_INST_0_i_10_n_0 ),
        .I4(\dout[4]_INST_0_i_11_n_5 ),
        .I5(\dout[15]_INST_0_i_19_n_0 ),
        .O(\dout[6]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00002020000A202A)) 
    \dout[6]_INST_0_i_5 
       (.I0(eqOp135_in),
        .I1(din[9]),
        .I2(p_2_in88_in),
        .I3(r_code[9]),
        .I4(din[7]),
        .I5(r_code[7]),
        .O(\dout[6]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h008800A800000020)) 
    \dout[6]_INST_0_i_6 
       (.I0(eqOp135_in),
        .I1(soc[2]),
        .I2(soc[0]),
        .I3(soc[1]),
        .I4(\dout[14]_INST_0_i_9_n_0 ),
        .I5(\dout[6]_INST_0_i_7_n_0_repN ),
        .O(\dout[6]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "dout[6]_INST_0_i_7_rewire" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \dout[6]_INST_0_i_7_rewire_replica 
       (.I0(\dout[5]_INST_0_i_11_n_0 ),
        .I1(\dout[5]_INST_0_i_5_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[6]_INST_0_i_7_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \dout[6]_INST_0_i_7_rewire_rewire_rewire 
       (.I0(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[6]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF444)) 
    \dout[6]_INST_0_i_8 
       (.I0(\dout[4]_INST_0_i_40_n_0 ),
        .I1(\dout[14]_INST_0_i_10_n_0 ),
        .I2(\dout[14]_INST_0_i_11_n_0 ),
        .I3(\dout[7]_INST_0_i_13_n_0 ),
        .I4(\dout[6]_INST_0_i_12_n_0 ),
        .O(\dout[6]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000411455554114)) 
    \dout[6]_INST_0_i_9 
       (.I0(bw),
        .I1(\dout[4]_INST_0_i_40_n_0 ),
        .I2(\dout[6]_INST_0_i_13_n_0 ),
        .I3(\dout[6]_INST_0_i_14_n_0 ),
        .I4(\dout[9]_INST_0_i_12_n_0 ),
        .I5(\dout[9]_INST_0_i_20_n_0 ),
        .O(\dout[6]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[7]_INST_0 
       (.I0(pc[7]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[7] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[7]_INST_0_i_1_n_0 ),
        .O(dout[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF54FFFFFF540000)) 
    \dout[7]_INST_0_i_1 
       (.I0(\dout[15]_INST_0_i_9_n_0 ),
        .I1(\dout[15]_INST_0_i_8_n_0 ),
        .I2(\dout[15]_INST_0_i_7_n_0 ),
        .I3(\dout[15]_INST_0_i_6_n_0 ),
        .I4(\dout[15]_INST_0_i_11_n_0 ),
        .I5(\dout[7]_INST_0_i_2_n_0 ),
        .O(\dout[7]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55404040)) 
    \dout[7]_INST_0_i_10 
       (.I0(bw),
        .I1(\dout[4]_INST_0_i_43_n_4 ),
        .I2(\dout[15]_INST_0_i_20_n_0 ),
        .I3(\dout[4]_INST_0_i_44_n_4 ),
        .I4(\dout[15]_INST_0_i_31_n_0 ),
        .O(\dout[7]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h953F)) 
    \dout[7]_INST_0_i_11_rewire_rewire 
       (.I0(\dout[15]_INST_0_i_33_n_0 ),
        .I1(\dout[15]_INST_0_i_82_n_0 ),
        .I2(\dout[9]_INST_0_i_22_n_0 ),
        .I3(\dout[7]_INST_0_i_7_n_0 ),
        .O(\dout[4]_INST_0_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0C0C0CFF04000400)) 
    \dout[7]_INST_0_i_12 
       (.I0(\dout[15]_INST_0_i_11_n_0 ),
        .I1(doc[0]),
        .I2(\dout[15]_INST_0_i_37_n_0 ),
        .I3(\dout[15]_INST_0_i_33_n_0 ),
        .I4(\dout[2]_INST_0_i_42_n_0 ),
        .I5(\dout[9]_INST_0_i_22_n_0_repN ),
        .O(\dout[7]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0400)) 
    \dout[7]_INST_0_i_13_rewire 
       (.I0(\dout[5]_INST_0_i_11_n_0 ),
        .I1(\dout[14]_INST_0_i_23_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .I3(\dout[5]_INST_0_i_5_n_0 ),
        .O(\dout[7]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h8E)) 
    \dout[7]_INST_0_i_14 
       (.I0(\dout[6]_INST_0_i_14_n_0 ),
        .I1(\dout[4]_INST_0_i_40_n_0 ),
        .I2(\dout[6]_INST_0_i_13_n_0 ),
        .O(\dout[7]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFEFEFEFEFEFEFE)) 
    \dout[7]_INST_0_i_2 
       (.I0(\dout[7]_INST_0_i_3_n_0 ),
        .I1(\dout[7]_INST_0_i_4_n_0 ),
        .I2(\dout[7]_INST_0_i_5_n_0 ),
        .I3(\dout[7]_INST_0_i_6_n_0 ),
        .I4(\dout[7]_INST_0_i_7_n_0_repN ),
        .I5(nstate1),
        .O(\dout[7]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \dout[7]_INST_0_i_3 
       (.I0(\dout[15]_INST_0_i_14_n_0 ),
        .I1(\dout[7]_INST_0_i_7_n_0_repN ),
        .I2(\dout[4]_INST_0_i_8_n_4 ),
        .I3(eqOp93_in),
        .I4(\dout[4]_INST_0_i_6_n_4 ),
        .I5(\dout[4]_INST_0_i_7_n_0 ),
        .O(\dout[7]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \dout[7]_INST_0_i_4 
       (.I0(\dout[7]_INST_0_i_8_n_0 ),
        .I1(\dout[7]_INST_0_i_9_n_0 ),
        .I2(\dout[15]_INST_0_i_23_n_0 ),
        .I3(\dout[7]_INST_0_i_10_n_0 ),
        .I4(\dout[4]_INST_0_i_11_n_4 ),
        .I5(\dout[15]_INST_0_i_19_n_0 ),
        .O(\dout[7]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000005000300050)) 
    \dout[7]_INST_0_i_5 
       (.I0(\dout[9]_INST_0_i_11_n_0 ),
        .I1(soc[1]),
        .I2(eqOp135_in),
        .I3(soc[2]),
        .I4(soc[0]),
        .I5(\dout[15]_INST_0_i_15_n_0 ),
        .O(\dout[7]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAA8A8AAAA08A80)) 
    \dout[7]_INST_0_i_6 
       (.I0(eqOp135_in),
        .I1(din[9]),
        .I2(p_2_in88_in),
        .I3(r_code[9]),
        .I4(din[7]),
        .I5(r_code[7]),
        .O(\dout[7]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "dout[7]_INST_0_i_7" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[7]_INST_0_i_7_replica 
       (.I0(\dout[15]_INST_0_i_33_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[7]_INST_0_i_7_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \dout[7]_INST_0_i_7_rewire 
       (.I0(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[7]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF444)) 
    \dout[7]_INST_0_i_8 
       (.I0(\dout[4]_INST_0_i_39_n_0 ),
        .I1(\dout[14]_INST_0_i_10_n_0 ),
        .I2(\dout[14]_INST_0_i_11_n_0 ),
        .I3(\dout[9]_INST_0_i_19_n_0 ),
        .I4(\dout[7]_INST_0_i_12_n_0 ),
        .O(\dout[7]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000AA695569)) 
    \dout[7]_INST_0_i_9 
       (.I0(\dout[4]_INST_0_i_39_n_0 ),
        .I1(\dout[7]_INST_0_i_13_n_0 ),
        .I2(\dout[7]_INST_0_i_14_n_0 ),
        .I3(\dout[9]_INST_0_i_12_n_0 ),
        .I4(\dout[9]_INST_0_i_23_n_0 ),
        .I5(bw),
        .O(\dout[7]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[8]_INST_0 
       (.I0(pc[8]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[8] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[8]_INST_0_i_1_n_0 ),
        .O(dout[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00A2)) 
    \dout[8]_INST_0_i_1 
       (.I0(\dout[8]_INST_0_i_2_n_0 ),
        .I1(\dout[13]_INST_0_i_3_n_0 ),
        .I2(\dout[8]_INST_0_i_3_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[8]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \dout[8]_INST_0_i_10 
       (.I0(\dout[15]_INST_0_i_20_n_0 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_39_n_7 ),
        .O(\dout[8]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABAAABBB)) 
    \dout[8]_INST_0_i_11 
       (.I0(\dout[15]_INST_0_i_37_n_0 ),
        .I1(\dout[9]_INST_0_i_11_n_0 ),
        .I2(din[12]),
        .I3(p_2_in88_in),
        .I4(r_code[12]),
        .O(\dout[8]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB800B800B800)) 
    \dout[8]_INST_0_i_12 
       (.I0(\dout[15]_INST_0_i_66_n_7 ),
        .I1(bw),
        .I2(\dout[15]_INST_0_i_71_n_7 ),
        .I3(\dout[15]_INST_0_i_31_n_0 ),
        .I4(\dout[4]_INST_0_i_7_n_0 ),
        .I5(\dout[15]_INST_0_i_61_n_7 ),
        .O(\dout[8]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \dout[8]_INST_0_i_13 
       (.I0(\dout[15]_INST_0_i_11_n_0 ),
        .I1(\dout[9]_INST_0_i_18_n_0 ),
        .O(\dout[2]_INST_0_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFBBBBABAA)) 
    \dout[8]_INST_0_i_2_rewire 
       (.I0(\dout[8]_INST_0_i_12_n_0 ),
        .I1(\dout[8]_INST_0_i_4_n_0 ),
        .I2(\dout[8]_INST_0_i_5_n_0 ),
        .I3(\dout[15]_INST_0_i_23_n_0 ),
        .I4(\dout[8]_INST_0_i_6_n_0 ),
        .I5(\dout[8]_INST_0_i_7_n_0 ),
        .O(\dout[8]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF8)) 
    \dout[8]_INST_0_i_3 
       (.I0(eqOp93_in),
        .I1(\dout[11]_INST_0_i_8_n_7 ),
        .I2(\dout[8]_INST_0_i_8_n_0 ),
        .I3(\dout[8]_INST_0_i_9_n_0 ),
        .O(\dout[8]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F444FFF44444444)) 
    \dout[8]_INST_0_i_4 
       (.I0(\dout[15]_INST_0_i_39_n_7 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_51_n_7 ),
        .I3(bw),
        .I4(\dout[15]_INST_0_i_56_n_7 ),
        .I5(\dout[15]_INST_0_i_20_n_0 ),
        .O(\dout[8]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h959A6A65)) 
    \dout[8]_INST_0_i_5 
       (.I0(L[8]),
        .I1(sr_reg_n_0_),
        .I2(bw),
        .I3(\dout[9]_INST_0_i_12_n_0 ),
        .I4(\dout[9]_INST_0_i_11_n_0 ),
        .O(\dout[8]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFAFCF0FAFFFFF0FF)) 
    \dout[8]_INST_0_i_6 
       (.I0(\dout[14]_INST_0_i_10_n_0 ),
        .I1(\dout[14]_INST_0_i_11_n_0 ),
        .I2(\dout[8]_INST_0_i_10_n_0 ),
        .I3(\dout[9]_INST_0_i_11_n_0 ),
        .I4(L[8]),
        .I5(\dout[8]_INST_0_i_11_n_0 ),
        .O(\dout[8]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAE)) 
    \dout[8]_INST_0_i_7_rewire 
       (.I0(\dout[8]_INST_0_i_3_n_0 ),
        .I1(\dout[15]_INST_0_i_14_n_0 ),
        .I2(\dout[9]_INST_0_i_11_n_0 ),
        .O(\dout[8]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000005000300050)) 
    \dout[8]_INST_0_i_8 
       (.I0(\dout[9]_INST_0_i_14_n_0 ),
        .I1(soc[1]),
        .I2(eqOp135_in),
        .I3(soc[2]),
        .I4(soc[0]),
        .I5(\dout[2]_INST_0_i_45_n_0 ),
        .O(\dout[8]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCC80CC8000000C00)) 
    \dout[8]_INST_0_i_9 
       (.I0(soc[0]),
        .I1(eqOp135_in),
        .I2(soc[1]),
        .I3(soc[2]),
        .I4(\dout[9]_INST_0_i_11_n_0 ),
        .I5(\dout[13]_INST_0_i_21_n_0 ),
        .O(\dout[8]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \dout[9]_INST_0 
       (.I0(pc[9]),
        .I1(\dout[15]_INST_0_i_1_n_0 ),
        .I2(\sr_reg_n_0_[9] ),
        .I3(\dout[15]_INST_0_i_2_n_0 ),
        .I4(\dout[9]_INST_0_i_1_n_0 ),
        .O(dout[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCC80CC8000000C00)) 
    \dout[9]_INST_0_i_10 
       (.I0(soc[0]),
        .I1(eqOp135_in),
        .I2(soc[1]),
        .I3(soc[2]),
        .I4(\dout[9]_INST_0_i_14_n_0 ),
        .I5(\dout[13]_INST_0_i_21_n_0 ),
        .O(\dout[9]_INST_0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00F4F4)) 
    \dout[9]_INST_0_i_11 
       (.I0(\rrs[0] [8]),
        .I1(\FSM_sequential_state[1]_i_12_n_0 ),
        .I2(\dout[9]_INST_0_i_17_n_0 ),
        .I3(\dout[9]_INST_0_i_18_n_0 ),
        .I4(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[9]_INST_0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000C550404FF)) 
    \dout[9]_INST_0_i_12 
       (.I0(\dout[9]_INST_0_i_19_n_0 ),
        .I1(\dout[9]_INST_0_i_20_n_0 ),
        .I2(\dout[9]_INST_0_i_21_n_0 ),
        .I3(\dout[7]_INST_0_i_7_n_0_repN ),
        .I4(\dout[9]_INST_0_i_22_n_0_repN ),
        .I5(\dout[9]_INST_0_i_23_n_0 ),
        .O(\dout[9]_INST_0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \dout[9]_INST_0_i_13 
       (.I0(\dout[15]_INST_0_i_20_n_0 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_39_n_6 ),
        .O(\dout[9]_INST_0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \dout[9]_INST_0_i_14 
       (.I0(\dout[0]_INST_0_i_10_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .I2(\dout[9]_INST_0_i_24_n_0 ),
        .O(\dout[9]_INST_0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABAAABBB)) 
    \dout[9]_INST_0_i_15 
       (.I0(\dout[15]_INST_0_i_37_n_0 ),
        .I1(\dout[9]_INST_0_i_14_n_0 ),
        .I2(din[12]),
        .I3(p_2_in88_in),
        .I4(r_code[12]),
        .O(\dout[9]_INST_0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFB800B800B800)) 
    \dout[9]_INST_0_i_16 
       (.I0(\dout[15]_INST_0_i_66_n_6 ),
        .I1(bw),
        .I2(\dout[15]_INST_0_i_71_n_6 ),
        .I3(\dout[15]_INST_0_i_31_n_0 ),
        .I4(\dout[4]_INST_0_i_7_n_0 ),
        .I5(\dout[15]_INST_0_i_61_n_6 ),
        .O(\dout[9]_INST_0_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0A3A3A3A0A0A0A0)) 
    \dout[9]_INST_0_i_17 
       (.I0(\addr[8]_INST_0_i_8_n_0 ),
        .I1(\FSM_sequential_state[1]_i_12_n_0 ),
        .I2(\dout[5]_INST_0_i_10_n_0 ),
        .I3(\dout[5]_INST_0_i_14_n_0 ),
        .I4(src__0[8]),
        .I5(\dout[9]_INST_0_i_25_n_0 ),
        .O(\dout[9]_INST_0_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1101F0001101FF0F)) 
    \dout[9]_INST_0_i_18 
       (.I0(lbe_INST_0_i_7_n_0),
        .I1(\dout[9]_INST_0_i_26_n_0 ),
        .I2(\dout[5]_INST_0_i_10_n_0 ),
        .I3(lbe_INST_0_i_11_n_0),
        .I4(\FSM_sequential_state[1]_i_12_n_0 ),
        .I5(\dout[9]_INST_0_i_27_n_0 ),
        .O(\dout[9]_INST_0_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \dout[9]_INST_0_i_19_rewire 
       (.I0(\dout[15]_INST_0_i_82_n_0 ),
        .I1(\dout[15]_INST_0_i_33_n_0 ),
        .I2(\dout[9]_INST_0_i_22_n_0 ),
        .O(\dout[9]_INST_0_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FEFE00FE)) 
    \dout[9]_INST_0_i_1_rewire_rewire 
       (.I0(\dout[9]_INST_0_i_16_n_0 ),
        .I1(\dout[9]_INST_0_i_8_n_0 ),
        .I2(\dout[9]_INST_0_i_2_n_0 ),
        .I3(\dout[13]_INST_0_i_3_n_0 ),
        .I4(\dout[9]_INST_0_i_3_n_0 ),
        .I5(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[9]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555665666666666)) 
    \dout[9]_INST_0_i_20 
       (.I0(\dout[4]_INST_0_i_40_n_0 ),
        .I1(\dout[6]_INST_0_i_13_n_0 ),
        .I2(\dout[4]_INST_0_i_35_n_0 ),
        .I3(\dout[9]_INST_0_i_28_n_0 ),
        .I4(\dout[4]_INST_0_i_32_n_0 ),
        .I5(\dout[9]_INST_0_i_29_n_0 ),
        .O(\dout[9]_INST_0_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9999999696969696)) 
    \dout[9]_INST_0_i_21 
       (.I0(\dout[5]_INST_0_i_12_n_0_repN ),
        .I1(\dout[13]_INST_0_i_20_n_0_repN ),
        .I2(\dout[4]_INST_0_i_32_n_0 ),
        .I3(\dout[4]_INST_0_i_20_n_0 ),
        .I4(\dout[4]_INST_0_i_5_n_0 ),
        .I5(\dout[4]_INST_0_i_35_n_0 ),
        .O(\dout[9]_INST_0_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "dout[9]_INST_0_i_22" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \dout[9]_INST_0_i_22_replica 
       (.I0(\dout[15]_INST_0_i_82_n_0 ),
        .I1(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[9]_INST_0_i_22_n_0_repN ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \dout[9]_INST_0_i_22_rewire 
       (.I0(\dout[15]_INST_0_i_11_n_0 ),
        .O(\dout[9]_INST_0_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAA8888AAA8)) 
    \dout[9]_INST_0_i_23 
       (.I0(\dout[9]_INST_0_i_30_n_0 ),
        .I1(\dout[7]_INST_0_i_13_n_0 ),
        .I2(\dout[5]_INST_0_i_12_n_0_repN ),
        .I3(\dout[13]_INST_0_i_20_n_0_repN ),
        .I4(\dout[9]_INST_0_i_31_n_0 ),
        .I5(\dout[6]_INST_0_i_13_n_0 ),
        .O(\dout[9]_INST_0_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00F3E2E2)) 
    \dout[9]_INST_0_i_24 
       (.I0(\dout[9]_INST_0_i_32_n_0 ),
        .I1(\dout[5]_INST_0_i_10_n_0 ),
        .I2(\addr[9]_INST_0_i_8_n_0 ),
        .I3(\rrs[0] [9]),
        .I4(\FSM_sequential_state[1]_i_12_n_0 ),
        .O(\dout[9]_INST_0_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7774747477777777)) 
    \dout[9]_INST_0_i_25 
       (.I0(soc[0]),
        .I1(eqOp93_in),
        .I2(\dout[5]_INST_0_i_14_n_0 ),
        .I3(bw),
        .I4(r_a0),
        .I5(din[8]),
        .O(\dout[9]_INST_0_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0880088AA880A88)) 
    \dout[9]_INST_0_i_26 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(\dout[11]_INST_0_i_42_n_0 ),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(as[0]),
        .I5(lbe_INST_0_i_23_n_0),
        .O(\dout[9]_INST_0_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000800080008FFFB)) 
    \dout[9]_INST_0_i_27 
       (.I0(src__0[0]),
        .I1(rd_INST_0_i_21_n_0),
        .I2(rd_INST_0_i_16_n_0),
        .I3(\dout[13]_INST_0_i_3_n_0 ),
        .I4(eqOp93_in),
        .I5(\dout[11]_INST_0_i_41_n_0 ),
        .O(\dout[9]_INST_0_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3233)) 
    \dout[9]_INST_0_i_28_rewire 
       (.I0(\dout[3]_INST_0_i_10_n_0 ),
        .I1(\dout[4]_INST_0_i_20_n_0 ),
        .I2(\dout[15]_INST_0_i_11_n_0 ),
        .I3(\dout[3]_INST_0_i_5_n_0 ),
        .O(\dout[9]_INST_0_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00F700F0)) 
    \dout[9]_INST_0_i_29_rewire_rewire 
       (.I0(\dout[5]_INST_0_i_15_n_0 ),
        .I1(\dout[4]_INST_0_i_46_n_0 ),
        .I2(\dout[15]_INST_0_i_84_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .I4(\dout[4]_INST_0_i_16_n_0 ),
        .O(\dout[9]_INST_0_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0F0F0900)) 
    \dout[9]_INST_0_i_2_rewire 
       (.I0(\dout[9]_INST_0_i_4_n_0 ),
        .I1(\dout[9]_INST_0_i_5_n_0 ),
        .I2(\dout[9]_INST_0_i_6_n_0 ),
        .I3(\dout[15]_INST_0_i_23_n_0 ),
        .I4(\dout[9]_INST_0_i_7_n_0 ),
        .O(\dout[9]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF8)) 
    \dout[9]_INST_0_i_3 
       (.I0(eqOp93_in),
        .I1(\dout[11]_INST_0_i_8_n_6 ),
        .I2(\dout[9]_INST_0_i_9_n_0 ),
        .I3(\dout[9]_INST_0_i_10_n_0 ),
        .O(\dout[9]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h44F400F0)) 
    \dout[9]_INST_0_i_30_rewire_rewire 
       (.I0(\dout[5]_INST_0_i_11_n_0 ),
        .I1(\dout[5]_INST_0_i_5_n_0 ),
        .I2(\dout[14]_INST_0_i_23_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .I4(\dout[6]_INST_0_i_7_n_0 ),
        .O(\dout[9]_INST_0_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5501555501010101)) 
    \dout[9]_INST_0_i_31 
       (.I0(\dout[4]_INST_0_i_32_n_0 ),
        .I1(\dout[4]_INST_0_i_20_n_0 ),
        .I2(\dout[4]_INST_0_i_5_n_0 ),
        .I3(\dout[4]_INST_0_i_47_n_0 ),
        .I4(\dout[3]_INST_0_i_12_n_0 ),
        .I5(\dout[9]_INST_0_i_33_n_0 ),
        .O(\dout[9]_INST_0_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000477777774777)) 
    \dout[9]_INST_0_i_32 
       (.I0(soc[1]),
        .I1(eqOp93_in),
        .I2(din[9]),
        .I3(\dout[15]_INST_0_i_109_n_0 ),
        .I4(\dout[5]_INST_0_i_14_n_0 ),
        .I5(src__0[9]),
        .O(\dout[9]_INST_0_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FF717371FFFF)) 
    \dout[9]_INST_0_i_33 
       (.I0(\dout[4]_INST_0_i_61_n_0 ),
        .I1(\dout[2]_INST_0_i_15_n_0 ),
        .I2(\dout[1]_INST_0_i_5_n_0 ),
        .I3(\dout[15]_INST_0_i_11_n_0 ),
        .I4(\dout[2]_INST_0_i_14_n_0 ),
        .I5(\dout[2]_INST_0_i_13_n_0 ),
        .O(\dout[9]_INST_0_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6565A665A6A6A665)) 
    \dout[9]_INST_0_i_4 
       (.I0(\dout[15]_INST_0_i_80_n_0 ),
        .I1(L[8]),
        .I2(\dout[9]_INST_0_i_11_n_0 ),
        .I3(\dout[9]_INST_0_i_12_n_0 ),
        .I4(bw),
        .I5(sr_reg_n_0_),
        .O(\dout[9]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFDF4DCFDFFFCFDF)) 
    \dout[9]_INST_0_i_5 
       (.I0(\dout[9]_INST_0_i_4_n_0 ),
        .I1(L[11]),
        .I2(\dout[11]_INST_0_i_16_n_0 ),
        .I3(\dout[11]_INST_0_i_14_n_0 ),
        .I4(L[10]),
        .I5(\dout[2]_INST_0_i_12_n_0 ),
        .O(\dout[9]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F444FFF44444444)) 
    \dout[9]_INST_0_i_6 
       (.I0(\dout[15]_INST_0_i_39_n_6 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_51_n_6 ),
        .I3(bw),
        .I4(\dout[15]_INST_0_i_56_n_6 ),
        .I5(\dout[15]_INST_0_i_20_n_0 ),
        .O(\dout[9]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFAFCF0FAFFFFF0FF)) 
    \dout[9]_INST_0_i_7 
       (.I0(\dout[14]_INST_0_i_10_n_0 ),
        .I1(\dout[14]_INST_0_i_11_n_0 ),
        .I2(\dout[9]_INST_0_i_13_n_0 ),
        .I3(\dout[9]_INST_0_i_14_n_0 ),
        .I4(L[9]),
        .I5(\dout[9]_INST_0_i_15_n_0 ),
        .O(\dout[9]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAE)) 
    \dout[9]_INST_0_i_8_rewire 
       (.I0(\dout[9]_INST_0_i_3_n_0 ),
        .I1(\dout[15]_INST_0_i_14_n_0 ),
        .I2(\dout[9]_INST_0_i_14_n_0 ),
        .O(\dout[9]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0030005000000050)) 
    \dout[9]_INST_0_i_9 
       (.I0(\dout[2]_INST_0_i_12_n_0 ),
        .I1(soc[1]),
        .I2(eqOp135_in),
        .I3(soc[2]),
        .I4(soc[0]),
        .I5(\dout[0]_INST_0_i_5_n_0 ),
        .O(\dout[9]_INST_0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBABB)) 
    hbe_INST_0
       (.I0(lbe_INST_0_i_4_n_0),
        .I1(lbe_INST_0_i_1_n_0),
        .I2(lbe_INST_0_i_3_n_0),
        .I3(bw),
        .O(hbe));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8FFF0F008000000)) 
    \iack[0]_i_1 
       (.I0(\iack[0]_i_2_n_0 ),
        .I1(\iack[8]_i_2_n_0 ),
        .I2(halt),
        .I3(\iack[0]_i_3_n_0 ),
        .I4(\iack[14]_i_4_n_0 ),
        .I5(iack[0]),
        .O(\iack[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \iack[0]_i_2 
       (.I0(irq[1]),
        .I1(irq[2]),
        .I2(irq[3]),
        .I3(irq[0]),
        .I4(\irqaddr[3]_i_2_n_0 ),
        .I5(irq[8]),
        .O(\iack[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \iack[0]_i_3 
       (.I0(\irqaddr[4]_i_2_n_0 ),
        .I1(\irqaddr[3]_i_2_n_0 ),
        .I2(irq[0]),
        .I3(irq[3]),
        .I4(irq[2]),
        .I5(irq[1]),
        .O(\iack[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFAAAA00400000)) 
    \iack[10]_i_1 
       (.I0(halt),
        .I1(\iack[11]_i_2_n_0 ),
        .I2(irq[10]),
        .I3(irq[11]),
        .I4(\iack[14]_i_4_n_0 ),
        .I5(iack[10]),
        .O(\iack[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFAA4000)) 
    \iack[11]_i_1 
       (.I0(halt),
        .I1(\iack[11]_i_2_n_0 ),
        .I2(irq[11]),
        .I3(\iack[14]_i_4_n_0 ),
        .I4(iack[11]),
        .O(\iack[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \iack[11]_i_2 
       (.I0(irq[13]),
        .I1(irq[12]),
        .I2(irq[14]),
        .O(\iack[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFAAAA00040000)) 
    \iack[12]_i_1 
       (.I0(halt),
        .I1(irq[12]),
        .I2(irq[14]),
        .I3(irq[13]),
        .I4(\iack[14]_i_4_n_0 ),
        .I5(iack[12]),
        .O(\iack[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFAA0400)) 
    \iack[13]_i_1 
       (.I0(halt),
        .I1(irq[13]),
        .I2(irq[14]),
        .I3(\iack[14]_i_4_n_0 ),
        .I4(iack[13]),
        .O(\iack[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFEC2020)) 
    \iack[14]_i_1 
       (.I0(\iack[14]_i_3_n_0 ),
        .I1(halt),
        .I2(irq[14]),
        .I3(\iack[14]_i_4_n_0 ),
        .I4(iack[14]),
        .O(\iack[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \iack[14]_i_2 
       (.I0(rst),
        .O(\iack[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000020)) 
    \iack[14]_i_3 
       (.I0(state[0]),
        .I1(state[1]),
        .I2(state[2]),
        .I3(state[4]),
        .I4(state[3]),
        .O(\iack[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \iack[14]_i_4 
       (.I0(state[3]),
        .I1(state[4]),
        .I2(state[2]),
        .I3(state[1]),
        .I4(state[0]),
        .I5(girq),
        .O(\iack[14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEFFAAAAAAAA)) 
    \iack[14]_i_5 
       (.I0(irq[14]),
        .I1(irq[4]),
        .I2(irq[0]),
        .I3(\iack[14]_i_6_n_0 ),
        .I4(\iack[14]_i_7_n_0 ),
        .I5(p_1_in108_in),
        .O(girq));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \iack[14]_i_6 
       (.I0(irq[1]),
        .I1(irq[2]),
        .I2(irq[3]),
        .O(\iack[14]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFFFFFFFFFF)) 
    \iack[14]_i_7 
       (.I0(irq[8]),
        .I1(irq[5]),
        .I2(irq[9]),
        .I3(\iack[14]_i_8_n_0 ),
        .I4(\iack[5]_i_2_n_0 ),
        .I5(\iack[9]_i_2_n_0 ),
        .O(\iack[14]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \iack[14]_i_8 
       (.I0(irq[12]),
        .I1(irq[13]),
        .O(\iack[14]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFA40)) 
    \iack[1]_i_1 
       (.I0(halt),
        .I1(\iack[1]_i_2_n_0 ),
        .I2(\iack[14]_i_4_n_0 ),
        .I3(iack[1]),
        .O(\iack[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000020)) 
    \iack[1]_i_2 
       (.I0(\iack[4]_i_2_n_0 ),
        .I1(irq[4]),
        .I2(irq[1]),
        .I3(irq[2]),
        .I4(irq[3]),
        .O(\iack[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFA40)) 
    \iack[2]_i_1 
       (.I0(halt),
        .I1(\iack[2]_i_2_n_0 ),
        .I2(\iack[14]_i_4_n_0 ),
        .I3(iack[2]),
        .O(\iack[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \iack[2]_i_2 
       (.I0(\irqaddr[4]_i_2_n_0 ),
        .I1(irq[7]),
        .I2(irq[3]),
        .I3(irq[2]),
        .I4(irq[6]),
        .I5(\iack[2]_i_3_n_0 ),
        .O(\iack[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \iack[2]_i_3 
       (.I0(irq[4]),
        .I1(irq[5]),
        .O(\iack[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8FFF0F008000000)) 
    \iack[3]_i_1 
       (.I0(\iack[3]_i_2_n_0 ),
        .I1(\iack[4]_i_2_n_0 ),
        .I2(halt),
        .I3(\iack[3]_i_3_n_0 ),
        .I4(\iack[14]_i_4_n_0 ),
        .I5(iack[3]),
        .O(\iack[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \iack[3]_i_2 
       (.I0(irq[3]),
        .I1(irq[4]),
        .O(\iack[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \iack[3]_i_3 
       (.I0(\irqaddr[4]_i_2_n_0 ),
        .I1(irq[6]),
        .I2(irq[7]),
        .I3(irq[5]),
        .I4(irq[3]),
        .I5(irq[4]),
        .O(\iack[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFAA4000)) 
    \iack[4]_i_1 
       (.I0(halt),
        .I1(\iack[4]_i_2_n_0 ),
        .I2(irq[4]),
        .I3(\iack[14]_i_4_n_0 ),
        .I4(iack[4]),
        .O(\iack[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000002)) 
    \iack[4]_i_2 
       (.I0(\iack[8]_i_2_n_0 ),
        .I1(irq[7]),
        .I2(irq[6]),
        .I3(irq[8]),
        .I4(irq[5]),
        .O(\iack[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFAAAA10000000)) 
    \iack[5]_i_1 
       (.I0(halt),
        .I1(\irqaddr[4]_i_2_n_0 ),
        .I2(\iack[5]_i_2_n_0 ),
        .I3(irq[5]),
        .I4(\iack[14]_i_4_n_0 ),
        .I5(iack[5]),
        .O(\iack[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \iack[5]_i_2 
       (.I0(irq[7]),
        .I1(irq[6]),
        .O(\iack[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFAAAA00040000)) 
    \iack[6]_i_1 
       (.I0(halt),
        .I1(irq[6]),
        .I2(\irqaddr[4]_i_2_n_0 ),
        .I3(irq[7]),
        .I4(\iack[14]_i_4_n_0 ),
        .I5(iack[6]),
        .O(\iack[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFAA0400)) 
    \iack[7]_i_1 
       (.I0(halt),
        .I1(irq[7]),
        .I2(\irqaddr[4]_i_2_n_0 ),
        .I3(\iack[14]_i_4_n_0 ),
        .I4(iack[7]),
        .O(\iack[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFAA4000)) 
    \iack[8]_i_1 
       (.I0(halt),
        .I1(\iack[8]_i_2_n_0 ),
        .I2(irq[8]),
        .I3(\iack[14]_i_4_n_0 ),
        .I4(iack[8]),
        .O(\iack[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \iack[8]_i_2 
       (.I0(irq[14]),
        .I1(irq[12]),
        .I2(irq[13]),
        .I3(irq[11]),
        .I4(irq[10]),
        .I5(irq[9]),
        .O(\iack[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFAAAA40000000)) 
    \iack[9]_i_1 
       (.I0(halt),
        .I1(\iack[11]_i_2_n_0 ),
        .I2(\iack[9]_i_2_n_0 ),
        .I3(irq[9]),
        .I4(\iack[14]_i_4_n_0 ),
        .I5(iack[9]),
        .O(\iack[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \iack[9]_i_2 
       (.I0(irq[11]),
        .I1(irq[10]),
        .O(\iack[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[0]_i_1_n_0 ),
        .Q(iack[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[10]_i_1_n_0 ),
        .Q(iack[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[11]_i_1_n_0 ),
        .Q(iack[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[12]_i_1_n_0 ),
        .Q(iack[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[13]_i_1_n_0 ),
        .Q(iack[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[14]_i_1_n_0 ),
        .Q(iack[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[1]_i_1_n_0 ),
        .Q(iack[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[2]_i_1_n_0 ),
        .Q(iack[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[3]_i_1_n_0 ),
        .Q(iack[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[4]_i_1_n_0 ),
        .Q(iack[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[5]_i_1_n_0 ),
        .Q(iack[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[6]_i_1_n_0 ),
        .Q(iack[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[7]_i_1_n_0 ),
        .Q(iack[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[8]_i_1_n_0 ),
        .Q(iack[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \iack_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\iack[14]_i_2_n_0 ),
        .D(\iack[9]_i_1_n_0 ),
        .Q(iack[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00AB)) 
    \irqaddr[1]_i_1 
       (.I0(irq[13]),
        .I1(\irqaddr[1]_i_2_n_0 ),
        .I2(irq[12]),
        .I3(irq[14]),
        .O(\irqaddr[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4545454544444544)) 
    \irqaddr[1]_i_2 
       (.I0(irq[11]),
        .I1(irq[10]),
        .I2(irq[9]),
        .I3(\irqaddr[1]_i_3_n_0 ),
        .I4(irq[7]),
        .I5(irq[8]),
        .O(\irqaddr[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAEEEEAAAAFFEF)) 
    \irqaddr[1]_i_3 
       (.I0(irq[6]),
        .I1(irq[4]),
        .I2(irq[1]),
        .I3(irq[2]),
        .I4(irq[5]),
        .I5(irq[3]),
        .O(\irqaddr[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAABBAAAAAAFB)) 
    \irqaddr[2]_i_1 
       (.I0(irq[14]),
        .I1(\iack[9]_i_2_n_0 ),
        .I2(\irqaddr[2]_i_2_n_0 ),
        .I3(irq[13]),
        .I4(irq[12]),
        .I5(irq[9]),
        .O(\irqaddr[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000005455555555)) 
    \irqaddr[2]_i_2 
       (.I0(irq[8]),
        .I1(irq[2]),
        .I2(irq[3]),
        .I3(irq[5]),
        .I4(irq[4]),
        .I5(\iack[5]_i_2_n_0 ),
        .O(\irqaddr[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555555555555557)) 
    \irqaddr[3]_i_1 
       (.I0(\iack[11]_i_2_n_0 ),
        .I1(irq[8]),
        .I2(irq[11]),
        .I3(irq[10]),
        .I4(irq[9]),
        .I5(\irqaddr[3]_i_2_n_0 ),
        .O(\irqaddr[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \irqaddr[3]_i_2 
       (.I0(irq[6]),
        .I1(irq[7]),
        .I2(irq[5]),
        .I3(irq[4]),
        .O(\irqaddr[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \irqaddr[4]_i_1 
       (.I0(\iack[14]_i_4_n_0 ),
        .I1(halt),
        .O(irqaddr0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFD)) 
    \irqaddr[4]_i_2 
       (.I0(\iack[11]_i_2_n_0 ),
        .I1(irq[9]),
        .I2(irq[10]),
        .I3(irq[11]),
        .I4(irq[8]),
        .O(\irqaddr[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \irqaddr_reg[1] 
       (.C(clk),
        .CE(irqaddr0),
        .D(\irqaddr[1]_i_1_n_0 ),
        .PRE(\iack[14]_i_2_n_0 ),
        .Q(irqaddr[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \irqaddr_reg[2] 
       (.C(clk),
        .CE(irqaddr0),
        .D(\irqaddr[2]_i_1_n_0 ),
        .PRE(\iack[14]_i_2_n_0 ),
        .Q(irqaddr[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \irqaddr_reg[3] 
       (.C(clk),
        .CE(irqaddr0),
        .D(\irqaddr[3]_i_1_n_0 ),
        .PRE(\iack[14]_i_2_n_0 ),
        .Q(irqaddr[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \irqaddr_reg[4] 
       (.C(clk),
        .CE(irqaddr0),
        .D(\irqaddr[4]_i_2_n_0 ),
        .PRE(\iack[14]_i_2_n_0 ),
        .Q(irqaddr[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF15)) 
    lbe_INST_0
       (.I0(lbe_INST_0_i_1_n_0),
        .I1(bw),
        .I2(lbe_INST_0_i_3_n_0),
        .I3(lbe_INST_0_i_4_n_0),
        .O(lbe));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5455555555515455)) 
    lbe_INST_0_i_1
       (.I0(rd_INST_0_i_1_n_0),
        .I1(state[0]),
        .I2(state[4]),
        .I3(state[3]),
        .I4(state[1]),
        .I5(state[2]),
        .O(lbe_INST_0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    lbe_INST_0_i_10
       (.I0(lbe_INST_0_i_18_n_0),
        .I1(\addr[15]_INST_0_i_31_n_0 ),
        .I2(plusOp3_out[0]),
        .I3(state[0]),
        .I4(plusOp4_out[0]),
        .O(lbe_INST_0_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFCFAFC0A0CFA0C0)) 
    lbe_INST_0_i_11
       (.I0(lbe_INST_0_i_19_n_0),
        .I1(lbe_INST_0_i_20_n_0),
        .I2(\r_code[11]_i_1_n_0 ),
        .I3(\r_code[10]_i_1_n_0 ),
        .I4(lbe_INST_0_i_21_n_0),
        .I5(lbe_INST_0_i_22_n_0),
        .O(lbe_INST_0_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00A000FC00A0000C)) 
    lbe_INST_0_i_12
       (.I0(\r_reg[7] [0]),
        .I1(\r_reg[4] [0]),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_9_n_0 ),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_reg[6] [0]),
        .O(lbe_INST_0_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABAAAAAA)) 
    lbe_INST_0_i_13
       (.I0(\r_code[3]_i_1_n_0 ),
        .I1(\addr[3]_INST_0_i_9_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_code[0]_i_1_n_0 ),
        .I4(\r_reg[5] [0]),
        .O(lbe_INST_0_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0C080008)) 
    lbe_INST_0_i_14
       (.I0(\r_reg[14] [0]),
        .I1(\r_code[1]_i_1_n_0 ),
        .I2(\addr[3]_INST_0_i_9_n_0 ),
        .I3(\r_code[0]_i_1_n_0 ),
        .I4(\r_reg[15] [0]),
        .O(lbe_INST_0_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h22200200FFFFFFFF)) 
    lbe_INST_0_i_15
       (.I0(\addr[3]_INST_0_i_9_n_0_repN ),
        .I1(\r_code[1]_i_1_n_0 ),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(\r_reg[8] [0]),
        .I4(\r_reg[9] [0]),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(lbe_INST_0_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF4FFF7)) 
    lbe_INST_0_i_16
       (.I0(\r_reg[13] [0]),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\addr[3]_INST_0_i_9_n_0 ),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(\r_reg[12] [0]),
        .O(lbe_INST_0_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAC000000)) 
    lbe_INST_0_i_17
       (.I0(\r_reg[11] [0]),
        .I1(\r_reg[10] [0]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_9_n_0 ),
        .I4(\r_code[1]_i_1_n_0 ),
        .O(lbe_INST_0_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    lbe_INST_0_i_18
       (.I0(\addr[3]_INST_0_i_23_n_7 ),
        .I1(p_4_in),
        .I2(pc[0]),
        .I3(\addr[15]_INST_0_i_40_n_0 ),
        .I4(plusOp2_out[0]),
        .O(lbe_INST_0_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    lbe_INST_0_i_19
       (.I0(\r_reg[15] [0]),
        .I1(\r_reg[14] [0]),
        .I2(soc[2]),
        .I3(\r_reg[13] [0]),
        .I4(soc[1]),
        .I5(\r_reg[12] [0]),
        .O(lbe_INST_0_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    lbe_INST_0_i_2
       (.I0(din[6]),
        .I1(p_2_in88_in),
        .I2(r_code[6]),
        .O(bw));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    lbe_INST_0_i_20
       (.I0(\r_reg[11] [0]),
        .I1(\r_reg[10] [0]),
        .I2(soc[2]),
        .I3(\r_reg[9] [0]),
        .I4(soc[1]),
        .I5(\r_reg[8] [0]),
        .O(lbe_INST_0_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3A003A0F3AF03AFF)) 
    lbe_INST_0_i_21
       (.I0(lbe_INST_0_i_23_n_0),
        .I1(as[0]),
        .I2(soc[1]),
        .I3(soc[2]),
        .I4(pc[0]),
        .I5(sp_reg[0]),
        .O(lbe_INST_0_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    lbe_INST_0_i_22
       (.I0(\r_reg[7] [0]),
        .I1(\r_reg[6] [0]),
        .I2(soc[2]),
        .I3(\r_reg[5] [0]),
        .I4(soc[1]),
        .I5(\r_reg[4] [0]),
        .O(lbe_INST_0_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFBBFCB8FFFFFFFF)) 
    lbe_INST_0_i_23
       (.I0(din[4]),
        .I1(p_2_in88_in),
        .I2(r_code[4]),
        .I3(din[5]),
        .I4(r_code[5]),
        .I5(sr_reg_n_0_),
        .O(lbe_INST_0_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFF4F44)) 
    lbe_INST_0_i_3
       (.I0(\addr[15]_INST_0_i_1_n_0 ),
        .I1(\rrs[0] [0]),
        .I2(\addr[15]_INST_0_i_3_n_0 ),
        .I3(sp_reg[0]),
        .I4(lbe_INST_0_i_6_n_0),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(lbe_INST_0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABEAAAAAAA)) 
    lbe_INST_0_i_4
       (.I0(rd_INST_0_i_2_n_0),
        .I1(state[2]),
        .I2(state[3]),
        .I3(state[0]),
        .I4(state[1]),
        .I5(state[4]),
        .O(lbe_INST_0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFAABAAAAAAAAA)) 
    lbe_INST_0_i_5
       (.I0(lbe_INST_0_i_7_n_0),
        .I1(lbe_INST_0_i_8_n_0),
        .I2(sr_reg_n_0_),
        .I3(\addr[15]_INST_0_i_8_n_0 ),
        .I4(lbe_INST_0_i_9_n_0),
        .I5(\addr[15]_INST_0_i_11_n_0 ),
        .O(\rrs[0] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000FFB8B8)) 
    lbe_INST_0_i_6
       (.I0(data3[0]),
        .I1(\addr[15]_INST_0_i_14_n_0 ),
        .I2(lbe_INST_0_i_10_n_0),
        .I3(lbe_INST_0_i_11_n_0),
        .I4(\addr[15]_INST_0_i_17_n_0 ),
        .I5(\addr[15]_INST_0_i_18_n_0 ),
        .O(lbe_INST_0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEEEEE0EEEE)) 
    lbe_INST_0_i_7
       (.I0(lbe_INST_0_i_12_n_0),
        .I1(lbe_INST_0_i_13_n_0),
        .I2(lbe_INST_0_i_14_n_0),
        .I3(lbe_INST_0_i_15_n_0),
        .I4(lbe_INST_0_i_16_n_0),
        .I5(lbe_INST_0_i_17_n_0),
        .O(lbe_INST_0_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFACCFA)) 
    lbe_INST_0_i_8
       (.I0(r_code[5]),
        .I1(din[5]),
        .I2(r_code[4]),
        .I3(p_2_in88_in),
        .I4(din[4]),
        .O(lbe_INST_0_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0AC00AC)) 
    lbe_INST_0_i_9
       (.I0(sp_reg[0]),
        .I1(pc[0]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(as[0]),
        .O(lbe_INST_0_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[0]_i_1 
       (.I0(din[0]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[3]_i_2_n_7 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[0]_INST_0_i_1_n_0 ),
        .O(\pc[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[10]_i_1 
       (.I0(din[10]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[11]_i_2_n_5 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[10]_INST_0_i_1_n_0 ),
        .O(\pc[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[11]_i_1 
       (.I0(din[11]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[11]_i_2_n_4 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[11]_INST_0_i_1_n_0 ),
        .O(\pc[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[12]_i_1 
       (.I0(din[12]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[15]_i_7_n_7 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[12]_INST_0_i_1_n_0 ),
        .O(\pc[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[13]_i_1 
       (.I0(din[13]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[15]_i_7_n_6 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[13]_INST_0_i_1_n_0 ),
        .O(\pc[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[14]_i_1 
       (.I0(din[14]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[15]_i_7_n_5 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[14]_INST_0_i_1_n_0 ),
        .O(\pc[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55545555)) 
    \pc[15]_i_1 
       (.I0(halt),
        .I1(\pc[15]_i_3_n_0 ),
        .I2(\pc[15]_i_4_n_0 ),
        .I3(rd_INST_0_i_10_n_0),
        .I4(\pc[15]_i_5_n_0 ),
        .O(\pc[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \pc[15]_i_10 
       (.I0(nstate1),
        .I1(soc[0]),
        .I2(state[1]),
        .I3(state[0]),
        .I4(rd_INST_0_i_37_n_0),
        .I5(state[2]),
        .O(\pc[15]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[15]_i_2 
       (.I0(din[15]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[15]_i_7_n_4 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[15]_INST_0_i_3_n_0 ),
        .O(\pc[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFF54FF54FF54)) 
    \pc[15]_i_3 
       (.I0(rd_INST_0_i_7_n_0),
        .I1(p_2_in88_in),
        .I2(rd_INST_0_i_18_n_0),
        .I3(\pc[15]_i_6_n_0 ),
        .I4(\pc[15]_i_8_n_0 ),
        .I5(\pc[15]_i_9_n_0 ),
        .O(\pc[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000002)) 
    \pc[15]_i_4 
       (.I0(\sp[0]_i_4_n_0 ),
        .I1(\r_code[11]_i_1_n_0 ),
        .I2(soc[2]),
        .I3(\r_code[10]_i_1_n_0 ),
        .I4(soc[1]),
        .O(\pc[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000DDD)) 
    \pc[15]_i_5 
       (.I0(\pc[15]_i_8_n_0 ),
        .I1(rd_INST_0_i_8_n_0),
        .I2(eqOp93_in),
        .I3(p_2_in88_in),
        .I4(\pc[15]_i_10_n_0 ),
        .O(\pc[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00024000)) 
    \pc[15]_i_6 
       (.I0(state[4]),
        .I1(state[2]),
        .I2(state[3]),
        .I3(state[0]),
        .I4(state[1]),
        .O(\pc[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \pc[15]_i_8 
       (.I0(\addr[15]_INST_0_i_11_n_0 ),
        .I1(\r_code[1]_i_1_n_0 ),
        .I2(\r_code[0]_i_1_n_0 ),
        .O(\pc[15]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000010010)) 
    \pc[15]_i_9 
       (.I0(state[1]),
        .I1(state[0]),
        .I2(state[2]),
        .I3(state[4]),
        .I4(state[3]),
        .I5(\addr[15]_INST_0_i_20_n_0 ),
        .O(\pc[15]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[1]_i_1 
       (.I0(din[1]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[3]_i_2_n_6 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[1]_INST_0_i_1_n_0 ),
        .O(\pc[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[2]_i_1 
       (.I0(din[2]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[3]_i_2_n_5 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[2]_INST_0_i_1_n_0 ),
        .O(\pc[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[3]_i_1 
       (.I0(din[3]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[3]_i_2_n_4 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[3]_INST_0_i_1_n_0 ),
        .O(\pc[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \pc[3]_i_5 
       (.I0(pc[1]),
        .O(\pc[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[4]_i_1 
       (.I0(din[4]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[7]_i_2_n_7 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[4]_INST_0_i_1_n_0 ),
        .O(\pc[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[5]_i_1 
       (.I0(din[5]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[7]_i_2_n_6 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[5]_INST_0_i_1_n_0 ),
        .O(\pc[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[6]_i_1 
       (.I0(din[6]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[7]_i_2_n_5 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[6]_INST_0_i_1_n_0 ),
        .O(\pc[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[7]_i_1 
       (.I0(din[7]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[7]_i_2_n_4 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[7]_INST_0_i_1_n_0 ),
        .O(\pc[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[8]_i_1 
       (.I0(din[8]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[11]_i_2_n_7 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[8]_INST_0_i_1_n_0 ),
        .O(\pc[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[9]_i_1 
       (.I0(din[9]),
        .I1(\pc[15]_i_6_n_0 ),
        .I2(\pc_reg[11]_i_2_n_6 ),
        .I3(\pc[15]_i_5_n_0 ),
        .I4(\dout[9]_INST_0_i_1_n_0 ),
        .O(\pc[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[0] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[0]_i_1_n_0 ),
        .Q(pc[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[10] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[10]_i_1_n_0 ),
        .Q(pc[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[11] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[11]_i_1_n_0 ),
        .Q(pc[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \pc_reg[11]_i_2 
       (.CI(\pc_reg[7]_i_2_n_0 ),
        .CO(pc_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\pc_reg[11]_i_2_n_4 ,\pc_reg[11]_i_2_n_5 ,\pc_reg[11]_i_2_n_6 ,\pc_reg[11]_i_2_n_7 }),
        .S(pc[11:8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[12] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[12]_i_1_n_0 ),
        .Q(pc[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[13] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[13]_i_1_n_0 ),
        .Q(pc[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[14] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[14]_i_1_n_0 ),
        .Q(pc[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[15] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[15]_i_2_n_0 ),
        .Q(pc[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \pc_reg[15]_i_7 
       (.CI(pc_reg[3]),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\pc_reg[15]_i_7_n_4 ,\pc_reg[15]_i_7_n_5 ,\pc_reg[15]_i_7_n_6 ,\pc_reg[15]_i_7_n_7 }),
        .S(pc[15:12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[1] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\pc[1]_i_1_n_0 ),
        .Q(pc[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[2] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[2]_i_1_n_0 ),
        .Q(pc[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[3] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[3]_i_1_n_0 ),
        .Q(pc[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \pc_reg[3]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\pc_reg[3]_i_2_n_0 ,\pc_reg[3]_i_2_n_1 ,\pc_reg[3]_i_2_n_2 ,\pc_reg[3]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,pc[1],\<const0>__0__0 }),
        .O({\pc_reg[3]_i_2_n_4 ,\pc_reg[3]_i_2_n_5 ,\pc_reg[3]_i_2_n_6 ,\pc_reg[3]_i_2_n_7 }),
        .S({pc[3:2],\pc[3]_i_5_n_0 ,pc[0]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[4] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[4]_i_1_n_0 ),
        .Q(pc[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[5] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[5]_i_1_n_0 ),
        .Q(pc[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[6] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[6]_i_1_n_0 ),
        .Q(pc[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[7] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[7]_i_1_n_0 ),
        .Q(pc[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \pc_reg[7]_i_2 
       (.CI(\pc_reg[3]_i_2_n_0 ),
        .CO({\pc_reg[7]_i_2_n_0 ,\pc_reg[7]_i_2_n_1 ,\pc_reg[7]_i_2_n_2 ,\pc_reg[7]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\pc_reg[7]_i_2_n_4 ,\pc_reg[7]_i_2_n_5 ,\pc_reg[7]_i_2_n_6 ,\pc_reg[7]_i_2_n_7 }),
        .S(pc[7:4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[8] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[8]_i_1_n_0 ),
        .Q(pc[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \pc_reg[9] 
       (.C(clk),
        .CE(\pc[15]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\pc[9]_i_1_n_0 ),
        .Q(pc[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4544454445445555)) 
    \r[10][0]_i_1 
       (.I0(halt),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r[10][0]_i_4_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(\r[8][0]_i_5_n_0 ),
        .I5(\r[10][0]_i_5_n_0 ),
        .O(\r[10][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF909)) 
    \r[10][0]_i_10 
       (.I0(bw),
        .I1(\r_reg[10] [1]),
        .I2(\r[10][0]_i_3_n_0 ),
        .I3(\dout[1]_INST_0_i_1_n_0 ),
        .O(r));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF606)) 
    \r[10][0]_i_11 
       (.I0(bw),
        .I1(\r_reg[10] [0]),
        .I2(\r[10][0]_i_3_n_0 ),
        .I3(\dout[0]_INST_0_i_1_n_0 ),
        .O(\r[10][0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00400000)) 
    \r[10][0]_i_3 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\addr[3]_INST_0_i_9_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\r_code[0]_i_1_n_0 ),
        .I4(\r_code[1]_i_1_n_0 ),
        .O(\r[10][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFDFFFFFFFDFDFDF)) 
    \r[10][0]_i_4 
       (.I0(\r_code[1]_i_1_n_0 ),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(din[2]),
        .I4(p_2_in88_in),
        .I5(r_code[2]),
        .O(\r[10][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCAFFFAF)) 
    \r[10][0]_i_5 
       (.I0(r_code[10]),
        .I1(din[10]),
        .I2(r_code[9]),
        .I3(p_2_in88_in),
        .I4(din[9]),
        .O(\r[10][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[10][0]_i_6 
       (.I0(bw),
        .I1(\r[10][0]_i_3_n_0 ),
        .O(\r[10][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[10][0]_i_7 
       (.I0(bw),
        .I1(\r[10][0]_i_3_n_0 ),
        .O(\r[10][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][0]_i_8 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [3]),
        .O(\r[10][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][0]_i_9 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [2]),
        .O(\r[10][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][12]_i_2 
       (.I0(\dout[15]_INST_0_i_3_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [15]),
        .O(\r[10][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [14]),
        .O(\r[10][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [13]),
        .O(\r[10][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [12]),
        .O(\r[10][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [7]),
        .O(\r[10][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [6]),
        .O(\r[10][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [5]),
        .O(\r[10][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [4]),
        .O(\r[10][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [11]),
        .O(\r[10][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [10]),
        .O(\r[10][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [9]),
        .O(\r[10][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[10][8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\r[10][0]_i_3_n_0 ),
        .I2(\r_reg[10] [8]),
        .O(\r[10][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4544454445445555)) 
    \r[11][0]_i_1 
       (.I0(halt),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r[11][0]_i_4_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(\r[9][0]_i_5_n_0 ),
        .I5(\r[10][0]_i_5_n_0 ),
        .O(\r[11][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF606)) 
    \r[11][0]_i_10 
       (.I0(bw),
        .I1(\r_reg[11] [0]),
        .I2(\r[11][0]_i_3_n_0 ),
        .I3(\dout[0]_INST_0_i_1_n_0 ),
        .O(\r[11][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h40000000)) 
    \r[11][0]_i_3 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\addr[3]_INST_0_i_9_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\r_code[0]_i_1_n_0 ),
        .I4(\r_code[1]_i_1_n_0 ),
        .O(\r[11][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF7FFFFFFF7F7F7F)) 
    \r[11][0]_i_4 
       (.I0(\r_code[1]_i_1_n_0 ),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(din[2]),
        .I4(p_2_in88_in),
        .I5(r_code[2]),
        .O(\r[11][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[11][0]_i_5 
       (.I0(bw),
        .I1(\r[11][0]_i_3_n_0 ),
        .O(\r[11][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[11][0]_i_6 
       (.I0(bw),
        .I1(\r[11][0]_i_3_n_0 ),
        .O(\r[11][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][0]_i_7 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [3]),
        .O(\r[11][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][0]_i_8 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [2]),
        .O(\r[11][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF909)) 
    \r[11][0]_i_9 
       (.I0(bw),
        .I1(\r_reg[11] [1]),
        .I2(\r[11][0]_i_3_n_0 ),
        .I3(\dout[1]_INST_0_i_1_n_0 ),
        .O(\r[11][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][12]_i_2 
       (.I0(\dout[15]_INST_0_i_3_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [15]),
        .O(\r[11][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [14]),
        .O(\r[11][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [13]),
        .O(\r[11][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [12]),
        .O(\r[11][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [7]),
        .O(\r[11][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [6]),
        .O(\r[11][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [5]),
        .O(\r[11][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [4]),
        .O(\r[11][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [11]),
        .O(\r[11][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [10]),
        .O(\r[11][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [9]),
        .O(\r[11][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[11][8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\r[11][0]_i_3_n_0 ),
        .I2(\r_reg[11] [8]),
        .O(\r[11][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4544555545444544)) 
    \r[12][0]_i_1 
       (.I0(halt),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r[12][0]_i_4_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(\r[4][0]_i_6_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\r[12][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF606)) 
    \r[12][0]_i_10 
       (.I0(bw),
        .I1(\r_reg[12] [0]),
        .I2(\r[12][0]_i_3_n_0 ),
        .I3(\dout[0]_INST_0_i_1_n_0 ),
        .O(\r[12][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000004)) 
    \r[12][0]_i_3 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\r_code[3]_i_1_n_0 ),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_9_n_0 ),
        .I4(\r_code[1]_i_1_n_0 ),
        .O(\r[12][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFABFBFFFFFFFF)) 
    \r[12][0]_i_4 
       (.I0(\r_code[1]_i_1_n_0 ),
        .I1(r_code[2]),
        .I2(p_2_in88_in),
        .I3(din[2]),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\r[12][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[12][0]_i_5 
       (.I0(bw),
        .I1(\r[12][0]_i_3_n_0 ),
        .O(\r[12][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[12][0]_i_6 
       (.I0(bw),
        .I1(\r[12][0]_i_3_n_0 ),
        .O(\r[12][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][0]_i_7 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [3]),
        .O(\r[12][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][0]_i_8 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [2]),
        .O(\r[12][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF909)) 
    \r[12][0]_i_9 
       (.I0(bw),
        .I1(\r_reg[12] [1]),
        .I2(\r[12][0]_i_3_n_0 ),
        .I3(\dout[1]_INST_0_i_1_n_0 ),
        .O(\r[12][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][12]_i_2 
       (.I0(\dout[15]_INST_0_i_3_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [15]),
        .O(\r[12][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [14]),
        .O(\r[12][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [13]),
        .O(\r[12][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [12]),
        .O(\r[12][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [7]),
        .O(\r[12][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [6]),
        .O(\r[12][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [5]),
        .O(\r[12][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [4]),
        .O(\r[12][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [11]),
        .O(\r[12][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [10]),
        .O(\r[12][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [9]),
        .O(\r[12][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[12][8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\r[12][0]_i_3_n_0 ),
        .I2(\r_reg[12] [8]),
        .O(\r[12][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4544555545444544)) 
    \r[13][0]_i_1 
       (.I0(halt),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r[13][0]_i_4_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(\r[5][0]_i_5_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\r[13][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF606)) 
    \r[13][0]_i_10 
       (.I0(bw),
        .I1(\r_reg[13] [0]),
        .I2(\r[13][0]_i_3_n_0 ),
        .I3(\dout[0]_INST_0_i_1_n_0 ),
        .O(\r[13][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \r[13][0]_i_3 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\r_code[3]_i_1_n_0 ),
        .I2(\addr[3]_INST_0_i_9_n_0 ),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(\r_code[0]_i_1_n_0 ),
        .O(\r[13][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDDFFFDFFFFFFFFF)) 
    \r[13][0]_i_4 
       (.I0(\r_code[0]_i_1_n_0 ),
        .I1(\r_code[1]_i_1_n_0 ),
        .I2(r_code[2]),
        .I3(p_2_in88_in),
        .I4(din[2]),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\r[13][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[13][0]_i_5 
       (.I0(bw),
        .I1(\r[13][0]_i_3_n_0 ),
        .O(\r[13][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[13][0]_i_6 
       (.I0(bw),
        .I1(\r[13][0]_i_3_n_0 ),
        .O(\r[13][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][0]_i_7 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [3]),
        .O(\r[13][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][0]_i_8 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [2]),
        .O(\r[13][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF909)) 
    \r[13][0]_i_9 
       (.I0(bw),
        .I1(\r_reg[13] [1]),
        .I2(\r[13][0]_i_3_n_0 ),
        .I3(\dout[1]_INST_0_i_1_n_0 ),
        .O(\r[13][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][12]_i_2 
       (.I0(\dout[15]_INST_0_i_3_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [15]),
        .O(\r[13][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [14]),
        .O(\r[13][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [13]),
        .O(\r[13][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [12]),
        .O(\r[13][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [7]),
        .O(\r[13][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [6]),
        .O(\r[13][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [5]),
        .O(\r[13][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [4]),
        .O(\r[13][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [11]),
        .O(\r[13][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [10]),
        .O(\r[13][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [9]),
        .O(\r[13][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[13][8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\r[13][0]_i_3_n_0 ),
        .I2(\r_reg[13] [8]),
        .O(\r[13][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4544555545444544)) 
    \r[14][0]_i_1 
       (.I0(halt),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r[14][0]_i_4_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(\r[6][0]_i_5_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\r[14][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF606)) 
    \r[14][0]_i_10 
       (.I0(bw),
        .I1(\r_reg[14] [0]),
        .I2(\r[14][0]_i_3_n_0 ),
        .I3(\dout[0]_INST_0_i_1_n_0 ),
        .O(\r[14][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \r[14][0]_i_3 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\r_code[3]_i_1_n_0 ),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(\addr[3]_INST_0_i_9_n_0 ),
        .O(\r[14][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF1DFFFFFFFFFF)) 
    \r[14][0]_i_4 
       (.I0(r_code[2]),
        .I1(p_2_in88_in),
        .I2(din[2]),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(\r_code[0]_i_1_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\r[14][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[14][0]_i_5 
       (.I0(bw),
        .I1(\r[14][0]_i_3_n_0 ),
        .O(\r[14][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[14][0]_i_6 
       (.I0(bw),
        .I1(\r[14][0]_i_3_n_0 ),
        .O(\r[14][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][0]_i_7 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [3]),
        .O(\r[14][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][0]_i_8 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [2]),
        .O(\r[14][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF909)) 
    \r[14][0]_i_9 
       (.I0(bw),
        .I1(\r_reg[14] [1]),
        .I2(\r[14][0]_i_3_n_0 ),
        .I3(\dout[1]_INST_0_i_1_n_0 ),
        .O(\r[14][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][12]_i_2 
       (.I0(\dout[15]_INST_0_i_3_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [15]),
        .O(\r[14][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [14]),
        .O(\r[14][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [13]),
        .O(\r[14][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [12]),
        .O(\r[14][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [7]),
        .O(\r[14][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [6]),
        .O(\r[14][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [5]),
        .O(\r[14][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [4]),
        .O(\r[14][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [11]),
        .O(\r[14][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [10]),
        .O(\r[14][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [9]),
        .O(\r[14][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[14][8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\r[14][0]_i_3_n_0 ),
        .I2(\r_reg[14] [8]),
        .O(\r[14][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4544555545444544)) 
    \r[15][0]_i_1 
       (.I0(halt),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r[15][0]_i_4_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(\r[7][0]_i_5_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\r[15][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF606)) 
    \r[15][0]_i_10 
       (.I0(bw),
        .I1(\r_reg[15] [0]),
        .I2(\r[15][0]_i_3_n_0 ),
        .I3(\dout[0]_INST_0_i_1_n_0 ),
        .O(\r[15][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00400000)) 
    \r[15][0]_i_3 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\r_code[3]_i_1_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_9_n_0 ),
        .I4(\r_code[0]_i_1_n_0 ),
        .O(\r[15][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h57F7FFFFFFFFFFFF)) 
    \r[15][0]_i_4 
       (.I0(\r_code[0]_i_1_n_0 ),
        .I1(r_code[2]),
        .I2(p_2_in88_in),
        .I3(din[2]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\r[15][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[15][0]_i_5 
       (.I0(bw),
        .I1(\r[15][0]_i_3_n_0 ),
        .O(\r[15][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[15][0]_i_6 
       (.I0(bw),
        .I1(\r[15][0]_i_3_n_0 ),
        .O(\r[15][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][0]_i_7 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [3]),
        .O(\r[15][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][0]_i_8 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [2]),
        .O(\r[15][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF909)) 
    \r[15][0]_i_9 
       (.I0(bw),
        .I1(\r_reg[15] [1]),
        .I2(\r[15][0]_i_3_n_0 ),
        .I3(\dout[1]_INST_0_i_1_n_0 ),
        .O(\r[15][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][12]_i_2 
       (.I0(\dout[15]_INST_0_i_3_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [15]),
        .O(\r[15][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [14]),
        .O(\r[15][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [13]),
        .O(\r[15][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [12]),
        .O(\r[15][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [7]),
        .O(\r[15][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0_repN ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [6]),
        .O(\r[15][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [5]),
        .O(\r[15][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [4]),
        .O(\r[15][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [11]),
        .O(\r[15][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [10]),
        .O(\r[15][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [9]),
        .O(\r[15][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[15][8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\r[15][0]_i_3_n_0 ),
        .I2(\r_reg[15] [8]),
        .O(\r[15][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4544454445445555)) 
    \r[4][0]_i_1 
       (.I0(halt),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r[4][0]_i_4_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(\r[4][0]_i_6_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\r[4][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][0]_i_10 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [2]),
        .O(\r[4][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF909)) 
    \r[4][0]_i_11 
       (.I0(bw),
        .I1(\r_reg[4] [1]),
        .I2(\r[4][0]_i_3_n_0 ),
        .I3(\dout[1]_INST_0_i_1_n_0 ),
        .O(\r[4][0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF606)) 
    \r[4][0]_i_12 
       (.I0(bw),
        .I1(\r_reg[4] [0]),
        .I2(\r[4][0]_i_3_n_0 ),
        .I3(\dout[0]_INST_0_i_1_n_0 ),
        .O(\r[4][0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \r[4][0]_i_3 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\addr[3]_INST_0_i_9_n_0 ),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(\r_code[3]_i_1_n_0 ),
        .O(\r[4][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEFFFEF)) 
    \r[4][0]_i_4 
       (.I0(\r_code[3]_i_1_n_0 ),
        .I1(\r_code[1]_i_1_n_0 ),
        .I2(r_code[2]),
        .I3(p_2_in88_in),
        .I4(din[2]),
        .I5(\r_code[0]_i_1_n_0 ),
        .O(\r[4][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h2A)) 
    \r[4][0]_i_5 
       (.I0(\pc[15]_i_9_n_0 ),
        .I1(\r_code[1]_i_1_n_0 ),
        .I2(\addr[15]_INST_0_i_11_n_0 ),
        .O(\r[4][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFBFF)) 
    \r[4][0]_i_6 
       (.I0(soc[2]),
        .I1(\r_code[10]_i_1_n_0 ),
        .I2(soc[1]),
        .I3(\sp[0]_i_4_n_0 ),
        .O(\r[4][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[4][0]_i_7 
       (.I0(bw),
        .I1(\r[4][0]_i_3_n_0 ),
        .O(\r[4][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[4][0]_i_8 
       (.I0(bw),
        .I1(\r[4][0]_i_3_n_0 ),
        .O(\r[4][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][0]_i_9 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [3]),
        .O(\r[4][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][12]_i_2 
       (.I0(\dout[15]_INST_0_i_3_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [15]),
        .O(\r[4][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [14]),
        .O(\r[4][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [13]),
        .O(\r[4][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [12]),
        .O(\r[4][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [7]),
        .O(\r[4][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [6]),
        .O(\r[4][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [5]),
        .O(\r[4][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [4]),
        .O(\r[4][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [11]),
        .O(\r[4][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [10]),
        .O(\r[4][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [9]),
        .O(\r[4][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[4][8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\r[4][0]_i_3_n_0 ),
        .I2(\r_reg[4] [8]),
        .O(\r[4][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4544454445445555)) 
    \r[5][0]_i_1 
       (.I0(halt),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r[5][0]_i_4_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(\r[5][0]_i_5_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\r[5][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF909)) 
    \r[5][0]_i_10 
       (.I0(bw),
        .I1(\r_reg[5] [1]),
        .I2(\r[5][0]_i_3_n_0 ),
        .I3(\dout[1]_INST_0_i_1_n_0 ),
        .O(\r[5][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF606)) 
    \r[5][0]_i_11 
       (.I0(bw),
        .I1(\r_reg[5] [0]),
        .I2(\r[5][0]_i_3_n_0 ),
        .I3(\dout[0]_INST_0_i_1_n_0 ),
        .O(\r[5][0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000100)) 
    \r[5][0]_i_3 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\addr[3]_INST_0_i_9_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_code[0]_i_1_n_0 ),
        .I4(\r_code[3]_i_1_n_0 ),
        .O(\r[5][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBFBFBFFFFFFFBFF)) 
    \r[5][0]_i_4 
       (.I0(\r_code[3]_i_1_n_0 ),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(r_code[2]),
        .I4(p_2_in88_in),
        .I5(din[2]),
        .O(\r[5][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hDFFF)) 
    \r[5][0]_i_5 
       (.I0(soc[1]),
        .I1(soc[2]),
        .I2(\r_code[10]_i_1_n_0 ),
        .I3(\sp[0]_i_4_n_0 ),
        .O(\r[5][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[5][0]_i_6 
       (.I0(bw),
        .I1(\r[5][0]_i_3_n_0 ),
        .O(\r[5][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[5][0]_i_7 
       (.I0(bw),
        .I1(\r[5][0]_i_3_n_0 ),
        .O(\r[5][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][0]_i_8 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [3]),
        .O(\r[5][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][0]_i_9 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [2]),
        .O(\r[5][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][12]_i_2 
       (.I0(\dout[15]_INST_0_i_3_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [15]),
        .O(\r[5][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [14]),
        .O(\r[5][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [13]),
        .O(\r[5][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [12]),
        .O(\r[5][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [7]),
        .O(\r[5][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [6]),
        .O(\r[5][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [5]),
        .O(\r[5][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [4]),
        .O(\r[5][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [11]),
        .O(\r[5][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [10]),
        .O(\r[5][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [9]),
        .O(\r[5][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[5][8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\r[5][0]_i_3_n_0 ),
        .I2(\r_reg[5] [8]),
        .O(\r[5][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4544454445445555)) 
    \r[6][0]_i_1 
       (.I0(halt),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r[6][0]_i_4_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(\r[6][0]_i_5_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\r[6][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF909)) 
    \r[6][0]_i_10 
       (.I0(bw),
        .I1(\r_reg[6] [1]),
        .I2(\r[6][0]_i_3_n_0 ),
        .I3(\dout[1]_INST_0_i_1_n_0 ),
        .O(\r[6][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF606)) 
    \r[6][0]_i_11 
       (.I0(bw),
        .I1(\r_reg[6] [0]),
        .I2(\r[6][0]_i_3_n_0 ),
        .I3(\dout[0]_INST_0_i_1_n_0 ),
        .O(\r[6][0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \r[6][0]_i_3 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\addr[3]_INST_0_i_9_n_0 ),
        .I4(\r_code[3]_i_1_n_0 ),
        .O(\r[6][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFABFBFFFF)) 
    \r[6][0]_i_4 
       (.I0(\r_code[3]_i_1_n_0 ),
        .I1(r_code[2]),
        .I2(p_2_in88_in),
        .I3(din[2]),
        .I4(\r_code[1]_i_1_n_0 ),
        .I5(\r_code[0]_i_1_n_0 ),
        .O(\r[6][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF7F)) 
    \r[6][0]_i_5 
       (.I0(\sp[0]_i_4_n_0 ),
        .I1(\r_code[10]_i_1_n_0 ),
        .I2(soc[2]),
        .I3(soc[1]),
        .O(\r[6][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[6][0]_i_6 
       (.I0(bw),
        .I1(\r[6][0]_i_3_n_0 ),
        .O(\r[6][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[6][0]_i_7 
       (.I0(bw),
        .I1(\r[6][0]_i_3_n_0 ),
        .O(\r[6][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][0]_i_8 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [3]),
        .O(\r[6][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][0]_i_9 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [2]),
        .O(\r[6][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][12]_i_2 
       (.I0(\dout[15]_INST_0_i_3_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [15]),
        .O(\r[6][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [14]),
        .O(\r[6][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [13]),
        .O(\r[6][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [12]),
        .O(\r[6][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [7]),
        .O(\r[6][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [6]),
        .O(\r[6][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [5]),
        .O(\r[6][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [4]),
        .O(\r[6][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [11]),
        .O(\r[6][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [10]),
        .O(\r[6][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [9]),
        .O(\r[6][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[6][8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\r[6][0]_i_3_n_0 ),
        .I2(\r_reg[6] [8]),
        .O(\r[6][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4544454445445555)) 
    \r[7][0]_i_1 
       (.I0(halt),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r[7][0]_i_4_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(\r[7][0]_i_5_n_0 ),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(\r[7][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF909)) 
    \r[7][0]_i_10 
       (.I0(bw),
        .I1(\r_reg[7] [1]),
        .I2(\r[7][0]_i_3_n_0 ),
        .I3(\dout[1]_INST_0_i_1_n_0 ),
        .O(\r[7][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF606)) 
    \r[7][0]_i_11 
       (.I0(bw),
        .I1(\r_reg[7] [0]),
        .I2(\r[7][0]_i_3_n_0 ),
        .I3(\dout[0]_INST_0_i_1_n_0 ),
        .O(\r[7][0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000400)) 
    \r[7][0]_i_3 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\r_code[1]_i_1_n_0 ),
        .I2(\addr[3]_INST_0_i_9_n_0 ),
        .I3(\r_code[0]_i_1_n_0 ),
        .I4(\r_code[3]_i_1_n_0 ),
        .O(\r[7][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBFFFBFFFFFFFFF)) 
    \r[7][0]_i_4 
       (.I0(\r_code[3]_i_1_n_0 ),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(r_code[2]),
        .I3(p_2_in88_in),
        .I4(din[2]),
        .I5(\r_code[1]_i_1_n_0 ),
        .O(\r[7][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \r[7][0]_i_5 
       (.I0(\sp[0]_i_4_n_0 ),
        .I1(soc[2]),
        .I2(soc[1]),
        .I3(\r_code[10]_i_1_n_0 ),
        .O(\r[7][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[7][0]_i_6 
       (.I0(bw),
        .I1(\r[7][0]_i_3_n_0 ),
        .O(\r[7][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[7][0]_i_7 
       (.I0(bw),
        .I1(\r[7][0]_i_3_n_0 ),
        .O(\r[7][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][0]_i_8 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [3]),
        .O(\r[7][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][0]_i_9 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [2]),
        .O(\r[7][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][12]_i_2 
       (.I0(\dout[15]_INST_0_i_3_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [15]),
        .O(\r[7][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [14]),
        .O(\r[7][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [13]),
        .O(\r[7][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [12]),
        .O(\r[7][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [7]),
        .O(\r[7][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [6]),
        .O(\r[7][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [5]),
        .O(\r[7][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [4]),
        .O(\r[7][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [11]),
        .O(\r[7][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [10]),
        .O(\r[7][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [9]),
        .O(\r[7][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[7][8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\r[7][0]_i_3_n_0 ),
        .I2(\r_reg[7] [8]),
        .O(\r[7][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4544454445445555)) 
    \r[8][0]_i_1 
       (.I0(halt),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r[8][0]_i_4_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(\r[8][0]_i_5_n_0 ),
        .I5(\r[8][0]_i_6_n_0 ),
        .O(\r[8][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][0]_i_10 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [2]),
        .O(\r[8][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF909)) 
    \r[8][0]_i_11 
       (.I0(bw),
        .I1(\r_reg[8] [1]),
        .I2(\r[8][0]_i_3_n_0 ),
        .I3(\dout[1]_INST_0_i_1_n_0 ),
        .O(\r[8][0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF606)) 
    \r[8][0]_i_12 
       (.I0(bw),
        .I1(\r_reg[8] [0]),
        .I2(\r[8][0]_i_3_n_0 ),
        .I3(\dout[0]_INST_0_i_1_n_0 ),
        .O(\r[8][0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \r[8][0]_i_3 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\addr[3]_INST_0_i_9_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(\r_code[0]_i_1_n_0 ),
        .I4(\r_code[1]_i_1_n_0 ),
        .O(\r[8][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFEFFFFFFFEFEFEF)) 
    \r[8][0]_i_4 
       (.I0(\r_code[1]_i_1_n_0 ),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\r_code[3]_i_1_n_0 ),
        .I3(din[2]),
        .I4(p_2_in88_in),
        .I5(r_code[2]),
        .O(\r[8][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \r[8][0]_i_5 
       (.I0(\sp[0]_i_4_n_0 ),
        .I1(soc[1]),
        .I2(\r_code[11]_i_1_n_0 ),
        .O(\r[8][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFACCFA)) 
    \r[8][0]_i_6 
       (.I0(r_code[10]),
        .I1(din[10]),
        .I2(r_code[9]),
        .I3(p_2_in88_in),
        .I4(din[9]),
        .O(\r[8][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[8][0]_i_7 
       (.I0(bw),
        .I1(\r[8][0]_i_3_n_0 ),
        .O(\r[8][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[8][0]_i_8 
       (.I0(bw),
        .I1(\r[8][0]_i_3_n_0 ),
        .O(\r[8][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][0]_i_9 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [3]),
        .O(\r[8][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][12]_i_2 
       (.I0(\dout[15]_INST_0_i_3_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [15]),
        .O(\r[8][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [14]),
        .O(\r[8][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [13]),
        .O(\r[8][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [12]),
        .O(\r[8][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [7]),
        .O(\r[8][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [6]),
        .O(\r[8][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [5]),
        .O(\r[8][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [4]),
        .O(\r[8][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [11]),
        .O(\r[8][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [10]),
        .O(\r[8][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [9]),
        .O(\r[8][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[8][8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\r[8][0]_i_3_n_0 ),
        .I2(\r_reg[8] [8]),
        .O(\r[8][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4544454445445555)) 
    \r[9][0]_i_1 
       (.I0(halt),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r[9][0]_i_4_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(\r[9][0]_i_5_n_0 ),
        .I5(\r[8][0]_i_6_n_0 ),
        .O(\r[9][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF909)) 
    \r[9][0]_i_10 
       (.I0(bw),
        .I1(\r_reg[9] [1]),
        .I2(\r[9][0]_i_3_n_0 ),
        .I3(\dout[1]_INST_0_i_1_n_0 ),
        .O(\r[9][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF606)) 
    \r[9][0]_i_11 
       (.I0(bw),
        .I1(\r_reg[9] [0]),
        .I2(\r[9][0]_i_3_n_0 ),
        .I3(\dout[0]_INST_0_i_1_n_0 ),
        .O(\r[9][0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00400000)) 
    \r[9][0]_i_3 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\r_code[3]_i_1_n_0 ),
        .I2(\addr[3]_INST_0_i_9_n_0 ),
        .I3(\r_code[1]_i_1_n_0 ),
        .I4(\r_code[0]_i_1_n_0 ),
        .O(\r[9][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFDDDFDFFFFFFFF)) 
    \r[9][0]_i_4 
       (.I0(\r_code[0]_i_1_n_0 ),
        .I1(\r_code[1]_i_1_n_0 ),
        .I2(r_code[2]),
        .I3(p_2_in88_in),
        .I4(din[2]),
        .I5(\r_code[3]_i_1_n_0 ),
        .O(\r[9][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \r[9][0]_i_5 
       (.I0(\sp[0]_i_4_n_0 ),
        .I1(soc[1]),
        .I2(\r_code[11]_i_1_n_0 ),
        .O(\r[9][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[9][0]_i_6 
       (.I0(bw),
        .I1(\r[9][0]_i_3_n_0 ),
        .O(\r[9][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r[9][0]_i_7 
       (.I0(bw),
        .I1(\r[9][0]_i_3_n_0 ),
        .O(\r[9][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][0]_i_8 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [3]),
        .O(\r[9][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][0]_i_9 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [2]),
        .O(\r[9][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][12]_i_2 
       (.I0(\dout[15]_INST_0_i_3_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [15]),
        .O(\r[9][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [14]),
        .O(\r[9][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [13]),
        .O(\r[9][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [12]),
        .O(\r[9][12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [7]),
        .O(\r[9][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [6]),
        .O(\r[9][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [5]),
        .O(\r[9][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [4]),
        .O(\r[9][4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [11]),
        .O(\r[9][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [10]),
        .O(\r[9][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [9]),
        .O(\r[9][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[9][8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\r[9][0]_i_3_n_0 ),
        .I2(\r_reg[9] [8]),
        .O(\r[9][8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    r_a0_reg
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(lbe_INST_0_i_3_n_0),
        .Q(r_a0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[0]_i_1 
       (.I0(din[0]),
        .I1(p_2_in88_in),
        .I2(r_code[0]),
        .O(\r_code[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[10]_i_1 
       (.I0(din[10]),
        .I1(p_2_in88_in),
        .I2(r_code[10]),
        .O(\r_code[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[11]_i_1 
       (.I0(din[11]),
        .I1(p_2_in88_in),
        .I2(r_code[11]),
        .O(\r_code[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[12]_i_1 
       (.I0(din[12]),
        .I1(p_2_in88_in),
        .I2(r_code[12]),
        .O(doc[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[13]_i_1 
       (.I0(din[13]),
        .I1(p_2_in88_in),
        .I2(r_code[13]),
        .O(doc[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[14]_i_1 
       (.I0(din[14]),
        .I1(p_2_in88_in),
        .I2(r_code[14]),
        .O(doc[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[15]_i_1 
       (.I0(din[15]),
        .I1(p_2_in88_in),
        .I2(r_code[15]),
        .O(doc[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[1]_i_1 
       (.I0(din[1]),
        .I1(p_2_in88_in),
        .I2(r_code[1]),
        .O(\r_code[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    \r_code[2]_i_1 
       (.I0(r_code[2]),
        .I1(p_2_in88_in),
        .I2(din[2]),
        .O(\r_code[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[3]_i_1 
       (.I0(din[3]),
        .I1(p_2_in88_in),
        .I2(r_code[3]),
        .O(\r_code[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[4]_i_1 
       (.I0(din[4]),
        .I1(p_2_in88_in),
        .I2(r_code[4]),
        .O(as[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[5]_i_1 
       (.I0(din[5]),
        .I1(p_2_in88_in),
        .I2(r_code[5]),
        .O(as[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[7]_i_1 
       (.I0(din[7]),
        .I1(p_2_in88_in),
        .I2(r_code[7]),
        .O(soc[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[8]_i_1 
       (.I0(din[8]),
        .I1(p_2_in88_in),
        .I2(r_code[8]),
        .O(soc[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_code[9]_i_1 
       (.I0(din[9]),
        .I1(p_2_in88_in),
        .I2(r_code[9]),
        .O(soc[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[0] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_code[0]_i_1_n_0 ),
        .Q(r_code[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[10] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_code[10]_i_1_n_0 ),
        .Q(r_code[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[11] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_code[11]_i_1_n_0 ),
        .Q(r_code[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[12] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(doc[0]),
        .Q(r_code[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[13] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(doc[1]),
        .Q(r_code[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[14] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(doc[2]),
        .Q(r_code[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[15] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(doc[3]),
        .Q(r_code[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[1] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_code[1]_i_1_n_0 ),
        .Q(r_code[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[2] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_code[2]_i_1_n_0 ),
        .Q(r_code[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[3] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_code[3]_i_1_n_0 ),
        .Q(r_code[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[4] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(as[0]),
        .Q(r_code[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[5] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(as[1]),
        .Q(r_code[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[6] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(bw),
        .Q(r_code[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[7] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(soc[0]),
        .Q(r_code[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[8] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(soc[1]),
        .Q(r_code[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_code_reg[9] 
       (.C(clk),
        .CE(\FSM_sequential_state[4]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(soc[2]),
        .Q(r_code[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][0] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[10][0]_i_2_n_7 ),
        .Q(\r_reg[10] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[10][0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO(r_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r[10][0]_i_6_n_0 ,\r[10][0]_i_7_n_0 }),
        .O({\r_reg[10][0]_i_2_n_4 ,\r_reg[10][0]_i_2_n_5 ,\r_reg[10][0]_i_2_n_6 ,\r_reg[10][0]_i_2_n_7 }),
        .S({\r[10][0]_i_8_n_0 ,\r[10][0]_i_9_n_0 ,r,\r[10][0]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][10] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[10][8]_i_1_n_5 ),
        .Q(\r_reg[10] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][11] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[10][8]_i_1_n_4 ),
        .Q(\r_reg[10] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][12] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[10][12]_i_1_n_7 ),
        .Q(\r_reg[10] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[10][12]_i_1 
       (.CI(\r_reg[10][8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[10][12]_i_1_n_4 ,\r_reg[10][12]_i_1_n_5 ,\r_reg[10][12]_i_1_n_6 ,\r_reg[10][12]_i_1_n_7 }),
        .S({\r[10][12]_i_2_n_0 ,\r[10][12]_i_3_n_0 ,\r[10][12]_i_4_n_0 ,\r[10][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][13] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[10][12]_i_1_n_6 ),
        .Q(\r_reg[10] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][14] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[10][12]_i_1_n_5 ),
        .Q(\r_reg[10] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][15] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[10][12]_i_1_n_4 ),
        .Q(\r_reg[10] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][1] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[10][0]_i_2_n_6 ),
        .Q(\r_reg[10] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][2] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[10][0]_i_2_n_5 ),
        .Q(\r_reg[10] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][3] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[10][0]_i_2_n_4 ),
        .Q(\r_reg[10] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][4] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[10][4]_i_1_n_7 ),
        .Q(\r_reg[10] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[10][4]_i_1 
       (.CI(r_reg[3]),
        .CO({\r_reg[10][4]_i_1_n_0 ,\r_reg[10][4]_i_1_n_1 ,\r_reg[10][4]_i_1_n_2 ,\r_reg[10][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[10][4]_i_1_n_4 ,\r_reg[10][4]_i_1_n_5 ,\r_reg[10][4]_i_1_n_6 ,\r_reg[10][4]_i_1_n_7 }),
        .S({\r[10][4]_i_2_n_0 ,\r[10][4]_i_3_n_0 ,\r[10][4]_i_4_n_0 ,\r[10][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][5] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[10][4]_i_1_n_6 ),
        .Q(\r_reg[10] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][6] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[10][4]_i_1_n_5 ),
        .Q(\r_reg[10] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][7] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[10][4]_i_1_n_4 ),
        .Q(\r_reg[10] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][8] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[10][8]_i_1_n_7 ),
        .Q(\r_reg[10] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[10][8]_i_1 
       (.CI(\r_reg[10][4]_i_1_n_0 ),
        .CO({\r_reg[10][8]_i_1_n_0 ,\r_reg[10][8]_i_1_n_1 ,\r_reg[10][8]_i_1_n_2 ,\r_reg[10][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[10][8]_i_1_n_4 ,\r_reg[10][8]_i_1_n_5 ,\r_reg[10][8]_i_1_n_6 ,\r_reg[10][8]_i_1_n_7 }),
        .S({\r[10][8]_i_2_n_0 ,\r[10][8]_i_3_n_0 ,\r[10][8]_i_4_n_0 ,\r[10][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[10][9] 
       (.C(clk),
        .CE(\r[10][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[10][8]_i_1_n_6 ),
        .Q(\r_reg[10] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][0] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[11][0]_i_2_n_7 ),
        .Q(\r_reg[11] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[11][0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[11][0]_i_2_n_0 ,\r_reg[11][0]_i_2_n_1 ,\r_reg[11][0]_i_2_n_2 ,\r_reg[11][0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r[11][0]_i_5_n_0 ,\r[11][0]_i_6_n_0 }),
        .O({\r_reg[11][0]_i_2_n_4 ,\r_reg[11][0]_i_2_n_5 ,\r_reg[11][0]_i_2_n_6 ,\r_reg[11][0]_i_2_n_7 }),
        .S({\r[11][0]_i_7_n_0 ,\r[11][0]_i_8_n_0 ,\r[11][0]_i_9_n_0 ,\r[11][0]_i_10_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][10] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[11][8]_i_1_n_5 ),
        .Q(\r_reg[11] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][11] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[11][8]_i_1_n_4 ),
        .Q(\r_reg[11] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][12] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[11][12]_i_1_n_7 ),
        .Q(\r_reg[11] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[11][12]_i_1 
       (.CI(\r_reg[11][8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[11][12]_i_1_n_4 ,\r_reg[11][12]_i_1_n_5 ,\r_reg[11][12]_i_1_n_6 ,\r_reg[11][12]_i_1_n_7 }),
        .S({\r[11][12]_i_2_n_0 ,\r[11][12]_i_3_n_0 ,\r[11][12]_i_4_n_0 ,\r[11][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][13] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[11][12]_i_1_n_6 ),
        .Q(\r_reg[11] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][14] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[11][12]_i_1_n_5 ),
        .Q(\r_reg[11] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][15] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[11][12]_i_1_n_4 ),
        .Q(\r_reg[11] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][1] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[11][0]_i_2_n_6 ),
        .Q(\r_reg[11] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][2] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[11][0]_i_2_n_5 ),
        .Q(\r_reg[11] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][3] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[11][0]_i_2_n_4 ),
        .Q(\r_reg[11] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][4] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[11][4]_i_1_n_7 ),
        .Q(\r_reg[11] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[11][4]_i_1 
       (.CI(\r_reg[11][0]_i_2_n_0 ),
        .CO({\r_reg[11][4]_i_1_n_0 ,\r_reg[11][4]_i_1_n_1 ,\r_reg[11][4]_i_1_n_2 ,\r_reg[11][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[11][4]_i_1_n_4 ,\r_reg[11][4]_i_1_n_5 ,\r_reg[11][4]_i_1_n_6 ,\r_reg[11][4]_i_1_n_7 }),
        .S({\r[11][4]_i_2_n_0 ,\r[11][4]_i_3_n_0 ,\r[11][4]_i_4_n_0 ,\r[11][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][5] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[11][4]_i_1_n_6 ),
        .Q(\r_reg[11] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][6] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[11][4]_i_1_n_5 ),
        .Q(\r_reg[11] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][7] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[11][4]_i_1_n_4 ),
        .Q(\r_reg[11] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][8] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[11][8]_i_1_n_7 ),
        .Q(\r_reg[11] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[11][8]_i_1 
       (.CI(\r_reg[11][4]_i_1_n_0 ),
        .CO({\r_reg[11][8]_i_1_n_0 ,\r_reg[11][8]_i_1_n_1 ,\r_reg[11][8]_i_1_n_2 ,\r_reg[11][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[11][8]_i_1_n_4 ,\r_reg[11][8]_i_1_n_5 ,\r_reg[11][8]_i_1_n_6 ,\r_reg[11][8]_i_1_n_7 }),
        .S({\r[11][8]_i_2_n_0 ,\r[11][8]_i_3_n_0 ,\r[11][8]_i_4_n_0 ,\r[11][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[11][9] 
       (.C(clk),
        .CE(\r[11][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[11][8]_i_1_n_6 ),
        .Q(\r_reg[11] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][0] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[12][0]_i_2_n_7 ),
        .Q(\r_reg[12] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[12][0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[12][0]_i_2_n_0 ,\r_reg[12][0]_i_2_n_1 ,\r_reg[12][0]_i_2_n_2 ,\r_reg[12][0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r[12][0]_i_5_n_0 ,\r[12][0]_i_6_n_0 }),
        .O({\r_reg[12][0]_i_2_n_4 ,\r_reg[12][0]_i_2_n_5 ,\r_reg[12][0]_i_2_n_6 ,\r_reg[12][0]_i_2_n_7 }),
        .S({\r[12][0]_i_7_n_0 ,\r[12][0]_i_8_n_0 ,\r[12][0]_i_9_n_0 ,\r[12][0]_i_10_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][10] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[12][8]_i_1_n_5 ),
        .Q(\r_reg[12] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][11] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[12][8]_i_1_n_4 ),
        .Q(\r_reg[12] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][12] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[12][12]_i_1_n_7 ),
        .Q(\r_reg[12] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[12][12]_i_1 
       (.CI(\r_reg[12][8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[12][12]_i_1_n_4 ,\r_reg[12][12]_i_1_n_5 ,\r_reg[12][12]_i_1_n_6 ,\r_reg[12][12]_i_1_n_7 }),
        .S({\r[12][12]_i_2_n_0 ,\r[12][12]_i_3_n_0 ,\r[12][12]_i_4_n_0 ,\r[12][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][13] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[12][12]_i_1_n_6 ),
        .Q(\r_reg[12] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][14] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[12][12]_i_1_n_5 ),
        .Q(\r_reg[12] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][15] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[12][12]_i_1_n_4 ),
        .Q(\r_reg[12] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][1] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[12][0]_i_2_n_6 ),
        .Q(\r_reg[12] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][2] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[12][0]_i_2_n_5 ),
        .Q(\r_reg[12] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][3] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[12][0]_i_2_n_4 ),
        .Q(\r_reg[12] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][4] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[12][4]_i_1_n_7 ),
        .Q(\r_reg[12] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[12][4]_i_1 
       (.CI(\r_reg[12][0]_i_2_n_0 ),
        .CO({\r_reg[12][4]_i_1_n_0 ,\r_reg[12][4]_i_1_n_1 ,\r_reg[12][4]_i_1_n_2 ,\r_reg[12][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[12][4]_i_1_n_4 ,\r_reg[12][4]_i_1_n_5 ,\r_reg[12][4]_i_1_n_6 ,\r_reg[12][4]_i_1_n_7 }),
        .S({\r[12][4]_i_2_n_0 ,\r[12][4]_i_3_n_0 ,\r[12][4]_i_4_n_0 ,\r[12][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][5] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[12][4]_i_1_n_6 ),
        .Q(\r_reg[12] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][6] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[12][4]_i_1_n_5 ),
        .Q(\r_reg[12] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][7] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[12][4]_i_1_n_4 ),
        .Q(\r_reg[12] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][8] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[12][8]_i_1_n_7 ),
        .Q(\r_reg[12] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[12][8]_i_1 
       (.CI(\r_reg[12][4]_i_1_n_0 ),
        .CO({\r_reg[12][8]_i_1_n_0 ,\r_reg[12][8]_i_1_n_1 ,\r_reg[12][8]_i_1_n_2 ,\r_reg[12][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[12][8]_i_1_n_4 ,\r_reg[12][8]_i_1_n_5 ,\r_reg[12][8]_i_1_n_6 ,\r_reg[12][8]_i_1_n_7 }),
        .S({\r[12][8]_i_2_n_0 ,\r[12][8]_i_3_n_0 ,\r[12][8]_i_4_n_0 ,\r[12][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[12][9] 
       (.C(clk),
        .CE(\r[12][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[12][8]_i_1_n_6 ),
        .Q(\r_reg[12] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][0] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[13][0]_i_2_n_7 ),
        .Q(\r_reg[13] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[13][0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[13][0]_i_2_n_0 ,\r_reg[13][0]_i_2_n_1 ,\r_reg[13][0]_i_2_n_2 ,\r_reg[13][0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r[13][0]_i_5_n_0 ,\r[13][0]_i_6_n_0 }),
        .O({\r_reg[13][0]_i_2_n_4 ,\r_reg[13][0]_i_2_n_5 ,\r_reg[13][0]_i_2_n_6 ,\r_reg[13][0]_i_2_n_7 }),
        .S({\r[13][0]_i_7_n_0 ,\r[13][0]_i_8_n_0 ,\r[13][0]_i_9_n_0 ,\r[13][0]_i_10_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][10] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[13][8]_i_1_n_5 ),
        .Q(\r_reg[13] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][11] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[13][8]_i_1_n_4 ),
        .Q(\r_reg[13] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][12] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[13][12]_i_1_n_7 ),
        .Q(\r_reg[13] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[13][12]_i_1 
       (.CI(\r_reg[13][8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[13][12]_i_1_n_4 ,\r_reg[13][12]_i_1_n_5 ,\r_reg[13][12]_i_1_n_6 ,\r_reg[13][12]_i_1_n_7 }),
        .S({\r[13][12]_i_2_n_0 ,\r[13][12]_i_3_n_0 ,\r[13][12]_i_4_n_0 ,\r[13][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][13] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[13][12]_i_1_n_6 ),
        .Q(\r_reg[13] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][14] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[13][12]_i_1_n_5 ),
        .Q(\r_reg[13] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][15] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[13][12]_i_1_n_4 ),
        .Q(\r_reg[13] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][1] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[13][0]_i_2_n_6 ),
        .Q(\r_reg[13] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][2] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[13][0]_i_2_n_5 ),
        .Q(\r_reg[13] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][3] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[13][0]_i_2_n_4 ),
        .Q(\r_reg[13] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][4] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[13][4]_i_1_n_7 ),
        .Q(\r_reg[13] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[13][4]_i_1 
       (.CI(\r_reg[13][0]_i_2_n_0 ),
        .CO({\r_reg[13][4]_i_1_n_0 ,\r_reg[13][4]_i_1_n_1 ,\r_reg[13][4]_i_1_n_2 ,\r_reg[13][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[13][4]_i_1_n_4 ,\r_reg[13][4]_i_1_n_5 ,\r_reg[13][4]_i_1_n_6 ,\r_reg[13][4]_i_1_n_7 }),
        .S({\r[13][4]_i_2_n_0 ,\r[13][4]_i_3_n_0 ,\r[13][4]_i_4_n_0 ,\r[13][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][5] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[13][4]_i_1_n_6 ),
        .Q(\r_reg[13] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][6] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[13][4]_i_1_n_5 ),
        .Q(\r_reg[13] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][7] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[13][4]_i_1_n_4 ),
        .Q(\r_reg[13] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][8] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[13][8]_i_1_n_7 ),
        .Q(\r_reg[13] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[13][8]_i_1 
       (.CI(\r_reg[13][4]_i_1_n_0 ),
        .CO({\r_reg[13][8]_i_1_n_0 ,\r_reg[13][8]_i_1_n_1 ,\r_reg[13][8]_i_1_n_2 ,\r_reg[13][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[13][8]_i_1_n_4 ,\r_reg[13][8]_i_1_n_5 ,\r_reg[13][8]_i_1_n_6 ,\r_reg[13][8]_i_1_n_7 }),
        .S({\r[13][8]_i_2_n_0 ,\r[13][8]_i_3_n_0 ,\r[13][8]_i_4_n_0 ,\r[13][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[13][9] 
       (.C(clk),
        .CE(\r[13][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[13][8]_i_1_n_6 ),
        .Q(\r_reg[13] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][0] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[14][0]_i_2_n_7 ),
        .Q(\r_reg[14] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[14][0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[14][0]_i_2_n_0 ,\r_reg[14][0]_i_2_n_1 ,\r_reg[14][0]_i_2_n_2 ,\r_reg[14][0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r[14][0]_i_5_n_0 ,\r[14][0]_i_6_n_0 }),
        .O({\r_reg[14][0]_i_2_n_4 ,\r_reg[14][0]_i_2_n_5 ,\r_reg[14][0]_i_2_n_6 ,\r_reg[14][0]_i_2_n_7 }),
        .S({\r[14][0]_i_7_n_0 ,\r[14][0]_i_8_n_0 ,\r[14][0]_i_9_n_0 ,\r[14][0]_i_10_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][10] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[14][8]_i_1_n_5 ),
        .Q(\r_reg[14] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][11] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[14][8]_i_1_n_4 ),
        .Q(\r_reg[14] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][12] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[14][12]_i_1_n_7 ),
        .Q(\r_reg[14] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[14][12]_i_1 
       (.CI(\r_reg[14][8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[14][12]_i_1_n_4 ,\r_reg[14][12]_i_1_n_5 ,\r_reg[14][12]_i_1_n_6 ,\r_reg[14][12]_i_1_n_7 }),
        .S({\r[14][12]_i_2_n_0 ,\r[14][12]_i_3_n_0 ,\r[14][12]_i_4_n_0 ,\r[14][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][13] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[14][12]_i_1_n_6 ),
        .Q(\r_reg[14] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][14] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[14][12]_i_1_n_5 ),
        .Q(\r_reg[14] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][15] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[14][12]_i_1_n_4 ),
        .Q(\r_reg[14] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][1] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[14][0]_i_2_n_6 ),
        .Q(\r_reg[14] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][2] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[14][0]_i_2_n_5 ),
        .Q(\r_reg[14] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][3] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[14][0]_i_2_n_4 ),
        .Q(\r_reg[14] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][4] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[14][4]_i_1_n_7 ),
        .Q(\r_reg[14] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[14][4]_i_1 
       (.CI(\r_reg[14][0]_i_2_n_0 ),
        .CO({\r_reg[14][4]_i_1_n_0 ,\r_reg[14][4]_i_1_n_1 ,\r_reg[14][4]_i_1_n_2 ,\r_reg[14][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[14][4]_i_1_n_4 ,\r_reg[14][4]_i_1_n_5 ,\r_reg[14][4]_i_1_n_6 ,\r_reg[14][4]_i_1_n_7 }),
        .S({\r[14][4]_i_2_n_0 ,\r[14][4]_i_3_n_0 ,\r[14][4]_i_4_n_0 ,\r[14][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][5] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[14][4]_i_1_n_6 ),
        .Q(\r_reg[14] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][6] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[14][4]_i_1_n_5 ),
        .Q(\r_reg[14] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][7] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[14][4]_i_1_n_4 ),
        .Q(\r_reg[14] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][8] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[14][8]_i_1_n_7 ),
        .Q(\r_reg[14] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[14][8]_i_1 
       (.CI(\r_reg[14][4]_i_1_n_0 ),
        .CO({\r_reg[14][8]_i_1_n_0 ,\r_reg[14][8]_i_1_n_1 ,\r_reg[14][8]_i_1_n_2 ,\r_reg[14][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[14][8]_i_1_n_4 ,\r_reg[14][8]_i_1_n_5 ,\r_reg[14][8]_i_1_n_6 ,\r_reg[14][8]_i_1_n_7 }),
        .S({\r[14][8]_i_2_n_0 ,\r[14][8]_i_3_n_0 ,\r[14][8]_i_4_n_0 ,\r[14][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[14][9] 
       (.C(clk),
        .CE(\r[14][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[14][8]_i_1_n_6 ),
        .Q(\r_reg[14] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][0] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[15][0]_i_2_n_7 ),
        .Q(\r_reg[15] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[15][0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[15][0]_i_2_n_0 ,\r_reg[15][0]_i_2_n_1 ,\r_reg[15][0]_i_2_n_2 ,\r_reg[15][0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r[15][0]_i_5_n_0 ,\r[15][0]_i_6_n_0 }),
        .O({\r_reg[15][0]_i_2_n_4 ,\r_reg[15][0]_i_2_n_5 ,\r_reg[15][0]_i_2_n_6 ,\r_reg[15][0]_i_2_n_7 }),
        .S({\r[15][0]_i_7_n_0 ,\r[15][0]_i_8_n_0 ,\r[15][0]_i_9_n_0 ,\r[15][0]_i_10_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][10] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[15][8]_i_1_n_5 ),
        .Q(\r_reg[15] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][11] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[15][8]_i_1_n_4 ),
        .Q(\r_reg[15] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][12] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[15][12]_i_1_n_7 ),
        .Q(\r_reg[15] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[15][12]_i_1 
       (.CI(\r_reg[15][8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[15][12]_i_1_n_4 ,\r_reg[15][12]_i_1_n_5 ,\r_reg[15][12]_i_1_n_6 ,\r_reg[15][12]_i_1_n_7 }),
        .S({\r[15][12]_i_2_n_0 ,\r[15][12]_i_3_n_0 ,\r[15][12]_i_4_n_0 ,\r[15][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][13] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[15][12]_i_1_n_6 ),
        .Q(\r_reg[15] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][14] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[15][12]_i_1_n_5 ),
        .Q(\r_reg[15] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][15] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[15][12]_i_1_n_4 ),
        .Q(\r_reg[15] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][1] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[15][0]_i_2_n_6 ),
        .Q(\r_reg[15] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][2] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[15][0]_i_2_n_5 ),
        .Q(\r_reg[15] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][3] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[15][0]_i_2_n_4 ),
        .Q(\r_reg[15] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][4] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[15][4]_i_1_n_7 ),
        .Q(\r_reg[15] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[15][4]_i_1 
       (.CI(\r_reg[15][0]_i_2_n_0 ),
        .CO({\r_reg[15][4]_i_1_n_0 ,\r_reg[15][4]_i_1_n_1 ,\r_reg[15][4]_i_1_n_2 ,\r_reg[15][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[15][4]_i_1_n_4 ,\r_reg[15][4]_i_1_n_5 ,\r_reg[15][4]_i_1_n_6 ,\r_reg[15][4]_i_1_n_7 }),
        .S({\r[15][4]_i_2_n_0 ,\r[15][4]_i_3_n_0 ,\r[15][4]_i_4_n_0 ,\r[15][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][5] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[15][4]_i_1_n_6 ),
        .Q(\r_reg[15] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][6] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[15][4]_i_1_n_5 ),
        .Q(\r_reg[15] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][7] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[15][4]_i_1_n_4 ),
        .Q(\r_reg[15] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][8] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[15][8]_i_1_n_7 ),
        .Q(\r_reg[15] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[15][8]_i_1 
       (.CI(\r_reg[15][4]_i_1_n_0 ),
        .CO({\r_reg[15][8]_i_1_n_0 ,\r_reg[15][8]_i_1_n_1 ,\r_reg[15][8]_i_1_n_2 ,\r_reg[15][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[15][8]_i_1_n_4 ,\r_reg[15][8]_i_1_n_5 ,\r_reg[15][8]_i_1_n_6 ,\r_reg[15][8]_i_1_n_7 }),
        .S({\r[15][8]_i_2_n_0 ,\r[15][8]_i_3_n_0 ,\r[15][8]_i_4_n_0 ,\r[15][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[15][9] 
       (.C(clk),
        .CE(\r[15][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[15][8]_i_1_n_6 ),
        .Q(\r_reg[15] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][0] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[4][0]_i_2_n_7 ),
        .Q(\r_reg[4] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[4][0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[4][0]_i_2_n_0 ,\r_reg[4][0]_i_2_n_1 ,\r_reg[4][0]_i_2_n_2 ,\r_reg[4][0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r[4][0]_i_7_n_0 ,\r[4][0]_i_8_n_0 }),
        .O({\r_reg[4][0]_i_2_n_4 ,\r_reg[4][0]_i_2_n_5 ,\r_reg[4][0]_i_2_n_6 ,\r_reg[4][0]_i_2_n_7 }),
        .S({\r[4][0]_i_9_n_0 ,\r[4][0]_i_10_n_0 ,\r[4][0]_i_11_n_0 ,\r[4][0]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][10] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[4][8]_i_1_n_5 ),
        .Q(\r_reg[4] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][11] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[4][8]_i_1_n_4 ),
        .Q(\r_reg[4] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][12] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[4][12]_i_1_n_7 ),
        .Q(\r_reg[4] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[4][12]_i_1 
       (.CI(\r_reg[4][8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[4][12]_i_1_n_4 ,\r_reg[4][12]_i_1_n_5 ,\r_reg[4][12]_i_1_n_6 ,\r_reg[4][12]_i_1_n_7 }),
        .S({\r[4][12]_i_2_n_0 ,\r[4][12]_i_3_n_0 ,\r[4][12]_i_4_n_0 ,\r[4][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][13] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[4][12]_i_1_n_6 ),
        .Q(\r_reg[4] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][14] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[4][12]_i_1_n_5 ),
        .Q(\r_reg[4] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][15] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[4][12]_i_1_n_4 ),
        .Q(\r_reg[4] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][1] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[4][0]_i_2_n_6 ),
        .Q(\r_reg[4] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][2] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[4][0]_i_2_n_5 ),
        .Q(\r_reg[4] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][3] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[4][0]_i_2_n_4 ),
        .Q(\r_reg[4] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][4] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[4][4]_i_1_n_7 ),
        .Q(\r_reg[4] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[4][4]_i_1 
       (.CI(\r_reg[4][0]_i_2_n_0 ),
        .CO({\r_reg[4][4]_i_1_n_0 ,\r_reg[4][4]_i_1_n_1 ,\r_reg[4][4]_i_1_n_2 ,\r_reg[4][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[4][4]_i_1_n_4 ,\r_reg[4][4]_i_1_n_5 ,\r_reg[4][4]_i_1_n_6 ,\r_reg[4][4]_i_1_n_7 }),
        .S({\r[4][4]_i_2_n_0 ,\r[4][4]_i_3_n_0 ,\r[4][4]_i_4_n_0 ,\r[4][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][5] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[4][4]_i_1_n_6 ),
        .Q(\r_reg[4] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][6] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[4][4]_i_1_n_5 ),
        .Q(\r_reg[4] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][7] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[4][4]_i_1_n_4 ),
        .Q(\r_reg[4] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][8] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[4][8]_i_1_n_7 ),
        .Q(\r_reg[4] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[4][8]_i_1 
       (.CI(\r_reg[4][4]_i_1_n_0 ),
        .CO({\r_reg[4][8]_i_1_n_0 ,\r_reg[4][8]_i_1_n_1 ,\r_reg[4][8]_i_1_n_2 ,\r_reg[4][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[4][8]_i_1_n_4 ,\r_reg[4][8]_i_1_n_5 ,\r_reg[4][8]_i_1_n_6 ,\r_reg[4][8]_i_1_n_7 }),
        .S({\r[4][8]_i_2_n_0 ,\r[4][8]_i_3_n_0 ,\r[4][8]_i_4_n_0 ,\r[4][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[4][9] 
       (.C(clk),
        .CE(\r[4][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[4][8]_i_1_n_6 ),
        .Q(\r_reg[4] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][0] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[5][0]_i_2_n_7 ),
        .Q(\r_reg[5] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[5][0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[5][0]_i_2_n_0 ,\r_reg[5][0]_i_2_n_1 ,\r_reg[5][0]_i_2_n_2 ,\r_reg[5][0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r[5][0]_i_6_n_0 ,\r[5][0]_i_7_n_0 }),
        .O({\r_reg[5][0]_i_2_n_4 ,\r_reg[5][0]_i_2_n_5 ,\r_reg[5][0]_i_2_n_6 ,\r_reg[5][0]_i_2_n_7 }),
        .S({\r[5][0]_i_8_n_0 ,\r[5][0]_i_9_n_0 ,\r[5][0]_i_10_n_0 ,\r[5][0]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][10] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[5][8]_i_1_n_5 ),
        .Q(\r_reg[5] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][11] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[5][8]_i_1_n_4 ),
        .Q(\r_reg[5] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][12] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[5][12]_i_1_n_7 ),
        .Q(\r_reg[5] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[5][12]_i_1 
       (.CI(\r_reg[5][8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[5][12]_i_1_n_4 ,\r_reg[5][12]_i_1_n_5 ,\r_reg[5][12]_i_1_n_6 ,\r_reg[5][12]_i_1_n_7 }),
        .S({\r[5][12]_i_2_n_0 ,\r[5][12]_i_3_n_0 ,\r[5][12]_i_4_n_0 ,\r[5][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][13] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[5][12]_i_1_n_6 ),
        .Q(\r_reg[5] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][14] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[5][12]_i_1_n_5 ),
        .Q(\r_reg[5] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][15] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[5][12]_i_1_n_4 ),
        .Q(\r_reg[5] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][1] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[5][0]_i_2_n_6 ),
        .Q(\r_reg[5] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][2] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[5][0]_i_2_n_5 ),
        .Q(\r_reg[5] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][3] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[5][0]_i_2_n_4 ),
        .Q(\r_reg[5] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][4] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[5][4]_i_1_n_7 ),
        .Q(\r_reg[5] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[5][4]_i_1 
       (.CI(\r_reg[5][0]_i_2_n_0 ),
        .CO({\r_reg[5][4]_i_1_n_0 ,\r_reg[5][4]_i_1_n_1 ,\r_reg[5][4]_i_1_n_2 ,\r_reg[5][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[5][4]_i_1_n_4 ,\r_reg[5][4]_i_1_n_5 ,\r_reg[5][4]_i_1_n_6 ,\r_reg[5][4]_i_1_n_7 }),
        .S({\r[5][4]_i_2_n_0 ,\r[5][4]_i_3_n_0 ,\r[5][4]_i_4_n_0 ,\r[5][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][5] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[5][4]_i_1_n_6 ),
        .Q(\r_reg[5] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][6] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[5][4]_i_1_n_5 ),
        .Q(\r_reg[5] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][7] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[5][4]_i_1_n_4 ),
        .Q(\r_reg[5] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][8] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[5][8]_i_1_n_7 ),
        .Q(\r_reg[5] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[5][8]_i_1 
       (.CI(\r_reg[5][4]_i_1_n_0 ),
        .CO({\r_reg[5][8]_i_1_n_0 ,\r_reg[5][8]_i_1_n_1 ,\r_reg[5][8]_i_1_n_2 ,\r_reg[5][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[5][8]_i_1_n_4 ,\r_reg[5][8]_i_1_n_5 ,\r_reg[5][8]_i_1_n_6 ,\r_reg[5][8]_i_1_n_7 }),
        .S({\r[5][8]_i_2_n_0 ,\r[5][8]_i_3_n_0 ,\r[5][8]_i_4_n_0 ,\r[5][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[5][9] 
       (.C(clk),
        .CE(\r[5][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[5][8]_i_1_n_6 ),
        .Q(\r_reg[5] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][0] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[6][0]_i_2_n_7 ),
        .Q(\r_reg[6] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[6][0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[6][0]_i_2_n_0 ,\r_reg[6][0]_i_2_n_1 ,\r_reg[6][0]_i_2_n_2 ,\r_reg[6][0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r[6][0]_i_6_n_0 ,\r[6][0]_i_7_n_0 }),
        .O({\r_reg[6][0]_i_2_n_4 ,\r_reg[6][0]_i_2_n_5 ,\r_reg[6][0]_i_2_n_6 ,\r_reg[6][0]_i_2_n_7 }),
        .S({\r[6][0]_i_8_n_0 ,\r[6][0]_i_9_n_0 ,\r[6][0]_i_10_n_0 ,\r[6][0]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][10] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[6][8]_i_1_n_5 ),
        .Q(\r_reg[6] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][11] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[6][8]_i_1_n_4 ),
        .Q(\r_reg[6] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][12] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[6][12]_i_1_n_7 ),
        .Q(\r_reg[6] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[6][12]_i_1 
       (.CI(\r_reg[6][8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[6][12]_i_1_n_4 ,\r_reg[6][12]_i_1_n_5 ,\r_reg[6][12]_i_1_n_6 ,\r_reg[6][12]_i_1_n_7 }),
        .S({\r[6][12]_i_2_n_0 ,\r[6][12]_i_3_n_0 ,\r[6][12]_i_4_n_0 ,\r[6][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][13] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[6][12]_i_1_n_6 ),
        .Q(\r_reg[6] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][14] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[6][12]_i_1_n_5 ),
        .Q(\r_reg[6] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][15] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[6][12]_i_1_n_4 ),
        .Q(\r_reg[6] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][1] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[6][0]_i_2_n_6 ),
        .Q(\r_reg[6] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][2] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[6][0]_i_2_n_5 ),
        .Q(\r_reg[6] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][3] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[6][0]_i_2_n_4 ),
        .Q(\r_reg[6] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][4] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[6][4]_i_1_n_7 ),
        .Q(\r_reg[6] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[6][4]_i_1 
       (.CI(\r_reg[6][0]_i_2_n_0 ),
        .CO({\r_reg[6][4]_i_1_n_0 ,\r_reg[6][4]_i_1_n_1 ,\r_reg[6][4]_i_1_n_2 ,\r_reg[6][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[6][4]_i_1_n_4 ,\r_reg[6][4]_i_1_n_5 ,\r_reg[6][4]_i_1_n_6 ,\r_reg[6][4]_i_1_n_7 }),
        .S({\r[6][4]_i_2_n_0 ,\r[6][4]_i_3_n_0 ,\r[6][4]_i_4_n_0 ,\r[6][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][5] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[6][4]_i_1_n_6 ),
        .Q(\r_reg[6] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][6] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[6][4]_i_1_n_5 ),
        .Q(\r_reg[6] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][7] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[6][4]_i_1_n_4 ),
        .Q(\r_reg[6] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][8] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[6][8]_i_1_n_7 ),
        .Q(\r_reg[6] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[6][8]_i_1 
       (.CI(\r_reg[6][4]_i_1_n_0 ),
        .CO({\r_reg[6][8]_i_1_n_0 ,\r_reg[6][8]_i_1_n_1 ,\r_reg[6][8]_i_1_n_2 ,\r_reg[6][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[6][8]_i_1_n_4 ,\r_reg[6][8]_i_1_n_5 ,\r_reg[6][8]_i_1_n_6 ,\r_reg[6][8]_i_1_n_7 }),
        .S({\r[6][8]_i_2_n_0 ,\r[6][8]_i_3_n_0 ,\r[6][8]_i_4_n_0 ,\r[6][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[6][9] 
       (.C(clk),
        .CE(\r[6][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[6][8]_i_1_n_6 ),
        .Q(\r_reg[6] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][0] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[7][0]_i_2_n_7 ),
        .Q(\r_reg[7] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[7][0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[7][0]_i_2_n_0 ,\r_reg[7][0]_i_2_n_1 ,\r_reg[7][0]_i_2_n_2 ,\r_reg[7][0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r[7][0]_i_6_n_0 ,\r[7][0]_i_7_n_0 }),
        .O({\r_reg[7][0]_i_2_n_4 ,\r_reg[7][0]_i_2_n_5 ,\r_reg[7][0]_i_2_n_6 ,\r_reg[7][0]_i_2_n_7 }),
        .S({\r[7][0]_i_8_n_0 ,\r[7][0]_i_9_n_0 ,\r[7][0]_i_10_n_0 ,\r[7][0]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][10] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[7][8]_i_1_n_5 ),
        .Q(\r_reg[7] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][11] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[7][8]_i_1_n_4 ),
        .Q(\r_reg[7] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][12] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[7][12]_i_1_n_7 ),
        .Q(\r_reg[7] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[7][12]_i_1 
       (.CI(\r_reg[7][8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[7][12]_i_1_n_4 ,\r_reg[7][12]_i_1_n_5 ,\r_reg[7][12]_i_1_n_6 ,\r_reg[7][12]_i_1_n_7 }),
        .S({\r[7][12]_i_2_n_0 ,\r[7][12]_i_3_n_0 ,\r[7][12]_i_4_n_0 ,\r[7][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][13] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[7][12]_i_1_n_6 ),
        .Q(\r_reg[7] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][14] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[7][12]_i_1_n_5 ),
        .Q(\r_reg[7] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][15] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[7][12]_i_1_n_4 ),
        .Q(\r_reg[7] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][1] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[7][0]_i_2_n_6 ),
        .Q(\r_reg[7] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][2] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[7][0]_i_2_n_5 ),
        .Q(\r_reg[7] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][3] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[7][0]_i_2_n_4 ),
        .Q(\r_reg[7] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][4] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[7][4]_i_1_n_7 ),
        .Q(\r_reg[7] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[7][4]_i_1 
       (.CI(\r_reg[7][0]_i_2_n_0 ),
        .CO({\r_reg[7][4]_i_1_n_0 ,\r_reg[7][4]_i_1_n_1 ,\r_reg[7][4]_i_1_n_2 ,\r_reg[7][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[7][4]_i_1_n_4 ,\r_reg[7][4]_i_1_n_5 ,\r_reg[7][4]_i_1_n_6 ,\r_reg[7][4]_i_1_n_7 }),
        .S({\r[7][4]_i_2_n_0 ,\r[7][4]_i_3_n_0 ,\r[7][4]_i_4_n_0 ,\r[7][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][5] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[7][4]_i_1_n_6 ),
        .Q(\r_reg[7] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][6] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[7][4]_i_1_n_5 ),
        .Q(\r_reg[7] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][7] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[7][4]_i_1_n_4 ),
        .Q(\r_reg[7] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][8] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[7][8]_i_1_n_7 ),
        .Q(\r_reg[7] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[7][8]_i_1 
       (.CI(\r_reg[7][4]_i_1_n_0 ),
        .CO({\r_reg[7][8]_i_1_n_0 ,\r_reg[7][8]_i_1_n_1 ,\r_reg[7][8]_i_1_n_2 ,\r_reg[7][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[7][8]_i_1_n_4 ,\r_reg[7][8]_i_1_n_5 ,\r_reg[7][8]_i_1_n_6 ,\r_reg[7][8]_i_1_n_7 }),
        .S({\r[7][8]_i_2_n_0 ,\r[7][8]_i_3_n_0 ,\r[7][8]_i_4_n_0 ,\r[7][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[7][9] 
       (.C(clk),
        .CE(\r[7][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[7][8]_i_1_n_6 ),
        .Q(\r_reg[7] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][0] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[8][0]_i_2_n_7 ),
        .Q(\r_reg[8] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[8][0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[8][0]_i_2_n_0 ,\r_reg[8][0]_i_2_n_1 ,\r_reg[8][0]_i_2_n_2 ,\r_reg[8][0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r[8][0]_i_7_n_0 ,\r[8][0]_i_8_n_0 }),
        .O({\r_reg[8][0]_i_2_n_4 ,\r_reg[8][0]_i_2_n_5 ,\r_reg[8][0]_i_2_n_6 ,\r_reg[8][0]_i_2_n_7 }),
        .S({\r[8][0]_i_9_n_0 ,\r[8][0]_i_10_n_0 ,\r[8][0]_i_11_n_0 ,\r[8][0]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][10] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[8][8]_i_1_n_5 ),
        .Q(\r_reg[8] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][11] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[8][8]_i_1_n_4 ),
        .Q(\r_reg[8] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][12] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[8][12]_i_1_n_7 ),
        .Q(\r_reg[8] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[8][12]_i_1 
       (.CI(\r_reg[8][8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[8][12]_i_1_n_4 ,\r_reg[8][12]_i_1_n_5 ,\r_reg[8][12]_i_1_n_6 ,\r_reg[8][12]_i_1_n_7 }),
        .S({\r[8][12]_i_2_n_0 ,\r[8][12]_i_3_n_0 ,\r[8][12]_i_4_n_0 ,\r[8][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][13] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[8][12]_i_1_n_6 ),
        .Q(\r_reg[8] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][14] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[8][12]_i_1_n_5 ),
        .Q(\r_reg[8] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][15] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[8][12]_i_1_n_4 ),
        .Q(\r_reg[8] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][1] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[8][0]_i_2_n_6 ),
        .Q(\r_reg[8] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][2] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[8][0]_i_2_n_5 ),
        .Q(\r_reg[8] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][3] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[8][0]_i_2_n_4 ),
        .Q(\r_reg[8] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][4] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[8][4]_i_1_n_7 ),
        .Q(\r_reg[8] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[8][4]_i_1 
       (.CI(\r_reg[8][0]_i_2_n_0 ),
        .CO({\r_reg[8][4]_i_1_n_0 ,\r_reg[8][4]_i_1_n_1 ,\r_reg[8][4]_i_1_n_2 ,\r_reg[8][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[8][4]_i_1_n_4 ,\r_reg[8][4]_i_1_n_5 ,\r_reg[8][4]_i_1_n_6 ,\r_reg[8][4]_i_1_n_7 }),
        .S({\r[8][4]_i_2_n_0 ,\r[8][4]_i_3_n_0 ,\r[8][4]_i_4_n_0 ,\r[8][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][5] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[8][4]_i_1_n_6 ),
        .Q(\r_reg[8] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][6] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[8][4]_i_1_n_5 ),
        .Q(\r_reg[8] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][7] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[8][4]_i_1_n_4 ),
        .Q(\r_reg[8] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][8] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[8][8]_i_1_n_7 ),
        .Q(\r_reg[8] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[8][8]_i_1 
       (.CI(\r_reg[8][4]_i_1_n_0 ),
        .CO({\r_reg[8][8]_i_1_n_0 ,\r_reg[8][8]_i_1_n_1 ,\r_reg[8][8]_i_1_n_2 ,\r_reg[8][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[8][8]_i_1_n_4 ,\r_reg[8][8]_i_1_n_5 ,\r_reg[8][8]_i_1_n_6 ,\r_reg[8][8]_i_1_n_7 }),
        .S({\r[8][8]_i_2_n_0 ,\r[8][8]_i_3_n_0 ,\r[8][8]_i_4_n_0 ,\r[8][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[8][9] 
       (.C(clk),
        .CE(\r[8][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[8][8]_i_1_n_6 ),
        .Q(\r_reg[8] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][0] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[9][0]_i_2_n_7 ),
        .Q(\r_reg[9] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[9][0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\r_reg[9][0]_i_2_n_0 ,\r_reg[9][0]_i_2_n_1 ,\r_reg[9][0]_i_2_n_2 ,\r_reg[9][0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\r[9][0]_i_6_n_0 ,\r[9][0]_i_7_n_0 }),
        .O({\r_reg[9][0]_i_2_n_4 ,\r_reg[9][0]_i_2_n_5 ,\r_reg[9][0]_i_2_n_6 ,\r_reg[9][0]_i_2_n_7 }),
        .S({\r[9][0]_i_8_n_0 ,\r[9][0]_i_9_n_0 ,\r[9][0]_i_10_n_0 ,\r[9][0]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][10] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[9][8]_i_1_n_5 ),
        .Q(\r_reg[9] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][11] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[9][8]_i_1_n_4 ),
        .Q(\r_reg[9] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][12] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[9][12]_i_1_n_7 ),
        .Q(\r_reg[9] [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[9][12]_i_1 
       (.CI(\r_reg[9][8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[9][12]_i_1_n_4 ,\r_reg[9][12]_i_1_n_5 ,\r_reg[9][12]_i_1_n_6 ,\r_reg[9][12]_i_1_n_7 }),
        .S({\r[9][12]_i_2_n_0 ,\r[9][12]_i_3_n_0 ,\r[9][12]_i_4_n_0 ,\r[9][12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][13] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[9][12]_i_1_n_6 ),
        .Q(\r_reg[9] [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][14] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[9][12]_i_1_n_5 ),
        .Q(\r_reg[9] [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][15] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[9][12]_i_1_n_4 ),
        .Q(\r_reg[9] [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][1] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[9][0]_i_2_n_6 ),
        .Q(\r_reg[9] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][2] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[9][0]_i_2_n_5 ),
        .Q(\r_reg[9] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][3] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\r_reg[9][0]_i_2_n_4 ),
        .Q(\r_reg[9] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][4] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[9][4]_i_1_n_7 ),
        .Q(\r_reg[9] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[9][4]_i_1 
       (.CI(\r_reg[9][0]_i_2_n_0 ),
        .CO({\r_reg[9][4]_i_1_n_0 ,\r_reg[9][4]_i_1_n_1 ,\r_reg[9][4]_i_1_n_2 ,\r_reg[9][4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[9][4]_i_1_n_4 ,\r_reg[9][4]_i_1_n_5 ,\r_reg[9][4]_i_1_n_6 ,\r_reg[9][4]_i_1_n_7 }),
        .S({\r[9][4]_i_2_n_0 ,\r[9][4]_i_3_n_0 ,\r[9][4]_i_4_n_0 ,\r[9][4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][5] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[9][4]_i_1_n_6 ),
        .Q(\r_reg[9] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][6] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\r_reg[9][4]_i_1_n_5 ),
        .Q(\r_reg[9] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][7] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[9][4]_i_1_n_4 ),
        .Q(\r_reg[9] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][8] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[9][8]_i_1_n_7 ),
        .Q(\r_reg[9] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \r_reg[9][8]_i_1 
       (.CI(\r_reg[9][4]_i_1_n_0 ),
        .CO({\r_reg[9][8]_i_1_n_0 ,\r_reg[9][8]_i_1_n_1 ,\r_reg[9][8]_i_1_n_2 ,\r_reg[9][8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\r_reg[9][8]_i_1_n_4 ,\r_reg[9][8]_i_1_n_5 ,\r_reg[9][8]_i_1_n_6 ,\r_reg[9][8]_i_1_n_7 }),
        .S({\r[9][8]_i_2_n_0 ,\r[9][8]_i_3_n_0 ,\r[9][8]_i_4_n_0 ,\r[9][8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \r_reg[9][9] 
       (.C(clk),
        .CE(\r[9][0]_i_1_n_0 ),
        .CLR(\src[8]_i_2_n_0 ),
        .D(\r_reg[9][8]_i_1_n_6 ),
        .Q(\r_reg[9] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    rd_INST_0
       (.I0(rd_INST_0_i_1_n_0),
        .I1(rd_INST_0_i_2_n_0),
        .O(rd));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF8A000000)) 
    rd_INST_0_i_1
       (.I0(rd_INST_0_i_3_n_0),
        .I1(soc[1]),
        .I2(soc[2]),
        .I3(eqOp135_in),
        .I4(p_2_in88_in),
        .I5(rd_INST_0_i_6_n_0),
        .O(rd_INST_0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0FFF1F0F0F0F0)) 
    rd_INST_0_i_10
       (.I0(rd_INST_0_i_21_n_0),
        .I1(rd_INST_0_i_16_n_0),
        .I2(rd_INST_0_i_22_n_0),
        .I3(eqOp105_in),
        .I4(\dout[13]_INST_0_i_3_n_0 ),
        .I5(p_2_in88_in),
        .O(rd_INST_0_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEEEEEFEEEE)) 
    rd_INST_0_i_11
       (.I0(rd_INST_0_i_23_n_0),
        .I1(rd_INST_0_i_24_n_0),
        .I2(state[1]),
        .I3(state[4]),
        .I4(\FSM_sequential_state[1]_i_5_n_0 ),
        .I5(rd_INST_0_i_25_n_0),
        .O(nstate[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0507)) 
    rd_INST_0_i_12
       (.I0(rd_INST_0_i_26_n_0),
        .I1(rd_INST_0_i_27_n_0),
        .I2(state[4]),
        .I3(state[3]),
        .O(nstate[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000040055555555)) 
    rd_INST_0_i_13
       (.I0(state[4]),
        .I1(rd_INST_0_i_28_n_0),
        .I2(state[1]),
        .I3(state[0]),
        .I4(state[2]),
        .I5(rd_INST_0_i_29_n_0),
        .O(rd_INST_0_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEFEFEFFFEFE)) 
    rd_INST_0_i_14
       (.I0(rd_INST_0_i_30_n_0),
        .I1(rd_INST_0_i_31_n_0),
        .I2(rd_INST_0_i_32_n_0),
        .I3(state[4]),
        .I4(state[3]),
        .I5(rd_INST_0_i_33_n_0),
        .O(nstate[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF0000F444)) 
    rd_INST_0_i_15
       (.I0(rd_INST_0_i_34_n_0),
        .I1(state[3]),
        .I2(\FSM_sequential_state[1]_i_8_n_0 ),
        .I3(rd_INST_0_i_35_n_0),
        .I4(state[4]),
        .I5(rd_INST_0_i_36_n_0),
        .O(nstate[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h808080FFFFFF80FF)) 
    rd_INST_0_i_16
       (.I0(\r_code[0]_i_1_n_0 ),
        .I1(\r_code[1]_i_1_n_0 ),
        .I2(\addr[15]_INST_0_i_11_n_0 ),
        .I3(r_code[7]),
        .I4(p_2_in88_in),
        .I5(din[7]),
        .O(rd_INST_0_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hAFBF)) 
    rd_INST_0_i_17
       (.I0(rd_INST_0_i_21_n_0),
        .I1(din[15]),
        .I2(p_2_in88_in),
        .I3(din[14]),
        .O(rd_INST_0_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000080)) 
    rd_INST_0_i_18
       (.I0(state[1]),
        .I1(state[0]),
        .I2(state[3]),
        .I3(state[4]),
        .I4(state[2]),
        .O(rd_INST_0_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02AAAAAA)) 
    rd_INST_0_i_19
       (.I0(lbe_INST_0_i_8_n_0),
        .I1(as[1]),
        .I2(\r_code[0]_i_1_n_0 ),
        .I3(\addr[15]_INST_0_i_11_n_0 ),
        .I4(\r_code[1]_i_1_n_0 ),
        .O(rd_INST_0_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF1)) 
    rd_INST_0_i_2
       (.I0(rd_INST_0_i_7_n_0),
        .I1(rd_INST_0_i_8_n_0),
        .I2(rd_INST_0_i_9_n_0),
        .I3(rd_INST_0_i_10_n_0),
        .O(rd_INST_0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFF7)) 
    rd_INST_0_i_20
       (.I0(state[2]),
        .I1(state[3]),
        .I2(state[4]),
        .I3(state[0]),
        .I4(state[1]),
        .O(rd_INST_0_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAA02AAAA)) 
    rd_INST_0_i_21
       (.I0(lbe_INST_0_i_8_n_0),
        .I1(as[1]),
        .I2(soc[1]),
        .I3(\r_code[11]_i_1_n_0 ),
        .I4(soc[2]),
        .I5(\r_code[10]_i_1_n_0 ),
        .O(rd_INST_0_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000008000F)) 
    rd_INST_0_i_22
       (.I0(eqOp113_in),
        .I1(eqOp135_in),
        .I2(rd_INST_0_i_37_n_0),
        .I3(state[2]),
        .I4(state[0]),
        .I5(state[1]),
        .O(rd_INST_0_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h02A800A802A000A0)) 
    rd_INST_0_i_23
       (.I0(rd_INST_0_i_38_n_0),
        .I1(state[0]),
        .I2(state[4]),
        .I3(state[3]),
        .I4(\FSM_sequential_state[1]_i_5_n_0 ),
        .I5(rd_INST_0_i_39_n_0),
        .O(rd_INST_0_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h02000C0002000000)) 
    rd_INST_0_i_24
       (.I0(rd_INST_0_i_40_n_0),
        .I1(state[0]),
        .I2(state[4]),
        .I3(state[1]),
        .I4(state[2]),
        .I5(rd_INST_0_i_41_n_0),
        .O(rd_INST_0_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    rd_INST_0_i_25
       (.I0(state[0]),
        .I1(state[2]),
        .O(rd_INST_0_i_25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h066F064F6F6F6F6F)) 
    rd_INST_0_i_26
       (.I0(state[0]),
        .I1(state[2]),
        .I2(state[1]),
        .I3(\FSM_sequential_state[1]_i_5_n_0 ),
        .I4(rd_INST_0_i_16_n_0),
        .I5(state[3]),
        .O(rd_INST_0_i_26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111333333033333)) 
    rd_INST_0_i_27
       (.I0(rd_INST_0_i_42_n_0),
        .I1(rd_INST_0_i_43_n_0),
        .I2(rd_INST_0_i_44_n_0),
        .I3(state[1]),
        .I4(state[0]),
        .I5(state[2]),
        .O(rd_INST_0_i_27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 rd_INST_0_i_28
       (.I0(rd_INST_0_i_45_n_0),
        .I1(rd_INST_0_i_46_n_0),
        .O(rd_INST_0_i_28_n_0),
        .S(eqOp135_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 rd_INST_0_i_29
       (.I0(rd_INST_0_i_47_n_0),
        .I1(rd_INST_0_i_48_n_0),
        .O(rd_INST_0_i_29_n_0),
        .S(state[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0C000CAACCAACCAA)) 
    rd_INST_0_i_3
       (.I0(r_code[5]),
        .I1(din[5]),
        .I2(din[1]),
        .I3(p_2_in88_in),
        .I4(r_code[1]),
        .I5(\addr[15]_INST_0_i_11_n_0 ),
        .O(rd_INST_0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1101110100010101)) 
    rd_INST_0_i_30
       (.I0(state[3]),
        .I1(state[4]),
        .I2(state[0]),
        .I3(state[1]),
        .I4(state[2]),
        .I5(girq),
        .O(rd_INST_0_i_30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F00000400040)) 
    rd_INST_0_i_31
       (.I0(state[3]),
        .I1(rd_INST_0_i_49_n_0),
        .I2(state[0]),
        .I3(state[1]),
        .I4(state[4]),
        .I5(state[2]),
        .O(rd_INST_0_i_31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000004340)) 
    rd_INST_0_i_32
       (.I0(state[3]),
        .I1(state[4]),
        .I2(state[0]),
        .I3(girq),
        .I4(state[1]),
        .I5(state[2]),
        .O(rd_INST_0_i_32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h023303FF02FFFFFF)) 
    rd_INST_0_i_33
       (.I0(rd_INST_0_i_16_n_0),
        .I1(girq),
        .I2(rd_INST_0_i_50_n_0),
        .I3(state[1]),
        .I4(state[0]),
        .I5(state[2]),
        .O(rd_INST_0_i_33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h043C3CFF)) 
    rd_INST_0_i_34
       (.I0(rd_INST_0_i_16_n_0),
        .I1(state[1]),
        .I2(state[2]),
        .I3(state[0]),
        .I4(girq),
        .O(rd_INST_0_i_34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 rd_INST_0_i_35
       (.I0(rd_INST_0_i_51_n_0),
        .I1(rd_INST_0_i_52_n_0),
        .O(rd_INST_0_i_35_n_0),
        .S(eqOp135_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000000060E6)) 
    rd_INST_0_i_36
       (.I0(state[2]),
        .I1(state[1]),
        .I2(girq),
        .I3(state[0]),
        .I4(state[4]),
        .I5(state[3]),
        .O(rd_INST_0_i_36_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    rd_INST_0_i_37
       (.I0(state[4]),
        .I1(state[3]),
        .O(rd_INST_0_i_37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    rd_INST_0_i_38
       (.I0(state[1]),
        .I1(state[2]),
        .O(rd_INST_0_i_38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 rd_INST_0_i_39
       (.I0(rd_INST_0_i_53_n_0),
        .I1(rd_INST_0_i_54_n_0),
        .O(rd_INST_0_i_39_n_0),
        .S(eqOp135_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00020000)) 
    rd_INST_0_i_4
       (.I0(\dout[13]_INST_0_i_3_n_0 ),
        .I1(\r_code[10]_i_1_n_0 ),
        .I2(\r_code[11]_i_1_n_0 ),
        .I3(doc[1]),
        .I4(doc[0]),
        .O(eqOp135_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    rd_INST_0_i_40
       (.I0(\sr_reg_n_0_[4] ),
        .I1(state[3]),
        .I2(state_reg[4]),
        .I3(girq),
        .O(rd_INST_0_i_40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B0)) 
    rd_INST_0_i_41
       (.I0(rd_INST_0_i_16_n_0),
        .I1(state[3]),
        .I2(\sr_reg_n_0_[4] ),
        .I3(girq),
        .O(rd_INST_0_i_41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    rd_INST_0_i_42
       (.I0(\sr_reg_n_0_[4] ),
        .I1(girq),
        .O(rd_INST_0_i_42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h54040000)) 
    rd_INST_0_i_43
       (.I0(girq),
        .I1(state_reg[1]),
        .I2(state[0]),
        .I3(\sr_reg_n_0_[4] ),
        .I4(state[1]),
        .O(rd_INST_0_i_43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 rd_INST_0_i_44
       (.I0(rd_INST_0_i_57_n_0),
        .I1(rd_INST_0_i_58_n_0),
        .O(rd_INST_0_i_44_n_0),
        .S(eqOp135_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFFFEFEFCF00CFCF)) 
    rd_INST_0_i_45
       (.I0(rd_INST_0_i_50_n_0),
        .I1(girq),
        .I2(\FSM_sequential_state[3]_i_6_n_0 ),
        .I3(doc[1]),
        .I4(\dout[13]_INST_0_i_3_n_0 ),
        .I5(state_reg[3]),
        .O(rd_INST_0_i_45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000000000EA)) 
    rd_INST_0_i_46
       (.I0(girq),
        .I1(rd_INST_0_i_50_n_0),
        .I2(state_reg[3]),
        .I3(nstate1),
        .I4(\FSM_sequential_state[3]_i_8_n_0 ),
        .I5(rd_INST_0_i_19_n_0),
        .O(rd_INST_0_i_46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF54FF55F5FFF5FFF)) 
    rd_INST_0_i_47
       (.I0(girq),
        .I1(state[4]),
        .I2(state[1]),
        .I3(state[0]),
        .I4(state[3]),
        .I5(state[2]),
        .O(rd_INST_0_i_47_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h050A0805)) 
    rd_INST_0_i_48
       (.I0(state[0]),
        .I1(rd_INST_0_i_16_n_0),
        .I2(girq),
        .I3(state[1]),
        .I4(state[2]),
        .O(rd_INST_0_i_48_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 rd_INST_0_i_49
       (.I0(rd_INST_0_i_60_n_0),
        .I1(rd_INST_0_i_61_n_0),
        .O(rd_INST_0_i_49_n_0),
        .S(eqOp135_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000004)) 
    rd_INST_0_i_5
       (.I0(state[1]),
        .I1(\state[0]_repN ),
        .I2(\state[2]_repN ),
        .I3(\state[3]_repN ),
        .I4(\state[4]_repN ),
        .O(p_2_in88_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5455)) 
    rd_INST_0_i_50
       (.I0(\sr_reg_n_0_[4] ),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\addr[15]_INST_0_i_11_n_0 ),
        .O(rd_INST_0_i_50_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8AAA8AA20A02000)) 
    rd_INST_0_i_51
       (.I0(\FSM_sequential_state[3]_i_6_n_0 ),
        .I1(doc[1]),
        .I2(state_reg[2]),
        .I3(\dout[13]_INST_0_i_3_n_0 ),
        .I4(rd_INST_0_i_50_n_0),
        .I5(girq),
        .O(rd_INST_0_i_51_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEFEFEEEFEFEEEE)) 
    rd_INST_0_i_52
       (.I0(\FSM_sequential_state[3]_i_8_n_0 ),
        .I1(nstate1),
        .I2(rd_INST_0_i_19_n_0),
        .I3(rd_INST_0_i_50_n_0),
        .I4(girq),
        .I5(state_reg[2]),
        .O(rd_INST_0_i_52_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBAAABFAA30003000)) 
    rd_INST_0_i_53
       (.I0(\sr_reg_n_0_[4] ),
        .I1(doc[1]),
        .I2(\dout[13]_INST_0_i_3_n_0 ),
        .I3(state_reg[4]),
        .I4(\pc[15]_i_8_n_0 ),
        .I5(rd_INST_0_i_63_n_0),
        .O(rd_INST_0_i_53_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001000100010000)) 
    rd_INST_0_i_54
       (.I0(girq),
        .I1(rd_INST_0_i_19_n_0),
        .I2(\FSM_sequential_state[3]_i_8_n_0 ),
        .I3(nstate1),
        .I4(\sr_reg_n_0_[4] ),
        .I5(rd_INST_0_i_64_n_0),
        .O(rd_INST_0_i_54_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000640)) 
    rd_INST_0_i_55
       (.I0(state[0]),
        .I1(state[1]),
        .I2(state[2]),
        .I3(state[4]),
        .I4(state[3]),
        .O(state_reg[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h50154502)) 
    rd_INST_0_i_56
       (.I0(state[4]),
        .I1(state[2]),
        .I2(state[0]),
        .I3(state[1]),
        .I4(state[3]),
        .O(state_reg[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF2000000)) 
    rd_INST_0_i_57
       (.I0(state_reg[1]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\sr_reg_n_0_[4] ),
        .I3(\dout[5]_INST_0_i_10_n_0 ),
        .I4(rd_INST_0_i_65_n_0),
        .I5(rd_INST_0_i_66_n_0),
        .O(rd_INST_0_i_57_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF40CF40CF40CFCF)) 
    rd_INST_0_i_58
       (.I0(soc[0]),
        .I1(soc[1]),
        .I2(soc[2]),
        .I3(rd_INST_0_i_19_n_0),
        .I4(rd_INST_0_i_67_n_0),
        .I5(girq),
        .O(rd_INST_0_i_58_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h54105402)) 
    rd_INST_0_i_59
       (.I0(state[4]),
        .I1(state[1]),
        .I2(state[0]),
        .I3(state[3]),
        .I4(state[2]),
        .O(state_reg[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAABBAEAAE)) 
    rd_INST_0_i_6
       (.I0(\addr[15]_INST_0_i_17_n_0 ),
        .I1(state[2]),
        .I2(state[1]),
        .I3(state[0]),
        .I4(state[3]),
        .I5(state[4]),
        .O(rd_INST_0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3300B00033B3B0B3)) 
    rd_INST_0_i_60
       (.I0(rd_INST_0_i_50_n_0),
        .I1(rd_INST_0_i_63_n_0),
        .I2(state_reg[0]),
        .I3(\dout[13]_INST_0_i_3_n_0 ),
        .I4(doc[1]),
        .I5(rd_INST_0_i_69_n_0),
        .O(rd_INST_0_i_60_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0404555504045554)) 
    rd_INST_0_i_61
       (.I0(\FSM_sequential_state[3]_i_8_n_0 ),
        .I1(rd_INST_0_i_3_n_0),
        .I2(nstate1),
        .I3(rd_INST_0_i_70_n_0),
        .I4(rd_INST_0_i_19_n_0),
        .I5(girq),
        .O(rd_INST_0_i_61_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h41045106)) 
    rd_INST_0_i_62
       (.I0(state[4]),
        .I1(state[1]),
        .I2(state[3]),
        .I3(state[2]),
        .I4(state[0]),
        .O(state_reg[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4440004044444444)) 
    rd_INST_0_i_63
       (.I0(girq),
        .I1(\FSM_sequential_state[3]_i_6_n_0 ),
        .I2(r_code[13]),
        .I3(p_2_in88_in),
        .I4(din[13]),
        .I5(\dout[13]_INST_0_i_3_n_0 ),
        .O(rd_INST_0_i_63_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000041400)) 
    rd_INST_0_i_64
       (.I0(state[3]),
        .I1(state[4]),
        .I2(state[2]),
        .I3(state[1]),
        .I4(state[0]),
        .I5(\pc[15]_i_8_n_0 ),
        .O(rd_INST_0_i_64_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    rd_INST_0_i_65
       (.I0(rd_INST_0_i_16_n_0),
        .I1(girq),
        .O(rd_INST_0_i_65_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF1F111F1F1111111)) 
    rd_INST_0_i_66
       (.I0(\FSM_sequential_state[3]_i_6_n_0 ),
        .I1(eqOp105_in),
        .I2(\dout[13]_INST_0_i_3_n_0 ),
        .I3(doc[1]),
        .I4(\FSM_sequential_state[1]_i_5_n_0 ),
        .I5(state_reg[1]),
        .O(rd_INST_0_i_66_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00045555)) 
    rd_INST_0_i_67
       (.I0(\sr_reg_n_0_[4] ),
        .I1(\addr[15]_INST_0_i_11_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_code[0]_i_1_n_0 ),
        .I4(state_reg[1]),
        .O(rd_INST_0_i_67_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00170570)) 
    rd_INST_0_i_68
       (.I0(state[2]),
        .I1(state[1]),
        .I2(state[0]),
        .I3(state[4]),
        .I4(state[3]),
        .O(state_reg[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hE2E2E2E2E200E2E2)) 
    rd_INST_0_i_69
       (.I0(r_code[5]),
        .I1(p_2_in88_in),
        .I2(din[5]),
        .I3(\r_code[10]_i_1_n_0 ),
        .I4(soc[2]),
        .I5(\r_code[11]_i_1_n_0 ),
        .O(rd_INST_0_i_69_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    rd_INST_0_i_7
       (.I0(nstate[4]),
        .I1(nstate[1]),
        .I2(rd_INST_0_i_13_n_0),
        .I3(nstate[0]),
        .I4(nstate[2]),
        .O(rd_INST_0_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000020802280A28)) 
    rd_INST_0_i_70
       (.I0(rd_INST_0_i_50_n_0),
        .I1(state[3]),
        .I2(state[4]),
        .I3(state[0]),
        .I4(state[1]),
        .I5(state[2]),
        .O(rd_INST_0_i_70_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5D005D5D5D5D5D5D)) 
    rd_INST_0_i_8
       (.I0(rd_INST_0_i_16_n_0),
        .I1(rd_INST_0_i_17_n_0),
        .I2(rd_INST_0_i_18_n_0),
        .I3(rd_INST_0_i_19_n_0),
        .I4(eqOp135_in),
        .I5(p_2_in88_in),
        .O(rd_INST_0_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF4544FFFF)) 
    rd_INST_0_i_9
       (.I0(rd_INST_0_i_16_n_0),
        .I1(rd_INST_0_i_18_n_0),
        .I2(\dout[13]_INST_0_i_3_n_0 ),
        .I3(p_2_in88_in),
        .I4(rd_INST_0_i_20_n_0),
        .I5(\addr[15]_INST_0_i_5_n_0 ),
        .O(rd_INST_0_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4444544455555555)) 
    \sp[0]_i_1 
       (.I0(halt),
        .I1(\sp[0]_i_3_n_0 ),
        .I2(soc[1]),
        .I3(\sp[0]_i_4_n_0 ),
        .I4(\sp[0]_i_5_n_0 ),
        .I5(\sp[0]_i_6_n_0 ),
        .O(\sp[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[0]_i_10 
       (.I0(\dout[1]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[1]),
        .I3(sp_reg[1]),
        .I4(sp19_out),
        .O(sp));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[0]_i_11 
       (.I0(sp_reg[0]),
        .I1(sp19_out),
        .I2(plusOp[0]),
        .I3(\sp[0]_i_6_n_0 ),
        .I4(\dout[0]_INST_0_i_1_n_0 ),
        .O(\sp[0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFACCFA)) 
    \sp[0]_i_12 
       (.I0(r_code[1]),
        .I1(din[1]),
        .I2(r_code[2]),
        .I3(p_2_in88_in),
        .I4(din[2]),
        .O(\sp[0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sp[0]_i_16 
       (.I0(sp_reg[1]),
        .O(\sp[0]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF0400FFFF)) 
    \sp[0]_i_3 
       (.I0(\r_code[3]_i_1_n_0 ),
        .I1(\r_code[0]_i_1_n_0 ),
        .I2(\sp[0]_i_12_n_0 ),
        .I3(\r[4][0]_i_5_n_0 ),
        .I4(rd_INST_0_i_20_n_0),
        .I5(sp19_out),
        .O(\sp[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEF000000000000)) 
    \sp[0]_i_4 
       (.I0(\r[10][0]_i_5_n_0 ),
        .I1(\r_code[11]_i_1_n_0 ),
        .I2(soc[1]),
        .I3(as[1]),
        .I4(as[0]),
        .I5(\addr[15]_INST_0_i_17_n_0 ),
        .O(\sp[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFCFFFFFFFCFAFA)) 
    \sp[0]_i_5 
       (.I0(r_code[11]),
        .I1(din[11]),
        .I2(soc[2]),
        .I3(din[10]),
        .I4(p_2_in88_in),
        .I5(r_code[10]),
        .O(\sp[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFBFF)) 
    \sp[0]_i_6 
       (.I0(rd_INST_0_i_8_n_0),
        .I1(\addr[3]_INST_0_i_9_n_0 ),
        .I2(\r_code[1]_i_1_n_0 ),
        .I3(\r_code[0]_i_1_n_0 ),
        .I4(\r_code[3]_i_1_n_0 ),
        .O(\sp[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0802)) 
    \sp[0]_i_7 
       (.I0(nstate[2]),
        .I1(nstate[1]),
        .I2(nstate[4]),
        .I3(rd_INST_0_i_13_n_0),
        .O(sp19_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[0]_i_8 
       (.I0(\dout[3]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[3]),
        .I3(sp_reg[3]),
        .I4(sp19_out),
        .O(\sp[0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[0]_i_9 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[2]),
        .I3(sp_reg[2]),
        .I4(sp19_out),
        .O(\sp[0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h74777444)) 
    \sp[12]_i_2 
       (.I0(sp_reg[15]),
        .I1(sp19_out),
        .I2(plusOp[15]),
        .I3(\sp[0]_i_6_n_0 ),
        .I4(\dout[15]_INST_0_i_3_n_0 ),
        .O(\sp[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[12]_i_3 
       (.I0(\dout[14]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[14]),
        .I3(sp_reg[14]),
        .I4(sp19_out),
        .O(\sp[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[12]_i_4 
       (.I0(\dout[13]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[13]),
        .I3(sp_reg[13]),
        .I4(sp19_out),
        .O(\sp[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[12]_i_5 
       (.I0(\dout[12]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[12]),
        .I3(sp_reg[12]),
        .I4(sp19_out),
        .O(\sp[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[4]_i_2 
       (.I0(\dout[7]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[7]),
        .I3(sp_reg[7]),
        .I4(sp19_out),
        .O(\sp[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[4]_i_3 
       (.I0(\dout[6]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[6]),
        .I3(sp_reg[6]),
        .I4(sp19_out),
        .O(\sp[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[4]_i_4 
       (.I0(\dout[5]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[5]),
        .I3(sp_reg[5]),
        .I4(sp19_out),
        .O(\sp[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[4]_i_5 
       (.I0(\dout[4]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[4]),
        .I3(sp_reg[4]),
        .I4(sp19_out),
        .O(\sp[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[8]_i_2 
       (.I0(\dout[11]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[11]),
        .I3(sp_reg[11]),
        .I4(sp19_out),
        .O(\sp[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[8]_i_3 
       (.I0(\dout[10]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[10]),
        .I3(sp_reg[10]),
        .I4(sp19_out),
        .O(\sp[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[8]_i_4 
       (.I0(\dout[9]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[9]),
        .I3(sp_reg[9]),
        .I4(sp19_out),
        .O(\sp[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FFE2E2)) 
    \sp[8]_i_5 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(\sp[0]_i_6_n_0 ),
        .I2(plusOp[8]),
        .I3(sp_reg[8]),
        .I4(sp19_out),
        .O(\sp[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[0] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[0]_i_2_n_7 ),
        .Q(sp_reg[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sp_reg[0]_i_13 
       (.CI(\<const0>__0__0 ),
        .CO({\sp_reg[0]_i_13_n_0 ,\sp_reg[0]_i_13_n_1 ,\sp_reg[0]_i_13_n_2 ,\sp_reg[0]_i_13_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,sp_reg[1],\<const0>__0__0 }),
        .O(plusOp[3:0]),
        .S({sp_reg[3:2],\sp[0]_i_16_n_0 ,sp_reg[0]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sp_reg[0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\sp_reg[0]_i_2_n_0 ,\sp_reg[0]_i_2_n_1 ,\sp_reg[0]_i_2_n_2 ,\sp_reg[0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({sp19_out,sp19_out,sp19_out,\<const0>__0__0 }),
        .O({\sp_reg[0]_i_2_n_4 ,\sp_reg[0]_i_2_n_5 ,\sp_reg[0]_i_2_n_6 ,\sp_reg[0]_i_2_n_7 }),
        .S({\sp[0]_i_8_n_0 ,\sp[0]_i_9_n_0 ,sp,\sp[0]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[10] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[8]_i_1_n_5 ),
        .Q(sp_reg[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[11] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[8]_i_1_n_4 ),
        .Q(sp_reg[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[12] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[12]_i_1_n_7 ),
        .Q(sp_reg[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sp_reg[12]_i_1 
       (.CI(\sp_reg[8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,sp19_out,sp19_out,sp19_out}),
        .O({\sp_reg[12]_i_1_n_4 ,\sp_reg[12]_i_1_n_5 ,\sp_reg[12]_i_1_n_6 ,\sp_reg[12]_i_1_n_7 }),
        .S({\sp[12]_i_2_n_0 ,\sp[12]_i_3_n_0 ,\sp[12]_i_4_n_0 ,\sp[12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sp_reg[12]_i_6 
       (.CI(\sp_reg[8]_i_6_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(plusOp[15:12]),
        .S(sp_reg[15:12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[13] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[12]_i_1_n_6 ),
        .Q(sp_reg[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[14] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[12]_i_1_n_5 ),
        .Q(sp_reg[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[15] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[12]_i_1_n_4 ),
        .Q(sp_reg[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[1] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[0]_i_2_n_6 ),
        .Q(sp_reg[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[2] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[0]_i_2_n_5 ),
        .Q(sp_reg[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[3] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[0]_i_2_n_4 ),
        .Q(sp_reg[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[4] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[4]_i_1_n_7 ),
        .Q(sp_reg[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sp_reg[4]_i_1 
       (.CI(\sp_reg[0]_i_2_n_0 ),
        .CO({\sp_reg[4]_i_1_n_0 ,\sp_reg[4]_i_1_n_1 ,\sp_reg[4]_i_1_n_2 ,\sp_reg[4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({sp19_out,sp19_out,sp19_out,sp19_out}),
        .O({\sp_reg[4]_i_1_n_4 ,\sp_reg[4]_i_1_n_5 ,\sp_reg[4]_i_1_n_6 ,\sp_reg[4]_i_1_n_7 }),
        .S({\sp[4]_i_2_n_0 ,\sp[4]_i_3_n_0 ,\sp[4]_i_4_n_0 ,\sp[4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sp_reg[4]_i_6 
       (.CI(\sp_reg[0]_i_13_n_0 ),
        .CO({\sp_reg[4]_i_6_n_0 ,\sp_reg[4]_i_6_n_1 ,\sp_reg[4]_i_6_n_2 ,\sp_reg[4]_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(plusOp[7:4]),
        .S(sp_reg[7:4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[5] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[4]_i_1_n_6 ),
        .Q(sp_reg[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[6] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[4]_i_1_n_5 ),
        .Q(sp_reg[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[7] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[4]_i_1_n_4 ),
        .Q(sp_reg[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[8] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[8]_i_1_n_7 ),
        .Q(sp_reg[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sp_reg[8]_i_1 
       (.CI(\sp_reg[4]_i_1_n_0 ),
        .CO({\sp_reg[8]_i_1_n_0 ,\sp_reg[8]_i_1_n_1 ,\sp_reg[8]_i_1_n_2 ,\sp_reg[8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({sp19_out,sp19_out,sp19_out,sp19_out}),
        .O({\sp_reg[8]_i_1_n_4 ,\sp_reg[8]_i_1_n_5 ,\sp_reg[8]_i_1_n_6 ,\sp_reg[8]_i_1_n_7 }),
        .S({\sp[8]_i_2_n_0 ,\sp[8]_i_3_n_0 ,\sp[8]_i_4_n_0 ,\sp[8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sp_reg[8]_i_6 
       (.CI(\sp_reg[4]_i_6_n_0 ),
        .CO({\sp_reg[8]_i_6_n_0 ,\sp_reg[8]_i_6_n_1 ,\sp_reg[8]_i_6_n_2 ,\sp_reg[8]_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(plusOp[11:8]),
        .S(sp_reg[11:8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sp_reg[9] 
       (.C(clk),
        .CE(\sp[0]_i_1_n_0 ),
        .CLR(\src[15]_i_3_n_0 ),
        .D(\sp_reg[8]_i_1_n_6 ),
        .Q(sp_reg[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \sr[0]_i_1 
       (.I0(din[0]),
        .I1(p_0_in6_in),
        .I2(\sr[0]_i_2_n_0 ),
        .I3(\sr[2]_i_3_n_0 ),
        .I4(sr_reg_n_0_),
        .O(sr));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000077477747)) 
    \sr[0]_i_2 
       (.I0(\sr[0]_i_3_n_0 ),
        .I1(eqOp135_in),
        .I2(\sr[0]_i_4_n_0 ),
        .I3(\sr[0]_i_5_n_0 ),
        .I4(\dout[0]_INST_0_i_1_n_0 ),
        .I5(sr1),
        .O(\sr[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000B8FFFFFFB8)) 
    \sr[0]_i_3 
       (.I0(\dout[2]_INST_0_i_45_n_0 ),
        .I1(bw),
        .I2(\dout[9]_INST_0_i_11_n_0 ),
        .I3(soc[0]),
        .I4(soc[2]),
        .I5(\dout[7]_INST_0_i_7_n_0_repN ),
        .O(\sr[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAFEFFAAAABABB)) 
    \sr[0]_i_4 
       (.I0(\sr[0]_i_6_n_0 ),
        .I1(\dout[15]_INST_0_i_23_n_0 ),
        .I2(\dout[15]_INST_0_i_19_n_0 ),
        .I3(\sr[1]_i_11_n_0 ),
        .I4(\sr[0]_i_7_n_0 ),
        .I5(\dout[14]_INST_0_i_18_n_0 ),
        .O(\sr[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF8FFF88888888888)) 
    \sr[0]_i_5 
       (.I0(\dout[4]_INST_0_i_7_n_0 ),
        .I1(\sr_reg[0]_i_8_n_3 ),
        .I2(\sr_reg[0]_i_9_n_3 ),
        .I3(bw),
        .I4(sr_reg[0]),
        .I5(\dout[15]_INST_0_i_31_n_0 ),
        .O(\sr[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \sr[0]_i_6 
       (.I0(\dout[15]_INST_0_i_31_n_0 ),
        .I1(\dout[4]_INST_0_i_7_n_0 ),
        .O(\sr[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F444FFF44444444)) 
    \sr[0]_i_7 
       (.I0(\sr_reg[0]_i_11_n_3 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\sr_reg[0]_i_12_n_3 ),
        .I3(bw),
        .I4(\sr_reg[0]_i_13_n_3 ),
        .I5(\dout[15]_INST_0_i_20_n_0 ),
        .O(\sr[0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[10]_i_1 
       (.I0(din[10]),
        .I1(p_0_in6_in),
        .I2(\dout[10]_INST_0_i_1_n_0 ),
        .O(\sr[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[11]_i_1 
       (.I0(din[11]),
        .I1(p_0_in6_in),
        .I2(\dout[11]_INST_0_i_1_n_0 ),
        .O(\sr[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[12]_i_1 
       (.I0(din[12]),
        .I1(p_0_in6_in),
        .I2(\dout[12]_INST_0_i_1_n_0 ),
        .O(\sr[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[13]_i_1 
       (.I0(din[13]),
        .I1(p_0_in6_in),
        .I2(\dout[13]_INST_0_i_1_n_0 ),
        .O(\sr[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[14]_i_1 
       (.I0(din[14]),
        .I1(p_0_in6_in),
        .I2(\dout[14]_INST_0_i_1_n_0 ),
        .O(\sr[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h0E)) 
    \sr[15]_i_1 
       (.I0(p_0_in6_in),
        .I1(sr1),
        .I2(halt),
        .O(\sr[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[15]_i_2 
       (.I0(din[15]),
        .I1(p_0_in6_in),
        .I2(\dout[15]_INST_0_i_3_n_0 ),
        .O(\sr[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000020)) 
    \sr[15]_i_3 
       (.I0(state[2]),
        .I1(state[1]),
        .I2(state[3]),
        .I3(state[4]),
        .I4(state[0]),
        .O(p_0_in6_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0040)) 
    \sr[15]_i_4 
       (.I0(\r_code[0]_i_1_n_0 ),
        .I1(\r_code[1]_i_1_n_0 ),
        .I2(\addr[15]_INST_0_i_11_n_0 ),
        .I3(rd_INST_0_i_8_n_0),
        .O(sr1));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88B8FFFF88B80000)) 
    \sr[1]_i_1 
       (.I0(din[1]),
        .I1(p_0_in6_in),
        .I2(\sr[1]_i_2_n_0 ),
        .I3(\sr[1]_i_3_n_0 ),
        .I4(\sr[2]_i_3_n_0 ),
        .I5(\sr_reg_n_0_[1] ),
        .O(\sr[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \sr[1]_i_10 
       (.I0(\dout[15]_INST_0_i_26_n_4 ),
        .I1(\dout[15]_INST_0_i_26_n_7 ),
        .I2(\sr[1]_i_23_n_0 ),
        .I3(\dout[15]_INST_0_i_56_n_4 ),
        .I4(\dout[15]_INST_0_i_26_n_6 ),
        .I5(\dout[15]_INST_0_i_26_n_5 ),
        .O(\sr[1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFFFFE)) 
    \sr[1]_i_11 
       (.I0(\sr[1]_i_24_n_0 ),
        .I1(\sr[1]_i_25_n_0 ),
        .I2(\dout[11]_INST_0_i_29_n_0 ),
        .I3(\sr[1]_i_26_n_0 ),
        .I4(\sr[1]_i_27_n_0 ),
        .I5(\sr[1]_i_28_n_0 ),
        .O(\sr[1]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[1]_i_12 
       (.I0(\sr[1]_i_29_n_0 ),
        .I1(\sr[1]_i_30_n_0 ),
        .I2(\sr[1]_i_31_n_0 ),
        .I3(\dout[2]_INST_0_i_11_n_6 ),
        .I4(\dout[4]_INST_0_i_11_n_4 ),
        .I5(\dout[2]_INST_0_i_11_n_5 ),
        .O(\sr[1]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF9FFFF)) 
    \sr[1]_i_13 
       (.I0(\dout[9]_INST_0_i_4_n_0 ),
        .I1(\dout[9]_INST_0_i_5_n_0 ),
        .I2(\sr[1]_i_32_n_0 ),
        .I3(\dout[10]_INST_0_i_5_n_0 ),
        .I4(\dout[12]_INST_0_i_5_n_0 ),
        .I5(\dout[11]_INST_0_i_5_n_0 ),
        .O(\sr[1]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA995A9A99595A995)) 
    \sr[1]_i_14 
       (.I0(\dout[15]_INST_0_i_44_n_0 ),
        .I1(\dout[14]_INST_0_i_27_n_0 ),
        .I2(L[13]),
        .I3(L[12]),
        .I4(\dout[4]_INST_0_i_13_n_0 ),
        .I5(\dout[9]_INST_0_i_5_n_0 ),
        .O(\sr[1]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4D00B2FFB2FF4D00)) 
    \sr[1]_i_15 
       (.I0(\dout[9]_INST_0_i_5_n_0 ),
        .I1(\dout[4]_INST_0_i_13_n_0 ),
        .I2(L[12]),
        .I3(\dout[15]_INST_0_i_45_n_0 ),
        .I4(\dout[14]_INST_0_i_16_n_0 ),
        .I5(\dout[15]_INST_0_i_44_n_0 ),
        .O(\sr[1]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[1]_i_16 
       (.I0(\sr[1]_i_33_n_0 ),
        .I1(\sr[1]_i_34_n_0 ),
        .I2(\sr[1]_i_35_n_0 ),
        .I3(\dout[4]_INST_0_i_44_n_6 ),
        .I4(\dout[15]_INST_0_i_30_n_7 ),
        .I5(\dout[15]_INST_0_i_71_n_5 ),
        .O(\sr[1]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \sr[1]_i_17 
       (.I0(\dout[15]_INST_0_i_66_n_4 ),
        .I1(\dout[15]_INST_0_i_29_n_4 ),
        .I2(\dout[15]_INST_0_i_66_n_5 ),
        .I3(\sr[1]_i_36_n_0 ),
        .O(\sr[1]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFD)) 
    \sr[1]_i_18 
       (.I0(\dout[4]_INST_0_i_7_n_0 ),
        .I1(\sr[1]_i_37_n_0 ),
        .I2(\dout[15]_INST_0_i_61_n_4 ),
        .I3(\dout[2]_INST_0_i_6_n_6 ),
        .I4(\dout[15]_INST_0_i_28_n_5 ),
        .I5(\dout[4]_INST_0_i_6_n_5 ),
        .O(\sr[1]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \sr[1]_i_19 
       (.I0(p_13_in),
        .I1(\dout[4]_INST_0_i_6_n_6 ),
        .I2(\dout[2]_INST_0_i_6_n_7 ),
        .I3(\dout[15]_INST_0_i_28_n_7 ),
        .I4(\sr[1]_i_38_n_0 ),
        .O(\sr[1]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \sr[1]_i_2 
       (.I0(\dout[1]_INST_0_i_1_n_0 ),
        .I1(sr1),
        .O(\sr[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \sr[1]_i_20 
       (.I0(\dout[6]_INST_0_i_5_n_0 ),
        .I1(sr_reg_n_0_),
        .I2(soc[1]),
        .O(\sr[1]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \sr[1]_i_21 
       (.I0(\dout[15]_INST_0_i_15_n_0 ),
        .I1(\dout[4]_INST_0_i_13_n_0 ),
        .I2(\dout[14]_INST_0_i_27_n_0 ),
        .I3(\sr[1]_i_39_n_0 ),
        .I4(\sr[1]_i_40_n_0 ),
        .I5(\sr[1]_i_41_n_0 ),
        .O(\sr[1]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[1]_i_22 
       (.I0(\dout[15]_INST_0_i_25_n_5 ),
        .I1(\dout[15]_INST_0_i_25_n_6 ),
        .I2(\dout[15]_INST_0_i_25_n_7 ),
        .I3(\dout[15]_INST_0_i_25_n_4 ),
        .O(\sr[1]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \sr[1]_i_23 
       (.I0(\dout[15]_INST_0_i_56_n_6 ),
        .I1(\sr[1]_i_42_n_0 ),
        .I2(\dout[2]_INST_0_i_30_n_7 ),
        .I3(\dout[2]_INST_0_i_30_n_5 ),
        .I4(\dout[15]_INST_0_i_56_n_7 ),
        .I5(\dout[15]_INST_0_i_56_n_5 ),
        .O(\sr[1]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \sr[1]_i_24 
       (.I0(L[11]),
        .I1(\dout[11]_INST_0_i_16_n_0 ),
        .O(\sr[1]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \sr[1]_i_25 
       (.I0(L[10]),
        .I1(\dout[2]_INST_0_i_12_n_0 ),
        .O(\sr[1]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[1]_i_26 
       (.I0(\sr[1]_i_43_n_0 ),
        .I1(\dout[9]_INST_0_i_19_n_0 ),
        .I2(\dout[4]_INST_0_i_32_n_0 ),
        .I3(\sr[1]_i_44_n_0 ),
        .I4(\dout[6]_INST_0_i_13_n_0 ),
        .I5(\dout[14]_INST_0_i_10_n_0 ),
        .O(\sr[1]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[1]_i_27 
       (.I0(\sr[1]_i_45_n_0 ),
        .I1(\dout[7]_INST_0_i_13_n_0 ),
        .I2(\dout[0]_INST_0_i_11_n_0 ),
        .I3(\dout[2]_INST_0_i_43_n_0 ),
        .I4(\dout[2]_INST_0_i_27_n_0 ),
        .I5(\dout[14]_INST_0_i_16_n_0 ),
        .O(\sr[1]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBAAA)) 
    \sr[1]_i_28 
       (.I0(\dout[15]_INST_0_i_20_n_0 ),
        .I1(\sr[1]_i_46_n_0 ),
        .I2(\dout[14]_INST_0_i_10_n_0 ),
        .I3(\dout[15]_INST_0_i_43_n_0 ),
        .O(\sr[1]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[1]_i_29 
       (.I0(\dout[15]_INST_0_i_39_n_7 ),
        .I1(\dout[4]_INST_0_i_11_n_5 ),
        .I2(\dout[15]_INST_0_i_21_n_6 ),
        .I3(\dout[15]_INST_0_i_39_n_6 ),
        .O(\sr[1]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFF00AE)) 
    \sr[1]_i_3 
       (.I0(\sr[1]_i_4_n_0 ),
        .I1(\sr[1]_i_5_n_0 ),
        .I2(\sr[1]_i_6_n_0 ),
        .I3(\sr[1]_i_7_n_0 ),
        .I4(eqOp135_in),
        .I5(\sr[1]_i_8_n_0 ),
        .O(\sr[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[1]_i_30 
       (.I0(\dout[15]_INST_0_i_21_n_7 ),
        .I1(\dout[15]_INST_0_i_39_n_4 ),
        .I2(\dout[15]_INST_0_i_39_n_5 ),
        .I3(\dout[4]_INST_0_i_11_n_6 ),
        .O(\sr[1]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[1]_i_31 
       (.I0(\dout[2]_INST_0_i_11_n_7 ),
        .I1(\dout[15]_INST_0_i_21_n_4 ),
        .I2(\dout[4]_INST_0_i_11_n_7 ),
        .I3(\dout[2]_INST_0_i_11_n_4 ),
        .O(\sr[1]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    \sr[1]_i_32 
       (.I0(\dout[6]_INST_0_i_9_n_0 ),
        .I1(\dout[5]_INST_0_i_8_n_0 ),
        .I2(\dout[7]_INST_0_i_9_n_0 ),
        .I3(\sr[1]_i_47_n_0 ),
        .I4(\dout[8]_INST_0_i_5_n_0 ),
        .O(\sr[1]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[1]_i_33 
       (.I0(\dout[15]_INST_0_i_30_n_4 ),
        .I1(bw),
        .I2(\dout[2]_INST_0_i_31_n_4 ),
        .I3(\dout[15]_INST_0_i_30_n_6 ),
        .I4(\dout[2]_INST_0_i_31_n_6 ),
        .I5(\dout[4]_INST_0_i_44_n_7 ),
        .O(\sr[1]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[1]_i_34 
       (.I0(\dout[15]_INST_0_i_71_n_7 ),
        .I1(\dout[4]_INST_0_i_44_n_4 ),
        .I2(\dout[15]_INST_0_i_71_n_6 ),
        .I3(\dout[2]_INST_0_i_31_n_5 ),
        .O(\sr[1]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[1]_i_35 
       (.I0(\dout[15]_INST_0_i_30_n_5 ),
        .I1(\dout[4]_INST_0_i_44_n_5 ),
        .I2(\dout[15]_INST_0_i_71_n_4 ),
        .I3(\dout[2]_INST_0_i_31_n_7 ),
        .O(\sr[1]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFD)) 
    \sr[1]_i_36 
       (.I0(bw),
        .I1(\dout[15]_INST_0_i_29_n_6 ),
        .I2(\dout[15]_INST_0_i_29_n_7 ),
        .I3(\dout[15]_INST_0_i_29_n_5 ),
        .I4(\dout[15]_INST_0_i_66_n_6 ),
        .I5(\dout[15]_INST_0_i_66_n_7 ),
        .O(\sr[1]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[1]_i_37 
       (.I0(\dout[15]_INST_0_i_28_n_6 ),
        .I1(\dout[4]_INST_0_i_6_n_7 ),
        .I2(\dout[15]_INST_0_i_61_n_7 ),
        .I3(\dout[4]_INST_0_i_6_n_4 ),
        .O(\sr[1]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[1]_i_38 
       (.I0(\dout[15]_INST_0_i_61_n_5 ),
        .I1(\dout[15]_INST_0_i_61_n_6 ),
        .I2(\dout[2]_INST_0_i_6_n_4 ),
        .I3(\dout[2]_INST_0_i_6_n_5 ),
        .O(\sr[1]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF4FFF0)) 
    \sr[1]_i_39_rewire_rewire 
       (.I0(\dout[5]_INST_0_i_11_n_0 ),
        .I1(\dout[5]_INST_0_i_5_n_0 ),
        .I2(\dout[4]_INST_0_i_5_n_0 ),
        .I3(\dout[0]_INST_0_i_5_n_0 ),
        .I4(\dout[6]_INST_0_i_7_n_0 ),
        .I5(\dout[2]_INST_0_i_5_n_0 ),
        .O(\sr[1]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEEEFFFEEEEEEEE)) 
    \sr[1]_i_4 
       (.I0(\dout[4]_INST_0_i_7_n_0 ),
        .I1(\dout[15]_INST_0_i_31_n_0 ),
        .I2(\sr[1]_i_9_n_0 ),
        .I3(bw),
        .I4(\sr[1]_i_10_n_0 ),
        .I5(\dout[15]_INST_0_i_20_n_0 ),
        .O(\sr[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFB3)) 
    \sr[1]_i_40_rewire 
       (.I0(\dout[4]_INST_0_i_16_n_0 ),
        .I1(\dout[9]_INST_0_i_11_n_0 ),
        .I2(\dout[13]_INST_0_i_20_n_0 ),
        .I3(\dout[11]_INST_0_i_26_n_0 ),
        .O(\sr[1]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \sr[1]_i_41 
       (.I0(\dout[14]_INST_0_i_9_n_0 ),
        .I1(\dout[2]_INST_0_i_12_n_0 ),
        .I2(\dout[11]_INST_0_i_16_n_0 ),
        .I3(\dout[9]_INST_0_i_14_n_0 ),
        .O(\sr[1]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[1]_i_42 
       (.I0(\dout[4]_INST_0_i_43_n_7 ),
        .I1(\dout[4]_INST_0_i_43_n_4 ),
        .I2(\dout[4]_INST_0_i_43_n_6 ),
        .I3(\dout[4]_INST_0_i_43_n_5 ),
        .I4(\dout[2]_INST_0_i_30_n_4 ),
        .I5(\dout[2]_INST_0_i_30_n_6 ),
        .O(\sr[1]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \sr[1]_i_43 
       (.I0(\dout[15]_INST_0_i_36_n_0 ),
        .I1(\dout[15]_INST_0_i_48_n_0 ),
        .O(\sr[1]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \sr[1]_i_44 
       (.I0(\dout[2]_INST_0_i_14_n_0 ),
        .I1(\dout[2]_INST_0_i_13_n_0 ),
        .O(\sr[1]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \sr[1]_i_45 
       (.I0(L[12]),
        .I1(\dout[4]_INST_0_i_13_n_0 ),
        .O(\sr[1]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFFFFFFFFFF)) 
    \sr[1]_i_46 
       (.I0(\sr[1]_i_48_n_0 ),
        .I1(\sr[1]_i_49_n_0 ),
        .I2(\sr[1]_i_50_n_0 ),
        .I3(\dout[4]_INST_0_i_40_n_0 ),
        .I4(\dout[15]_INST_0_i_80_n_0 ),
        .I5(\dout[2]_INST_0_i_33_n_0 ),
        .O(\sr[1]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \sr[1]_i_47 
       (.I0(\dout[0]_INST_0_i_8_n_0 ),
        .I1(\dout[1]_INST_0_i_8_n_0 ),
        .I2(\dout[2]_INST_0_i_9_n_0 ),
        .I3(\dout[4]_INST_0_i_10_n_0 ),
        .I4(\dout[15]_INST_0_i_23_n_0 ),
        .I5(\dout[3]_INST_0_i_8_n_0 ),
        .O(\sr[1]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FFFFFFF)) 
    \sr[1]_i_48 
       (.I0(\dout[4]_INST_0_i_20_n_0 ),
        .I1(\dout[4]_INST_0_i_5_n_0 ),
        .I2(\dout[15]_INST_0_i_45_n_0 ),
        .I3(\dout[4]_INST_0_i_39_n_0 ),
        .I4(\dout[15]_INST_0_i_79_n_0 ),
        .O(\sr[1]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h6FFFFFFFFFFF6FFF)) 
    \sr[1]_i_49 
       (.I0(\dout[5]_INST_0_i_12_n_0_repN ),
        .I1(\dout[13]_INST_0_i_20_n_0_repN ),
        .I2(\dout[2]_INST_0_i_35_n_0 ),
        .I3(\dout[15]_INST_0_i_78_n_0 ),
        .I4(\dout[2]_INST_0_i_14_n_0 ),
        .I5(\dout[11]_INST_0_i_26_n_0 ),
        .O(\sr[1]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEEF0EE)) 
    \sr[1]_i_5 
       (.I0(\sr[1]_i_11_n_0 ),
        .I1(\dout[15]_INST_0_i_23_n_0 ),
        .I2(\sr[1]_i_12_n_0 ),
        .I3(\dout[15]_INST_0_i_19_n_0 ),
        .I4(\dout[15]_INST_0_i_21_n_5 ),
        .O(\sr[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF99FFFFFFFFFFFFF)) 
    \sr[1]_i_50 
       (.I0(L[8]),
        .I1(\dout[9]_INST_0_i_11_n_0 ),
        .I2(L[12]),
        .I3(\dout[4]_INST_0_i_13_n_0 ),
        .I4(\dout[15]_INST_0_i_44_n_0 ),
        .I5(\dout[2]_INST_0_i_34_n_0 ),
        .O(\sr[1]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001000000010202)) 
    \sr[1]_i_6 
       (.I0(\dout[14]_INST_0_i_29_n_0 ),
        .I1(\dout[15]_INST_0_i_22_n_0 ),
        .I2(\sr[1]_i_13_n_0 ),
        .I3(\sr[1]_i_14_n_0 ),
        .I4(\dout[14]_INST_0_i_18_n_0 ),
        .I5(\sr[1]_i_15_n_0 ),
        .O(\sr[1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hD0FFD0D0)) 
    \sr[1]_i_7 
       (.I0(\sr[1]_i_16_n_0 ),
        .I1(\sr[1]_i_17_n_0 ),
        .I2(\dout[15]_INST_0_i_31_n_0 ),
        .I3(\sr[1]_i_18_n_0 ),
        .I4(\sr[1]_i_19_n_0 ),
        .O(\sr[1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAABAAABAAABAAAAA)) 
    \sr[1]_i_8 
       (.I0(sr1),
        .I1(\dout[7]_INST_0_i_7_n_0_repN ),
        .I2(eqOp135_in),
        .I3(\sr[1]_i_20_n_0 ),
        .I4(\dout[7]_INST_0_i_6_n_0 ),
        .I5(\sr[1]_i_21_n_0 ),
        .O(\sr[1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \sr[1]_i_9 
       (.I0(\dout[15]_INST_0_i_51_n_6 ),
        .I1(\dout[15]_INST_0_i_51_n_4 ),
        .I2(\dout[15]_INST_0_i_51_n_7 ),
        .I3(\dout[15]_INST_0_i_51_n_5 ),
        .I4(\sr[1]_i_22_n_0 ),
        .O(\sr[1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \sr[2]_i_1 
       (.I0(din[2]),
        .I1(p_0_in6_in),
        .I2(\sr[2]_i_2_n_0 ),
        .I3(\sr[2]_i_3_n_0 ),
        .I4(p_1_in122_in),
        .O(\sr[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \sr[2]_i_2 
       (.I0(\dout[2]_INST_0_i_1_n_0 ),
        .I1(sr1),
        .I2(\sr[2]_i_4_n_0 ),
        .I3(\sr[2]_i_5_n_0 ),
        .I4(\sr[2]_i_6_n_0 ),
        .I5(\dout[15]_INST_0_i_13_n_0 ),
        .O(\sr[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00FE)) 
    \sr[2]_i_3 
       (.I0(p_0_in6_in),
        .I1(\sr[8]_i_7_n_0 ),
        .I2(\sr[2]_i_7_n_0 ),
        .I3(halt),
        .O(\sr[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0AAA88880A008888)) 
    \sr[2]_i_4 
       (.I0(eqOp135_in),
        .I1(\dout[7]_INST_0_i_7_n_0_repN ),
        .I2(\dout[15]_INST_0_i_15_n_0 ),
        .I3(soc[1]),
        .I4(\sr[2]_i_8_n_0 ),
        .I5(sr_reg_n_0_),
        .O(\sr[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEECCEECCEECCEEFC)) 
    \sr[2]_i_5 
       (.I0(\dout[15]_INST_0_i_22_n_0 ),
        .I1(\sr[2]_i_9_n_0 ),
        .I2(\dout[15]_INST_0_i_16_n_0 ),
        .I3(\dout[15]_INST_0_i_23_n_0 ),
        .I4(\dout[15]_INST_0_i_19_n_0 ),
        .I5(\dout[15]_INST_0_i_20_n_0 ),
        .O(\sr[2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[2]_i_6 
       (.I0(eqOp135_in),
        .I1(\dout[4]_INST_0_i_7_n_0 ),
        .I2(\dout[15]_INST_0_i_31_n_0 ),
        .O(\sr[2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAA008A0)) 
    \sr[2]_i_7 
       (.I0(\sr[8]_i_6_n_0 ),
        .I1(doc[0]),
        .I2(doc[3]),
        .I3(doc[2]),
        .I4(doc[1]),
        .O(\sr[2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00053305)) 
    \sr[2]_i_8 
       (.I0(r_code[7]),
        .I1(din[7]),
        .I2(r_code[9]),
        .I3(p_2_in88_in),
        .I4(din[9]),
        .O(\sr[2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0FFF00088888888)) 
    \sr[2]_i_9 
       (.I0(\dout[15]_INST_0_i_21_n_4 ),
        .I1(\dout[15]_INST_0_i_19_n_0 ),
        .I2(\dout[15]_INST_0_i_25_n_4 ),
        .I3(bw),
        .I4(\dout[15]_INST_0_i_26_n_4 ),
        .I5(\dout[15]_INST_0_i_20_n_0 ),
        .O(\sr[2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[3]_i_1 
       (.I0(din[3]),
        .I1(p_0_in6_in),
        .I2(\dout[3]_INST_0_i_1_n_0 ),
        .O(\sr[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[4]_i_1 
       (.I0(din[4]),
        .I1(p_0_in6_in),
        .I2(\dout[4]_INST_0_i_1_n_0 ),
        .O(\sr[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[5]_i_1 
       (.I0(din[5]),
        .I1(p_0_in6_in),
        .I2(\dout[5]_INST_0_i_1_n_0 ),
        .O(\sr[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[6]_i_1 
       (.I0(din[6]),
        .I1(p_0_in6_in),
        .I2(\dout[6]_INST_0_i_1_n_0 ),
        .O(\sr[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[7]_i_1 
       (.I0(din[7]),
        .I1(p_0_in6_in),
        .I2(\dout[7]_INST_0_i_1_n_0 ),
        .O(\sr[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFACAF0000ACA0)) 
    \sr[8]_i_1 
       (.I0(din[8]),
        .I1(\sr[8]_i_2_n_0 ),
        .I2(p_0_in6_in),
        .I3(\sr[8]_i_3_n_0 ),
        .I4(halt),
        .I5(\sr_reg_n_0_[8] ),
        .O(\sr[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[8]_i_10 
       (.I0(\dout[15]_INST_0_i_29_n_4 ),
        .I1(bw),
        .I2(\dout[15]_INST_0_i_30_n_4 ),
        .O(\sr[8]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8B8B8B8B88BB8888)) 
    \sr[8]_i_2 
       (.I0(\dout[8]_INST_0_i_1_n_0 ),
        .I1(sr1),
        .I2(\sr[8]_i_4_n_0 ),
        .I3(\sr[8]_i_5_n_0 ),
        .I4(doc[2]),
        .I5(doc[3]),
        .O(\sr[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFE3C80000)) 
    \sr[8]_i_3 
       (.I0(doc[0]),
        .I1(doc[2]),
        .I2(doc[1]),
        .I3(doc[3]),
        .I4(\sr[8]_i_6_n_0 ),
        .I5(\sr[8]_i_7_n_0 ),
        .O(\sr[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F3F3F3F3F3F3F2A)) 
    \sr[8]_i_4 
       (.I0(\dout[15]_INST_0_i_43_n_0 ),
        .I1(\dout[15]_INST_0_i_36_n_0 ),
        .I2(\dout[14]_INST_0_i_10_n_0 ),
        .I3(\dout[15]_INST_0_i_21_n_4 ),
        .I4(doc[1]),
        .I5(doc[2]),
        .O(\sr[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FFFF757F757F)) 
    \sr[8]_i_5 
       (.I0(doc[0]),
        .I1(\dout[15]_INST_0_i_38_n_0 ),
        .I2(p_13_in),
        .I3(\dout[15]_INST_0_i_36_n_0 ),
        .I4(\sr[8]_i_8_n_0 ),
        .I5(doc[1]),
        .O(\sr[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000090FFFFFFFF)) 
    \sr[8]_i_6 
       (.I0(state[2]),
        .I1(state[1]),
        .I2(state[3]),
        .I3(state[4]),
        .I4(state[0]),
        .I5(rd_INST_0_i_8_n_0),
        .O(\sr[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8888A8AA88888888)) 
    \sr[8]_i_7 
       (.I0(\sr[8]_i_6_n_0 ),
        .I1(sr1),
        .I2(soc[1]),
        .I3(soc[0]),
        .I4(soc[2]),
        .I5(eqOp135_in),
        .O(\sr[8]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1F101F1F1F101010)) 
    \sr[8]_i_8 
       (.I0(\dout[15]_INST_0_i_43_n_0 ),
        .I1(\sr[8]_i_9_n_0 ),
        .I2(doc[0]),
        .I3(\dout[15]_INST_0_i_38_n_0 ),
        .I4(\sr[8]_i_10_n_0 ),
        .I5(\dout[15]_INST_0_i_36_n_0 ),
        .O(\sr[8]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[8]_i_9 
       (.I0(\dout[15]_INST_0_i_25_n_4 ),
        .I1(bw),
        .I2(\dout[15]_INST_0_i_26_n_4 ),
        .O(\sr[8]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[9]_i_1 
       (.I0(din[9]),
        .I1(p_0_in6_in),
        .I2(\dout[9]_INST_0_i_1_n_0 ),
        .O(\sr[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(sr),
        .Q(sr_reg_n_0_));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sr_reg[0]_i_10 
       (.CI(\dout[15]_INST_0_i_30_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(sr_reg),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\sr_reg[0]_i_8_n_3 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sr_reg[0]_i_11 
       (.CI(\dout[15]_INST_0_i_21_n_0 ),
        .CO({\sr_reg[0]_i_11_n_0 ,\sr_reg[0]_i_11_n_1 ,\sr_reg[0]_i_11_n_2 ,\sr_reg[0]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sr_reg[0]_i_12 
       (.CI(\dout[15]_INST_0_i_25_n_0 ),
        .CO({\sr_reg[0]_i_12_n_0 ,\sr_reg[0]_i_12_n_1 ,\sr_reg[0]_i_12_n_2 ,\sr_reg[0]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sr_reg[0]_i_13 
       (.CI(\dout[15]_INST_0_i_26_n_0 ),
        .CO({\sr_reg[0]_i_13_n_0 ,\sr_reg[0]_i_13_n_1 ,\sr_reg[0]_i_13_n_2 ,\sr_reg[0]_i_13_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sr_reg[0]_i_8 
       (.CI(\dout[15]_INST_0_i_28_n_0 ),
        .CO({\sr_reg[0]_i_8_n_0 ,\sr_reg[0]_i_8_n_1 ,\sr_reg[0]_i_8_n_2 ,\sr_reg[0]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \sr_reg[0]_i_9 
       (.CI(\dout[15]_INST_0_i_29_n_0 ),
        .CO({\sr_reg[0]_i_9_n_0 ,\sr_reg[0]_i_9_n_1 ,\sr_reg[0]_i_9_n_2 ,\sr_reg[0]_i_9_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[10] 
       (.C(clk),
        .CE(\sr[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[10]_i_1_n_0 ),
        .Q(\sr_reg_n_0_[10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[11] 
       (.C(clk),
        .CE(\sr[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[11]_i_1_n_0 ),
        .Q(\sr_reg_n_0_[11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[12] 
       (.C(clk),
        .CE(\sr[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[12]_i_1_n_0 ),
        .Q(\sr_reg_n_0_[12] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[13] 
       (.C(clk),
        .CE(\sr[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[13]_i_1_n_0 ),
        .Q(\sr_reg_n_0_[13] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[14] 
       (.C(clk),
        .CE(\sr[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[14]_i_1_n_0 ),
        .Q(\sr_reg_n_0_[14] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[15] 
       (.C(clk),
        .CE(\sr[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[15]_i_2_n_0 ),
        .Q(\sr_reg_n_0_[15] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[1]_i_1_n_0 ),
        .Q(\sr_reg_n_0_[1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[2]_i_1_n_0 ),
        .Q(p_1_in122_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[3] 
       (.C(clk),
        .CE(\sr[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[3]_i_1_n_0 ),
        .Q(p_1_in108_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[4] 
       (.C(clk),
        .CE(\sr[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[4]_i_1_n_0 ),
        .Q(\sr_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[5] 
       (.C(clk),
        .CE(\sr[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[5]_i_1_n_0 ),
        .Q(\sr_reg_n_0_[5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[6] 
       (.C(clk),
        .CE(\sr[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[6]_i_1_n_0 ),
        .Q(\sr_reg_n_0_[6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[7] 
       (.C(clk),
        .CE(\sr[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[7]_i_1_n_0 ),
        .Q(\sr_reg_n_0_[7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[8]_i_1_n_0 ),
        .Q(\sr_reg_n_0_[8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[9] 
       (.C(clk),
        .CE(\sr[15]_i_1_n_0 ),
        .CLR(\FSM_sequential_state[4]_i_3_n_0 ),
        .D(\sr[9]_i_1_n_0 ),
        .Q(\sr_reg_n_0_[9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBF80)) 
    \src[0]_i_1 
       (.I0(din[8]),
        .I1(r_a0),
        .I2(bw),
        .I3(din[0]),
        .O(data4[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h2A)) 
    \src[10]_i_1 
       (.I0(din[10]),
        .I1(r_a0),
        .I2(bw),
        .O(data4[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h2A)) 
    \src[11]_i_1 
       (.I0(din[11]),
        .I1(r_a0),
        .I2(bw),
        .O(data4[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h2A)) 
    \src[12]_i_1 
       (.I0(din[12]),
        .I1(r_a0),
        .I2(bw),
        .O(data4[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h2A)) 
    \src[13]_i_1 
       (.I0(din[13]),
        .I1(r_a0),
        .I2(bw),
        .O(data4[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h2A)) 
    \src[14]_i_1 
       (.I0(din[14]),
        .I1(r_a0),
        .I2(bw),
        .O(data4[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \src[15]_i_1 
       (.I0(state[2]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[0]),
        .I4(state[1]),
        .I5(halt),
        .O(src0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h70)) 
    \src[15]_i_2 
       (.I0(r_a0),
        .I1(bw),
        .I2(din[15]),
        .O(src));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \src[15]_i_3 
       (.I0(rst),
        .O(\src[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBF80)) 
    \src[1]_i_1 
       (.I0(din[9]),
        .I1(r_a0),
        .I2(bw),
        .I3(din[1]),
        .O(data4[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEA2A)) 
    \src[2]_i_1 
       (.I0(din[2]),
        .I1(bw),
        .I2(r_a0),
        .I3(din[10]),
        .O(data4[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEA2A)) 
    \src[3]_i_1 
       (.I0(din[3]),
        .I1(bw),
        .I2(r_a0),
        .I3(din[11]),
        .O(data4[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEA2A)) 
    \src[4]_i_1 
       (.I0(din[4]),
        .I1(bw),
        .I2(r_a0),
        .I3(din[12]),
        .O(data4[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEA2A)) 
    \src[5]_i_1 
       (.I0(din[5]),
        .I1(bw),
        .I2(r_a0),
        .I3(din[13]),
        .O(data4[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEA2A)) 
    \src[6]_i_1 
       (.I0(din[6]),
        .I1(bw),
        .I2(r_a0),
        .I3(din[14]),
        .O(data4[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEA2A)) 
    \src[7]_i_1 
       (.I0(din[7]),
        .I1(bw),
        .I2(r_a0),
        .I3(din[15]),
        .O(data4[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h2A)) 
    \src[8]_i_1 
       (.I0(din[8]),
        .I1(r_a0),
        .I2(bw),
        .O(data4[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \src[8]_i_2 
       (.I0(rst),
        .O(\src[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h2A)) 
    \src[9]_i_1 
       (.I0(din[9]),
        .I1(r_a0),
        .I2(bw),
        .O(data4[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[0] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[0]),
        .Q(src__0[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[10] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[10]),
        .Q(src__0[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[11] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[11]),
        .Q(src__0[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[12] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[12]),
        .Q(src__0[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[13] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[13]),
        .Q(src__0[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[14] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[14]),
        .Q(src__0[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[15] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(src),
        .Q(src__0[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[1] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[1]),
        .Q(src__0[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[2] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[2]),
        .Q(src__0[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[3] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[3]),
        .Q(src__0[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[4] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[4]),
        .Q(src__0[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[5] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[5]),
        .Q(src__0[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[6] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[6]),
        .Q(src__0[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[7] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[7]),
        .Q(src__0[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[8] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[8]_i_2_n_0 ),
        .D(data4[8]),
        .Q(src__0[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \src_reg[9] 
       (.C(clk),
        .CE(src0),
        .CLR(\src[15]_i_3_n_0 ),
        .D(data4[9]),
        .Q(src__0[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30000214)) 
    wr_INST_0
       (.I0(state[0]),
        .I1(state[4]),
        .I2(state[3]),
        .I3(state[1]),
        .I4(state[2]),
        .O(wr));
endmodule
